// Benchmark "TreeLUT" written by ABC on Fri Sep  5 17:09:39 2025

module TreeLUT ( 
    \all_features[0] , \all_features[1] , \all_features[2] ,
    \all_features[3] , \all_features[4] , \all_features[5] ,
    \all_features[6] , \all_features[7] , \all_features[8] ,
    \all_features[9] , \all_features[10] , \all_features[11] ,
    \all_features[12] , \all_features[13] , \all_features[14] ,
    \all_features[15] , \all_features[16] , \all_features[17] ,
    \all_features[18] , \all_features[19] , \all_features[20] ,
    \all_features[21] , \all_features[22] , \all_features[23] ,
    \all_features[24] , \all_features[25] , \all_features[26] ,
    \all_features[27] , \all_features[28] , \all_features[29] ,
    \all_features[30] , \all_features[31] , \all_features[32] ,
    \all_features[33] , \all_features[34] , \all_features[35] ,
    \all_features[36] , \all_features[37] , \all_features[38] ,
    \all_features[39] , \all_features[40] , \all_features[41] ,
    \all_features[42] , \all_features[43] , \all_features[44] ,
    \all_features[45] , \all_features[46] , \all_features[47] ,
    \all_features[48] , \all_features[49] , \all_features[50] ,
    \all_features[51] , \all_features[52] , \all_features[53] ,
    \all_features[54] , \all_features[55] , \all_features[56] ,
    \all_features[57] , \all_features[58] , \all_features[59] ,
    \all_features[60] , \all_features[61] , \all_features[62] ,
    \all_features[63] , \all_features[64] , \all_features[65] ,
    \all_features[66] , \all_features[67] , \all_features[68] ,
    \all_features[69] , \all_features[70] , \all_features[71] ,
    \all_features[72] , \all_features[73] , \all_features[74] ,
    \all_features[75] , \all_features[76] , \all_features[77] ,
    \all_features[78] , \all_features[79] , \all_features[80] ,
    \all_features[81] , \all_features[82] , \all_features[83] ,
    \all_features[84] , \all_features[85] , \all_features[86] ,
    \all_features[87] , \all_features[88] , \all_features[89] ,
    \all_features[90] , \all_features[91] , \all_features[92] ,
    \all_features[93] , \all_features[94] , \all_features[95] ,
    \all_features[96] , \all_features[97] , \all_features[98] ,
    \all_features[99] , \all_features[100] , \all_features[101] ,
    \all_features[102] , \all_features[103] , \all_features[104] ,
    \all_features[105] , \all_features[106] , \all_features[107] ,
    \all_features[108] , \all_features[109] , \all_features[110] ,
    \all_features[111] , \all_features[112] , \all_features[113] ,
    \all_features[114] , \all_features[115] , \all_features[116] ,
    \all_features[117] , \all_features[118] , \all_features[119] ,
    \all_features[120] , \all_features[121] , \all_features[122] ,
    \all_features[123] , \all_features[124] , \all_features[125] ,
    \all_features[126] , \all_features[127] , \all_features[128] ,
    \all_features[129] , \all_features[130] , \all_features[131] ,
    \all_features[132] , \all_features[133] , \all_features[134] ,
    \all_features[135] , \all_features[136] , \all_features[137] ,
    \all_features[138] , \all_features[139] , \all_features[140] ,
    \all_features[141] , \all_features[142] , \all_features[143] ,
    \all_features[144] , \all_features[145] , \all_features[146] ,
    \all_features[147] , \all_features[148] , \all_features[149] ,
    \all_features[150] , \all_features[151] , \all_features[152] ,
    \all_features[153] , \all_features[154] , \all_features[155] ,
    \all_features[156] , \all_features[157] , \all_features[158] ,
    \all_features[159] , \all_features[160] , \all_features[161] ,
    \all_features[162] , \all_features[163] , \all_features[164] ,
    \all_features[165] , \all_features[166] , \all_features[167] ,
    \all_features[168] , \all_features[169] , \all_features[170] ,
    \all_features[171] , \all_features[172] , \all_features[173] ,
    \all_features[174] , \all_features[175] , \all_features[176] ,
    \all_features[177] , \all_features[178] , \all_features[179] ,
    \all_features[180] , \all_features[181] , \all_features[182] ,
    \all_features[183] , \all_features[184] , \all_features[185] ,
    \all_features[186] , \all_features[187] , \all_features[188] ,
    \all_features[189] , \all_features[190] , \all_features[191] ,
    \all_features[192] , \all_features[193] , \all_features[194] ,
    \all_features[195] , \all_features[196] , \all_features[197] ,
    \all_features[198] , \all_features[199] , \all_features[200] ,
    \all_features[201] , \all_features[202] , \all_features[203] ,
    \all_features[204] , \all_features[205] , \all_features[206] ,
    \all_features[207] , \all_features[208] , \all_features[209] ,
    \all_features[210] , \all_features[211] , \all_features[212] ,
    \all_features[213] , \all_features[214] , \all_features[215] ,
    \all_features[216] , \all_features[217] , \all_features[218] ,
    \all_features[219] , \all_features[220] , \all_features[221] ,
    \all_features[222] , \all_features[223] , \all_features[224] ,
    \all_features[225] , \all_features[226] , \all_features[227] ,
    \all_features[228] , \all_features[229] , \all_features[230] ,
    \all_features[231] , \all_features[232] , \all_features[233] ,
    \all_features[234] , \all_features[235] , \all_features[236] ,
    \all_features[237] , \all_features[238] , \all_features[239] ,
    \all_features[240] , \all_features[241] , \all_features[242] ,
    \all_features[243] , \all_features[244] , \all_features[245] ,
    \all_features[246] , \all_features[247] , \all_features[248] ,
    \all_features[249] , \all_features[250] , \all_features[251] ,
    \all_features[252] , \all_features[253] , \all_features[254] ,
    \all_features[255] , \all_features[256] , \all_features[257] ,
    \all_features[258] , \all_features[259] , \all_features[260] ,
    \all_features[261] , \all_features[262] , \all_features[263] ,
    \all_features[264] , \all_features[265] , \all_features[266] ,
    \all_features[267] , \all_features[268] , \all_features[269] ,
    \all_features[270] , \all_features[271] , \all_features[272] ,
    \all_features[273] , \all_features[274] , \all_features[275] ,
    \all_features[276] , \all_features[277] , \all_features[278] ,
    \all_features[279] , \all_features[280] , \all_features[281] ,
    \all_features[282] , \all_features[283] , \all_features[284] ,
    \all_features[285] , \all_features[286] , \all_features[287] ,
    \all_features[288] , \all_features[289] , \all_features[290] ,
    \all_features[291] , \all_features[292] , \all_features[293] ,
    \all_features[294] , \all_features[295] , \all_features[296] ,
    \all_features[297] , \all_features[298] , \all_features[299] ,
    \all_features[300] , \all_features[301] , \all_features[302] ,
    \all_features[303] , \all_features[304] , \all_features[305] ,
    \all_features[306] , \all_features[307] , \all_features[308] ,
    \all_features[309] , \all_features[310] , \all_features[311] ,
    \all_features[312] , \all_features[313] , \all_features[314] ,
    \all_features[315] , \all_features[316] , \all_features[317] ,
    \all_features[318] , \all_features[319] , \all_features[320] ,
    \all_features[321] , \all_features[322] , \all_features[323] ,
    \all_features[324] , \all_features[325] , \all_features[326] ,
    \all_features[327] , \all_features[328] , \all_features[329] ,
    \all_features[330] , \all_features[331] , \all_features[332] ,
    \all_features[333] , \all_features[334] , \all_features[335] ,
    \all_features[336] , \all_features[337] , \all_features[338] ,
    \all_features[339] , \all_features[340] , \all_features[341] ,
    \all_features[342] , \all_features[343] , \all_features[344] ,
    \all_features[345] , \all_features[346] , \all_features[347] ,
    \all_features[348] , \all_features[349] , \all_features[350] ,
    \all_features[351] , \all_features[352] , \all_features[353] ,
    \all_features[354] , \all_features[355] , \all_features[356] ,
    \all_features[357] , \all_features[358] , \all_features[359] ,
    \all_features[360] , \all_features[361] , \all_features[362] ,
    \all_features[363] , \all_features[364] , \all_features[365] ,
    \all_features[366] , \all_features[367] , \all_features[368] ,
    \all_features[369] , \all_features[370] , \all_features[371] ,
    \all_features[372] , \all_features[373] , \all_features[374] ,
    \all_features[375] , \all_features[376] , \all_features[377] ,
    \all_features[378] , \all_features[379] , \all_features[380] ,
    \all_features[381] , \all_features[382] , \all_features[383] ,
    \all_features[384] , \all_features[385] , \all_features[386] ,
    \all_features[387] , \all_features[388] , \all_features[389] ,
    \all_features[390] , \all_features[391] , \all_features[392] ,
    \all_features[393] , \all_features[394] , \all_features[395] ,
    \all_features[396] , \all_features[397] , \all_features[398] ,
    \all_features[399] , \all_features[400] , \all_features[401] ,
    \all_features[402] , \all_features[403] , \all_features[404] ,
    \all_features[405] , \all_features[406] , \all_features[407] ,
    \all_features[408] , \all_features[409] , \all_features[410] ,
    \all_features[411] , \all_features[412] , \all_features[413] ,
    \all_features[414] , \all_features[415] , \all_features[416] ,
    \all_features[417] , \all_features[418] , \all_features[419] ,
    \all_features[420] , \all_features[421] , \all_features[422] ,
    \all_features[423] , \all_features[424] , \all_features[425] ,
    \all_features[426] , \all_features[427] , \all_features[428] ,
    \all_features[429] , \all_features[430] , \all_features[431] ,
    \all_features[432] , \all_features[433] , \all_features[434] ,
    \all_features[435] , \all_features[436] , \all_features[437] ,
    \all_features[438] , \all_features[439] , \all_features[440] ,
    \all_features[441] , \all_features[442] , \all_features[443] ,
    \all_features[444] , \all_features[445] , \all_features[446] ,
    \all_features[447] , \all_features[448] , \all_features[449] ,
    \all_features[450] , \all_features[451] , \all_features[452] ,
    \all_features[453] , \all_features[454] , \all_features[455] ,
    \all_features[456] , \all_features[457] , \all_features[458] ,
    \all_features[459] , \all_features[460] , \all_features[461] ,
    \all_features[462] , \all_features[463] , \all_features[464] ,
    \all_features[465] , \all_features[466] , \all_features[467] ,
    \all_features[468] , \all_features[469] , \all_features[470] ,
    \all_features[471] , \all_features[472] , \all_features[473] ,
    \all_features[474] , \all_features[475] , \all_features[476] ,
    \all_features[477] , \all_features[478] , \all_features[479] ,
    \all_features[480] , \all_features[481] , \all_features[482] ,
    \all_features[483] , \all_features[484] , \all_features[485] ,
    \all_features[486] , \all_features[487] , \all_features[488] ,
    \all_features[489] , \all_features[490] , \all_features[491] ,
    \all_features[492] , \all_features[493] , \all_features[494] ,
    \all_features[495] , \all_features[496] , \all_features[497] ,
    \all_features[498] , \all_features[499] , \all_features[500] ,
    \all_features[501] , \all_features[502] , \all_features[503] ,
    \all_features[504] , \all_features[505] , \all_features[506] ,
    \all_features[507] , \all_features[508] , \all_features[509] ,
    \all_features[510] , \all_features[511] , \all_features[512] ,
    \all_features[513] , \all_features[514] , \all_features[515] ,
    \all_features[516] , \all_features[517] , \all_features[518] ,
    \all_features[519] , \all_features[520] , \all_features[521] ,
    \all_features[522] , \all_features[523] , \all_features[524] ,
    \all_features[525] , \all_features[526] , \all_features[527] ,
    \all_features[528] , \all_features[529] , \all_features[530] ,
    \all_features[531] , \all_features[532] , \all_features[533] ,
    \all_features[534] , \all_features[535] , \all_features[536] ,
    \all_features[537] , \all_features[538] , \all_features[539] ,
    \all_features[540] , \all_features[541] , \all_features[542] ,
    \all_features[543] , \all_features[544] , \all_features[545] ,
    \all_features[546] , \all_features[547] , \all_features[548] ,
    \all_features[549] , \all_features[550] , \all_features[551] ,
    \all_features[552] , \all_features[553] , \all_features[554] ,
    \all_features[555] , \all_features[556] , \all_features[557] ,
    \all_features[558] , \all_features[559] , \all_features[560] ,
    \all_features[561] , \all_features[562] , \all_features[563] ,
    \all_features[564] , \all_features[565] , \all_features[566] ,
    \all_features[567] , \all_features[568] , \all_features[569] ,
    \all_features[570] , \all_features[571] , \all_features[572] ,
    \all_features[573] , \all_features[574] , \all_features[575] ,
    \all_features[576] , \all_features[577] , \all_features[578] ,
    \all_features[579] , \all_features[580] , \all_features[581] ,
    \all_features[582] , \all_features[583] , \all_features[584] ,
    \all_features[585] , \all_features[586] , \all_features[587] ,
    \all_features[588] , \all_features[589] , \all_features[590] ,
    \all_features[591] , \all_features[592] , \all_features[593] ,
    \all_features[594] , \all_features[595] , \all_features[596] ,
    \all_features[597] , \all_features[598] , \all_features[599] ,
    \all_features[600] , \all_features[601] , \all_features[602] ,
    \all_features[603] , \all_features[604] , \all_features[605] ,
    \all_features[606] , \all_features[607] , \all_features[608] ,
    \all_features[609] , \all_features[610] , \all_features[611] ,
    \all_features[612] , \all_features[613] , \all_features[614] ,
    \all_features[615] , \all_features[616] , \all_features[617] ,
    \all_features[618] , \all_features[619] , \all_features[620] ,
    \all_features[621] , \all_features[622] , \all_features[623] ,
    \all_features[624] , \all_features[625] , \all_features[626] ,
    \all_features[627] , \all_features[628] , \all_features[629] ,
    \all_features[630] , \all_features[631] , \all_features[632] ,
    \all_features[633] , \all_features[634] , \all_features[635] ,
    \all_features[636] , \all_features[637] , \all_features[638] ,
    \all_features[639] , \all_features[640] , \all_features[641] ,
    \all_features[642] , \all_features[643] , \all_features[644] ,
    \all_features[645] , \all_features[646] , \all_features[647] ,
    \all_features[648] , \all_features[649] , \all_features[650] ,
    \all_features[651] , \all_features[652] , \all_features[653] ,
    \all_features[654] , \all_features[655] , \all_features[656] ,
    \all_features[657] , \all_features[658] , \all_features[659] ,
    \all_features[660] , \all_features[661] , \all_features[662] ,
    \all_features[663] , \all_features[664] , \all_features[665] ,
    \all_features[666] , \all_features[667] , \all_features[668] ,
    \all_features[669] , \all_features[670] , \all_features[671] ,
    \all_features[672] , \all_features[673] , \all_features[674] ,
    \all_features[675] , \all_features[676] , \all_features[677] ,
    \all_features[678] , \all_features[679] , \all_features[680] ,
    \all_features[681] , \all_features[682] , \all_features[683] ,
    \all_features[684] , \all_features[685] , \all_features[686] ,
    \all_features[687] , \all_features[688] , \all_features[689] ,
    \all_features[690] , \all_features[691] , \all_features[692] ,
    \all_features[693] , \all_features[694] , \all_features[695] ,
    \all_features[696] , \all_features[697] , \all_features[698] ,
    \all_features[699] , \all_features[700] , \all_features[701] ,
    \all_features[702] , \all_features[703] , \all_features[704] ,
    \all_features[705] , \all_features[706] , \all_features[707] ,
    \all_features[708] , \all_features[709] , \all_features[710] ,
    \all_features[711] , \all_features[712] , \all_features[713] ,
    \all_features[714] , \all_features[715] , \all_features[716] ,
    \all_features[717] , \all_features[718] , \all_features[719] ,
    \all_features[720] , \all_features[721] , \all_features[722] ,
    \all_features[723] , \all_features[724] , \all_features[725] ,
    \all_features[726] , \all_features[727] , \all_features[728] ,
    \all_features[729] , \all_features[730] , \all_features[731] ,
    \all_features[732] , \all_features[733] , \all_features[734] ,
    \all_features[735] , \all_features[736] , \all_features[737] ,
    \all_features[738] , \all_features[739] , \all_features[740] ,
    \all_features[741] , \all_features[742] , \all_features[743] ,
    \all_features[744] , \all_features[745] , \all_features[746] ,
    \all_features[747] , \all_features[748] , \all_features[749] ,
    \all_features[750] , \all_features[751] , \all_features[752] ,
    \all_features[753] , \all_features[754] , \all_features[755] ,
    \all_features[756] , \all_features[757] , \all_features[758] ,
    \all_features[759] , \all_features[760] , \all_features[761] ,
    \all_features[762] , \all_features[763] , \all_features[764] ,
    \all_features[765] , \all_features[766] , \all_features[767] ,
    \all_features[768] , \all_features[769] , \all_features[770] ,
    \all_features[771] , \all_features[772] , \all_features[773] ,
    \all_features[774] , \all_features[775] , \all_features[776] ,
    \all_features[777] , \all_features[778] , \all_features[779] ,
    \all_features[780] , \all_features[781] , \all_features[782] ,
    \all_features[783] , \all_features[784] , \all_features[785] ,
    \all_features[786] , \all_features[787] , \all_features[788] ,
    \all_features[789] , \all_features[790] , \all_features[791] ,
    \all_features[792] , \all_features[793] , \all_features[794] ,
    \all_features[795] , \all_features[796] , \all_features[797] ,
    \all_features[798] , \all_features[799] , \all_features[800] ,
    \all_features[801] , \all_features[802] , \all_features[803] ,
    \all_features[804] , \all_features[805] , \all_features[806] ,
    \all_features[807] , \all_features[808] , \all_features[809] ,
    \all_features[810] , \all_features[811] , \all_features[812] ,
    \all_features[813] , \all_features[814] , \all_features[815] ,
    \all_features[816] , \all_features[817] , \all_features[818] ,
    \all_features[819] , \all_features[820] , \all_features[821] ,
    \all_features[822] , \all_features[823] , \all_features[824] ,
    \all_features[825] , \all_features[826] , \all_features[827] ,
    \all_features[828] , \all_features[829] , \all_features[830] ,
    \all_features[831] , \all_features[832] , \all_features[833] ,
    \all_features[834] , \all_features[835] , \all_features[836] ,
    \all_features[837] , \all_features[838] , \all_features[839] ,
    \all_features[840] , \all_features[841] , \all_features[842] ,
    \all_features[843] , \all_features[844] , \all_features[845] ,
    \all_features[846] , \all_features[847] , \all_features[848] ,
    \all_features[849] , \all_features[850] , \all_features[851] ,
    \all_features[852] , \all_features[853] , \all_features[854] ,
    \all_features[855] , \all_features[856] , \all_features[857] ,
    \all_features[858] , \all_features[859] , \all_features[860] ,
    \all_features[861] , \all_features[862] , \all_features[863] ,
    \all_features[864] , \all_features[865] , \all_features[866] ,
    \all_features[867] , \all_features[868] , \all_features[869] ,
    \all_features[870] , \all_features[871] , \all_features[872] ,
    \all_features[873] , \all_features[874] , \all_features[875] ,
    \all_features[876] , \all_features[877] , \all_features[878] ,
    \all_features[879] , \all_features[880] , \all_features[881] ,
    \all_features[882] , \all_features[883] , \all_features[884] ,
    \all_features[885] , \all_features[886] , \all_features[887] ,
    \all_features[888] , \all_features[889] , \all_features[890] ,
    \all_features[891] , \all_features[892] , \all_features[893] ,
    \all_features[894] , \all_features[895] , \all_features[896] ,
    \all_features[897] , \all_features[898] , \all_features[899] ,
    \all_features[900] , \all_features[901] , \all_features[902] ,
    \all_features[903] , \all_features[904] , \all_features[905] ,
    \all_features[906] , \all_features[907] , \all_features[908] ,
    \all_features[909] , \all_features[910] , \all_features[911] ,
    \all_features[912] , \all_features[913] , \all_features[914] ,
    \all_features[915] , \all_features[916] , \all_features[917] ,
    \all_features[918] , \all_features[919] , \all_features[920] ,
    \all_features[921] , \all_features[922] , \all_features[923] ,
    \all_features[924] , \all_features[925] , \all_features[926] ,
    \all_features[927] , \all_features[928] , \all_features[929] ,
    \all_features[930] , \all_features[931] , \all_features[932] ,
    \all_features[933] , \all_features[934] , \all_features[935] ,
    \all_features[936] , \all_features[937] , \all_features[938] ,
    \all_features[939] , \all_features[940] , \all_features[941] ,
    \all_features[942] , \all_features[943] , \all_features[944] ,
    \all_features[945] , \all_features[946] , \all_features[947] ,
    \all_features[948] , \all_features[949] , \all_features[950] ,
    \all_features[951] , \all_features[952] , \all_features[953] ,
    \all_features[954] , \all_features[955] , \all_features[956] ,
    \all_features[957] , \all_features[958] , \all_features[959] ,
    \all_features[960] , \all_features[961] , \all_features[962] ,
    \all_features[963] , \all_features[964] , \all_features[965] ,
    \all_features[966] , \all_features[967] , \all_features[968] ,
    \all_features[969] , \all_features[970] , \all_features[971] ,
    \all_features[972] , \all_features[973] , \all_features[974] ,
    \all_features[975] , \all_features[976] , \all_features[977] ,
    \all_features[978] , \all_features[979] , \all_features[980] ,
    \all_features[981] , \all_features[982] , \all_features[983] ,
    \all_features[984] , \all_features[985] , \all_features[986] ,
    \all_features[987] , \all_features[988] , \all_features[989] ,
    \all_features[990] , \all_features[991] , \all_features[992] ,
    \all_features[993] , \all_features[994] , \all_features[995] ,
    \all_features[996] , \all_features[997] , \all_features[998] ,
    \all_features[999] , \all_features[1000] , \all_features[1001] ,
    \all_features[1002] , \all_features[1003] , \all_features[1004] ,
    \all_features[1005] , \all_features[1006] , \all_features[1007] ,
    \all_features[1008] , \all_features[1009] , \all_features[1010] ,
    \all_features[1011] , \all_features[1012] , \all_features[1013] ,
    \all_features[1014] , \all_features[1015] , \all_features[1016] ,
    \all_features[1017] , \all_features[1018] , \all_features[1019] ,
    \all_features[1020] , \all_features[1021] , \all_features[1022] ,
    \all_features[1023] , \all_features[1024] , \all_features[1025] ,
    \all_features[1026] , \all_features[1027] , \all_features[1028] ,
    \all_features[1029] , \all_features[1030] , \all_features[1031] ,
    \all_features[1032] , \all_features[1033] , \all_features[1034] ,
    \all_features[1035] , \all_features[1036] , \all_features[1037] ,
    \all_features[1038] , \all_features[1039] , \all_features[1040] ,
    \all_features[1041] , \all_features[1042] , \all_features[1043] ,
    \all_features[1044] , \all_features[1045] , \all_features[1046] ,
    \all_features[1047] , \all_features[1048] , \all_features[1049] ,
    \all_features[1050] , \all_features[1051] , \all_features[1052] ,
    \all_features[1053] , \all_features[1054] , \all_features[1055] ,
    \all_features[1056] , \all_features[1057] , \all_features[1058] ,
    \all_features[1059] , \all_features[1060] , \all_features[1061] ,
    \all_features[1062] , \all_features[1063] , \all_features[1064] ,
    \all_features[1065] , \all_features[1066] , \all_features[1067] ,
    \all_features[1068] , \all_features[1069] , \all_features[1070] ,
    \all_features[1071] , \all_features[1072] , \all_features[1073] ,
    \all_features[1074] , \all_features[1075] , \all_features[1076] ,
    \all_features[1077] , \all_features[1078] , \all_features[1079] ,
    \all_features[1080] , \all_features[1081] , \all_features[1082] ,
    \all_features[1083] , \all_features[1084] , \all_features[1085] ,
    \all_features[1086] , \all_features[1087] , \all_features[1088] ,
    \all_features[1089] , \all_features[1090] , \all_features[1091] ,
    \all_features[1092] , \all_features[1093] , \all_features[1094] ,
    \all_features[1095] , \all_features[1096] , \all_features[1097] ,
    \all_features[1098] , \all_features[1099] , \all_features[1100] ,
    \all_features[1101] , \all_features[1102] , \all_features[1103] ,
    \all_features[1104] , \all_features[1105] , \all_features[1106] ,
    \all_features[1107] , \all_features[1108] , \all_features[1109] ,
    \all_features[1110] , \all_features[1111] , \all_features[1112] ,
    \all_features[1113] , \all_features[1114] , \all_features[1115] ,
    \all_features[1116] , \all_features[1117] , \all_features[1118] ,
    \all_features[1119] , \all_features[1120] , \all_features[1121] ,
    \all_features[1122] , \all_features[1123] , \all_features[1124] ,
    \all_features[1125] , \all_features[1126] , \all_features[1127] ,
    \all_features[1128] , \all_features[1129] , \all_features[1130] ,
    \all_features[1131] , \all_features[1132] , \all_features[1133] ,
    \all_features[1134] , \all_features[1135] , \all_features[1136] ,
    \all_features[1137] , \all_features[1138] , \all_features[1139] ,
    \all_features[1140] , \all_features[1141] , \all_features[1142] ,
    \all_features[1143] , \all_features[1144] , \all_features[1145] ,
    \all_features[1146] , \all_features[1147] , \all_features[1148] ,
    \all_features[1149] , \all_features[1150] , \all_features[1151] ,
    \all_features[1152] , \all_features[1153] , \all_features[1154] ,
    \all_features[1155] , \all_features[1156] , \all_features[1157] ,
    \all_features[1158] , \all_features[1159] , \all_features[1160] ,
    \all_features[1161] , \all_features[1162] , \all_features[1163] ,
    \all_features[1164] , \all_features[1165] , \all_features[1166] ,
    \all_features[1167] , \all_features[1168] , \all_features[1169] ,
    \all_features[1170] , \all_features[1171] , \all_features[1172] ,
    \all_features[1173] , \all_features[1174] , \all_features[1175] ,
    \all_features[1176] , \all_features[1177] , \all_features[1178] ,
    \all_features[1179] , \all_features[1180] , \all_features[1181] ,
    \all_features[1182] , \all_features[1183] , \all_features[1184] ,
    \all_features[1185] , \all_features[1186] , \all_features[1187] ,
    \all_features[1188] , \all_features[1189] , \all_features[1190] ,
    \all_features[1191] , \all_features[1192] , \all_features[1193] ,
    \all_features[1194] , \all_features[1195] , \all_features[1196] ,
    \all_features[1197] , \all_features[1198] , \all_features[1199] ,
    \all_features[1200] , \all_features[1201] , \all_features[1202] ,
    \all_features[1203] , \all_features[1204] , \all_features[1205] ,
    \all_features[1206] , \all_features[1207] , \all_features[1208] ,
    \all_features[1209] , \all_features[1210] , \all_features[1211] ,
    \all_features[1212] , \all_features[1213] , \all_features[1214] ,
    \all_features[1215] , \all_features[1216] , \all_features[1217] ,
    \all_features[1218] , \all_features[1219] , \all_features[1220] ,
    \all_features[1221] , \all_features[1222] , \all_features[1223] ,
    \all_features[1224] , \all_features[1225] , \all_features[1226] ,
    \all_features[1227] , \all_features[1228] , \all_features[1229] ,
    \all_features[1230] , \all_features[1231] , \all_features[1232] ,
    \all_features[1233] , \all_features[1234] , \all_features[1235] ,
    \all_features[1236] , \all_features[1237] , \all_features[1238] ,
    \all_features[1239] , \all_features[1240] , \all_features[1241] ,
    \all_features[1242] , \all_features[1243] , \all_features[1244] ,
    \all_features[1245] , \all_features[1246] , \all_features[1247] ,
    \all_features[1248] , \all_features[1249] , \all_features[1250] ,
    \all_features[1251] , \all_features[1252] , \all_features[1253] ,
    \all_features[1254] , \all_features[1255] , \all_features[1256] ,
    \all_features[1257] , \all_features[1258] , \all_features[1259] ,
    \all_features[1260] , \all_features[1261] , \all_features[1262] ,
    \all_features[1263] , \all_features[1264] , \all_features[1265] ,
    \all_features[1266] , \all_features[1267] , \all_features[1268] ,
    \all_features[1269] , \all_features[1270] , \all_features[1271] ,
    \all_features[1272] , \all_features[1273] , \all_features[1274] ,
    \all_features[1275] , \all_features[1276] , \all_features[1277] ,
    \all_features[1278] , \all_features[1279] , \all_features[1280] ,
    \all_features[1281] , \all_features[1282] , \all_features[1283] ,
    \all_features[1284] , \all_features[1285] , \all_features[1286] ,
    \all_features[1287] , \all_features[1288] , \all_features[1289] ,
    \all_features[1290] , \all_features[1291] , \all_features[1292] ,
    \all_features[1293] , \all_features[1294] , \all_features[1295] ,
    \all_features[1296] , \all_features[1297] , \all_features[1298] ,
    \all_features[1299] , \all_features[1300] , \all_features[1301] ,
    \all_features[1302] , \all_features[1303] , \all_features[1304] ,
    \all_features[1305] , \all_features[1306] , \all_features[1307] ,
    \all_features[1308] , \all_features[1309] , \all_features[1310] ,
    \all_features[1311] , \all_features[1312] , \all_features[1313] ,
    \all_features[1314] , \all_features[1315] , \all_features[1316] ,
    \all_features[1317] , \all_features[1318] , \all_features[1319] ,
    \all_features[1320] , \all_features[1321] , \all_features[1322] ,
    \all_features[1323] , \all_features[1324] , \all_features[1325] ,
    \all_features[1326] , \all_features[1327] , \all_features[1328] ,
    \all_features[1329] , \all_features[1330] , \all_features[1331] ,
    \all_features[1332] , \all_features[1333] , \all_features[1334] ,
    \all_features[1335] , \all_features[1336] , \all_features[1337] ,
    \all_features[1338] , \all_features[1339] , \all_features[1340] ,
    \all_features[1341] , \all_features[1342] , \all_features[1343] ,
    \all_features[1344] , \all_features[1345] , \all_features[1346] ,
    \all_features[1347] , \all_features[1348] , \all_features[1349] ,
    \all_features[1350] , \all_features[1351] , \all_features[1352] ,
    \all_features[1353] , \all_features[1354] , \all_features[1355] ,
    \all_features[1356] , \all_features[1357] , \all_features[1358] ,
    \all_features[1359] , \all_features[1360] , \all_features[1361] ,
    \all_features[1362] , \all_features[1363] , \all_features[1364] ,
    \all_features[1365] , \all_features[1366] , \all_features[1367] ,
    \all_features[1368] , \all_features[1369] , \all_features[1370] ,
    \all_features[1371] , \all_features[1372] , \all_features[1373] ,
    \all_features[1374] , \all_features[1375] , \all_features[1376] ,
    \all_features[1377] , \all_features[1378] , \all_features[1379] ,
    \all_features[1380] , \all_features[1381] , \all_features[1382] ,
    \all_features[1383] , \all_features[1384] , \all_features[1385] ,
    \all_features[1386] , \all_features[1387] , \all_features[1388] ,
    \all_features[1389] , \all_features[1390] , \all_features[1391] ,
    \all_features[1392] , \all_features[1393] , \all_features[1394] ,
    \all_features[1395] , \all_features[1396] , \all_features[1397] ,
    \all_features[1398] , \all_features[1399] , \all_features[1400] ,
    \all_features[1401] , \all_features[1402] , \all_features[1403] ,
    \all_features[1404] , \all_features[1405] , \all_features[1406] ,
    \all_features[1407] , \all_features[1408] , \all_features[1409] ,
    \all_features[1410] , \all_features[1411] , \all_features[1412] ,
    \all_features[1413] , \all_features[1414] , \all_features[1415] ,
    \all_features[1416] , \all_features[1417] , \all_features[1418] ,
    \all_features[1419] , \all_features[1420] , \all_features[1421] ,
    \all_features[1422] , \all_features[1423] , \all_features[1424] ,
    \all_features[1425] , \all_features[1426] , \all_features[1427] ,
    \all_features[1428] , \all_features[1429] , \all_features[1430] ,
    \all_features[1431] , \all_features[1432] , \all_features[1433] ,
    \all_features[1434] , \all_features[1435] , \all_features[1436] ,
    \all_features[1437] , \all_features[1438] , \all_features[1439] ,
    \all_features[1440] , \all_features[1441] , \all_features[1442] ,
    \all_features[1443] , \all_features[1444] , \all_features[1445] ,
    \all_features[1446] , \all_features[1447] , \all_features[1448] ,
    \all_features[1449] , \all_features[1450] , \all_features[1451] ,
    \all_features[1452] , \all_features[1453] , \all_features[1454] ,
    \all_features[1455] , \all_features[1456] , \all_features[1457] ,
    \all_features[1458] , \all_features[1459] , \all_features[1460] ,
    \all_features[1461] , \all_features[1462] , \all_features[1463] ,
    \all_features[1464] , \all_features[1465] , \all_features[1466] ,
    \all_features[1467] , \all_features[1468] , \all_features[1469] ,
    \all_features[1470] , \all_features[1471] , \all_features[1472] ,
    \all_features[1473] , \all_features[1474] , \all_features[1475] ,
    \all_features[1476] , \all_features[1477] , \all_features[1478] ,
    \all_features[1479] , \all_features[1480] , \all_features[1481] ,
    \all_features[1482] , \all_features[1483] , \all_features[1484] ,
    \all_features[1485] , \all_features[1486] , \all_features[1487] ,
    \all_features[1488] , \all_features[1489] , \all_features[1490] ,
    \all_features[1491] , \all_features[1492] , \all_features[1493] ,
    \all_features[1494] , \all_features[1495] , \all_features[1496] ,
    \all_features[1497] , \all_features[1498] , \all_features[1499] ,
    \all_features[1500] , \all_features[1501] , \all_features[1502] ,
    \all_features[1503] , \all_features[1504] , \all_features[1505] ,
    \all_features[1506] , \all_features[1507] , \all_features[1508] ,
    \all_features[1509] , \all_features[1510] , \all_features[1511] ,
    \all_features[1512] , \all_features[1513] , \all_features[1514] ,
    \all_features[1515] , \all_features[1516] , \all_features[1517] ,
    \all_features[1518] , \all_features[1519] , \all_features[1520] ,
    \all_features[1521] , \all_features[1522] , \all_features[1523] ,
    \all_features[1524] , \all_features[1525] , \all_features[1526] ,
    \all_features[1527] , \all_features[1528] , \all_features[1529] ,
    \all_features[1530] , \all_features[1531] , \all_features[1532] ,
    \all_features[1533] , \all_features[1534] , \all_features[1535] ,
    \all_features[1536] , \all_features[1537] , \all_features[1538] ,
    \all_features[1539] , \all_features[1540] , \all_features[1541] ,
    \all_features[1542] , \all_features[1543] , \all_features[1544] ,
    \all_features[1545] , \all_features[1546] , \all_features[1547] ,
    \all_features[1548] , \all_features[1549] , \all_features[1550] ,
    \all_features[1551] , \all_features[1552] , \all_features[1553] ,
    \all_features[1554] , \all_features[1555] , \all_features[1556] ,
    \all_features[1557] , \all_features[1558] , \all_features[1559] ,
    \all_features[1560] , \all_features[1561] , \all_features[1562] ,
    \all_features[1563] , \all_features[1564] , \all_features[1565] ,
    \all_features[1566] , \all_features[1567] , \all_features[1568] ,
    \all_features[1569] , \all_features[1570] , \all_features[1571] ,
    \all_features[1572] , \all_features[1573] , \all_features[1574] ,
    \all_features[1575] , \all_features[1576] , \all_features[1577] ,
    \all_features[1578] , \all_features[1579] , \all_features[1580] ,
    \all_features[1581] , \all_features[1582] , \all_features[1583] ,
    \all_features[1584] , \all_features[1585] , \all_features[1586] ,
    \all_features[1587] , \all_features[1588] , \all_features[1589] ,
    \all_features[1590] , \all_features[1591] , \all_features[1592] ,
    \all_features[1593] , \all_features[1594] , \all_features[1595] ,
    \all_features[1596] , \all_features[1597] , \all_features[1598] ,
    \all_features[1599] , \all_features[1600] , \all_features[1601] ,
    \all_features[1602] , \all_features[1603] , \all_features[1604] ,
    \all_features[1605] , \all_features[1606] , \all_features[1607] ,
    \all_features[1608] , \all_features[1609] , \all_features[1610] ,
    \all_features[1611] , \all_features[1612] , \all_features[1613] ,
    \all_features[1614] , \all_features[1615] , \all_features[1616] ,
    \all_features[1617] , \all_features[1618] , \all_features[1619] ,
    \all_features[1620] , \all_features[1621] , \all_features[1622] ,
    \all_features[1623] , \all_features[1624] , \all_features[1625] ,
    \all_features[1626] , \all_features[1627] , \all_features[1628] ,
    \all_features[1629] , \all_features[1630] , \all_features[1631] ,
    \all_features[1632] , \all_features[1633] , \all_features[1634] ,
    \all_features[1635] , \all_features[1636] , \all_features[1637] ,
    \all_features[1638] , \all_features[1639] , \all_features[1640] ,
    \all_features[1641] , \all_features[1642] , \all_features[1643] ,
    \all_features[1644] , \all_features[1645] , \all_features[1646] ,
    \all_features[1647] , \all_features[1648] , \all_features[1649] ,
    \all_features[1650] , \all_features[1651] , \all_features[1652] ,
    \all_features[1653] , \all_features[1654] , \all_features[1655] ,
    \all_features[1656] , \all_features[1657] , \all_features[1658] ,
    \all_features[1659] , \all_features[1660] , \all_features[1661] ,
    \all_features[1662] , \all_features[1663] , \all_features[1664] ,
    \all_features[1665] , \all_features[1666] , \all_features[1667] ,
    \all_features[1668] , \all_features[1669] , \all_features[1670] ,
    \all_features[1671] , \all_features[1672] , \all_features[1673] ,
    \all_features[1674] , \all_features[1675] , \all_features[1676] ,
    \all_features[1677] , \all_features[1678] , \all_features[1679] ,
    \all_features[1680] , \all_features[1681] , \all_features[1682] ,
    \all_features[1683] , \all_features[1684] , \all_features[1685] ,
    \all_features[1686] , \all_features[1687] , \all_features[1688] ,
    \all_features[1689] , \all_features[1690] , \all_features[1691] ,
    \all_features[1692] , \all_features[1693] , \all_features[1694] ,
    \all_features[1695] , \all_features[1696] , \all_features[1697] ,
    \all_features[1698] , \all_features[1699] , \all_features[1700] ,
    \all_features[1701] , \all_features[1702] , \all_features[1703] ,
    \all_features[1704] , \all_features[1705] , \all_features[1706] ,
    \all_features[1707] , \all_features[1708] , \all_features[1709] ,
    \all_features[1710] , \all_features[1711] , \all_features[1712] ,
    \all_features[1713] , \all_features[1714] , \all_features[1715] ,
    \all_features[1716] , \all_features[1717] , \all_features[1718] ,
    \all_features[1719] , \all_features[1720] , \all_features[1721] ,
    \all_features[1722] , \all_features[1723] , \all_features[1724] ,
    \all_features[1725] , \all_features[1726] , \all_features[1727] ,
    \all_features[1728] , \all_features[1729] , \all_features[1730] ,
    \all_features[1731] , \all_features[1732] , \all_features[1733] ,
    \all_features[1734] , \all_features[1735] , \all_features[1736] ,
    \all_features[1737] , \all_features[1738] , \all_features[1739] ,
    \all_features[1740] , \all_features[1741] , \all_features[1742] ,
    \all_features[1743] , \all_features[1744] , \all_features[1745] ,
    \all_features[1746] , \all_features[1747] , \all_features[1748] ,
    \all_features[1749] , \all_features[1750] , \all_features[1751] ,
    \all_features[1752] , \all_features[1753] , \all_features[1754] ,
    \all_features[1755] , \all_features[1756] , \all_features[1757] ,
    \all_features[1758] , \all_features[1759] , \all_features[1760] ,
    \all_features[1761] , \all_features[1762] , \all_features[1763] ,
    \all_features[1764] , \all_features[1765] , \all_features[1766] ,
    \all_features[1767] , \all_features[1768] , \all_features[1769] ,
    \all_features[1770] , \all_features[1771] , \all_features[1772] ,
    \all_features[1773] , \all_features[1774] , \all_features[1775] ,
    \all_features[1776] , \all_features[1777] , \all_features[1778] ,
    \all_features[1779] , \all_features[1780] , \all_features[1781] ,
    \all_features[1782] , \all_features[1783] , \all_features[1784] ,
    \all_features[1785] , \all_features[1786] , \all_features[1787] ,
    \all_features[1788] , \all_features[1789] , \all_features[1790] ,
    \all_features[1791] , \all_features[1792] , \all_features[1793] ,
    \all_features[1794] , \all_features[1795] , \all_features[1796] ,
    \all_features[1797] , \all_features[1798] , \all_features[1799] ,
    \all_features[1800] , \all_features[1801] , \all_features[1802] ,
    \all_features[1803] , \all_features[1804] , \all_features[1805] ,
    \all_features[1806] , \all_features[1807] , \all_features[1808] ,
    \all_features[1809] , \all_features[1810] , \all_features[1811] ,
    \all_features[1812] , \all_features[1813] , \all_features[1814] ,
    \all_features[1815] , \all_features[1816] , \all_features[1817] ,
    \all_features[1818] , \all_features[1819] , \all_features[1820] ,
    \all_features[1821] , \all_features[1822] , \all_features[1823] ,
    \all_features[1824] , \all_features[1825] , \all_features[1826] ,
    \all_features[1827] , \all_features[1828] , \all_features[1829] ,
    \all_features[1830] , \all_features[1831] , \all_features[1832] ,
    \all_features[1833] , \all_features[1834] , \all_features[1835] ,
    \all_features[1836] , \all_features[1837] , \all_features[1838] ,
    \all_features[1839] , \all_features[1840] , \all_features[1841] ,
    \all_features[1842] , \all_features[1843] , \all_features[1844] ,
    \all_features[1845] , \all_features[1846] , \all_features[1847] ,
    \all_features[1848] , \all_features[1849] , \all_features[1850] ,
    \all_features[1851] , \all_features[1852] , \all_features[1853] ,
    \all_features[1854] , \all_features[1855] , \all_features[1856] ,
    \all_features[1857] , \all_features[1858] , \all_features[1859] ,
    \all_features[1860] , \all_features[1861] , \all_features[1862] ,
    \all_features[1863] , \all_features[1864] , \all_features[1865] ,
    \all_features[1866] , \all_features[1867] , \all_features[1868] ,
    \all_features[1869] , \all_features[1870] , \all_features[1871] ,
    \all_features[1872] , \all_features[1873] , \all_features[1874] ,
    \all_features[1875] , \all_features[1876] , \all_features[1877] ,
    \all_features[1878] , \all_features[1879] , \all_features[1880] ,
    \all_features[1881] , \all_features[1882] , \all_features[1883] ,
    \all_features[1884] , \all_features[1885] , \all_features[1886] ,
    \all_features[1887] , \all_features[1888] , \all_features[1889] ,
    \all_features[1890] , \all_features[1891] , \all_features[1892] ,
    \all_features[1893] , \all_features[1894] , \all_features[1895] ,
    \all_features[1896] , \all_features[1897] , \all_features[1898] ,
    \all_features[1899] , \all_features[1900] , \all_features[1901] ,
    \all_features[1902] , \all_features[1903] , \all_features[1904] ,
    \all_features[1905] , \all_features[1906] , \all_features[1907] ,
    \all_features[1908] , \all_features[1909] , \all_features[1910] ,
    \all_features[1911] , \all_features[1912] , \all_features[1913] ,
    \all_features[1914] , \all_features[1915] , \all_features[1916] ,
    \all_features[1917] , \all_features[1918] , \all_features[1919] ,
    \all_features[1920] , \all_features[1921] , \all_features[1922] ,
    \all_features[1923] , \all_features[1924] , \all_features[1925] ,
    \all_features[1926] , \all_features[1927] , \all_features[1928] ,
    \all_features[1929] , \all_features[1930] , \all_features[1931] ,
    \all_features[1932] , \all_features[1933] , \all_features[1934] ,
    \all_features[1935] , \all_features[1936] , \all_features[1937] ,
    \all_features[1938] , \all_features[1939] , \all_features[1940] ,
    \all_features[1941] , \all_features[1942] , \all_features[1943] ,
    \all_features[1944] , \all_features[1945] , \all_features[1946] ,
    \all_features[1947] , \all_features[1948] , \all_features[1949] ,
    \all_features[1950] , \all_features[1951] , \all_features[1952] ,
    \all_features[1953] , \all_features[1954] , \all_features[1955] ,
    \all_features[1956] , \all_features[1957] , \all_features[1958] ,
    \all_features[1959] , \all_features[1960] , \all_features[1961] ,
    \all_features[1962] , \all_features[1963] , \all_features[1964] ,
    \all_features[1965] , \all_features[1966] , \all_features[1967] ,
    \all_features[1968] , \all_features[1969] , \all_features[1970] ,
    \all_features[1971] , \all_features[1972] , \all_features[1973] ,
    \all_features[1974] , \all_features[1975] , \all_features[1976] ,
    \all_features[1977] , \all_features[1978] , \all_features[1979] ,
    \all_features[1980] , \all_features[1981] , \all_features[1982] ,
    \all_features[1983] , \all_features[1984] , \all_features[1985] ,
    \all_features[1986] , \all_features[1987] , \all_features[1988] ,
    \all_features[1989] , \all_features[1990] , \all_features[1991] ,
    \all_features[1992] , \all_features[1993] , \all_features[1994] ,
    \all_features[1995] , \all_features[1996] , \all_features[1997] ,
    \all_features[1998] , \all_features[1999] , \all_features[2000] ,
    \all_features[2001] , \all_features[2002] , \all_features[2003] ,
    \all_features[2004] , \all_features[2005] , \all_features[2006] ,
    \all_features[2007] , \all_features[2008] , \all_features[2009] ,
    \all_features[2010] , \all_features[2011] , \all_features[2012] ,
    \all_features[2013] , \all_features[2014] , \all_features[2015] ,
    \all_features[2016] , \all_features[2017] , \all_features[2018] ,
    \all_features[2019] , \all_features[2020] , \all_features[2021] ,
    \all_features[2022] , \all_features[2023] , \all_features[2024] ,
    \all_features[2025] , \all_features[2026] , \all_features[2027] ,
    \all_features[2028] , \all_features[2029] , \all_features[2030] ,
    \all_features[2031] , \all_features[2032] , \all_features[2033] ,
    \all_features[2034] , \all_features[2035] , \all_features[2036] ,
    \all_features[2037] , \all_features[2038] , \all_features[2039] ,
    \all_features[2040] , \all_features[2041] , \all_features[2042] ,
    \all_features[2043] , \all_features[2044] , \all_features[2045] ,
    \all_features[2046] , \all_features[2047] , \all_features[2048] ,
    \all_features[2049] , \all_features[2050] , \all_features[2051] ,
    \all_features[2052] , \all_features[2053] , \all_features[2054] ,
    \all_features[2055] , \all_features[2056] , \all_features[2057] ,
    \all_features[2058] , \all_features[2059] , \all_features[2060] ,
    \all_features[2061] , \all_features[2062] , \all_features[2063] ,
    \all_features[2064] , \all_features[2065] , \all_features[2066] ,
    \all_features[2067] , \all_features[2068] , \all_features[2069] ,
    \all_features[2070] , \all_features[2071] , \all_features[2072] ,
    \all_features[2073] , \all_features[2074] , \all_features[2075] ,
    \all_features[2076] , \all_features[2077] , \all_features[2078] ,
    \all_features[2079] , \all_features[2080] , \all_features[2081] ,
    \all_features[2082] , \all_features[2083] , \all_features[2084] ,
    \all_features[2085] , \all_features[2086] , \all_features[2087] ,
    \all_features[2088] , \all_features[2089] , \all_features[2090] ,
    \all_features[2091] , \all_features[2092] , \all_features[2093] ,
    \all_features[2094] , \all_features[2095] , \all_features[2096] ,
    \all_features[2097] , \all_features[2098] , \all_features[2099] ,
    \all_features[2100] , \all_features[2101] , \all_features[2102] ,
    \all_features[2103] , \all_features[2104] , \all_features[2105] ,
    \all_features[2106] , \all_features[2107] , \all_features[2108] ,
    \all_features[2109] , \all_features[2110] , \all_features[2111] ,
    \all_features[2112] , \all_features[2113] , \all_features[2114] ,
    \all_features[2115] , \all_features[2116] , \all_features[2117] ,
    \all_features[2118] , \all_features[2119] , \all_features[2120] ,
    \all_features[2121] , \all_features[2122] , \all_features[2123] ,
    \all_features[2124] , \all_features[2125] , \all_features[2126] ,
    \all_features[2127] , \all_features[2128] , \all_features[2129] ,
    \all_features[2130] , \all_features[2131] , \all_features[2132] ,
    \all_features[2133] , \all_features[2134] , \all_features[2135] ,
    \all_features[2136] , \all_features[2137] , \all_features[2138] ,
    \all_features[2139] , \all_features[2140] , \all_features[2141] ,
    \all_features[2142] , \all_features[2143] , \all_features[2144] ,
    \all_features[2145] , \all_features[2146] , \all_features[2147] ,
    \all_features[2148] , \all_features[2149] , \all_features[2150] ,
    \all_features[2151] , \all_features[2152] , \all_features[2153] ,
    \all_features[2154] , \all_features[2155] , \all_features[2156] ,
    \all_features[2157] , \all_features[2158] , \all_features[2159] ,
    \all_features[2160] , \all_features[2161] , \all_features[2162] ,
    \all_features[2163] , \all_features[2164] , \all_features[2165] ,
    \all_features[2166] , \all_features[2167] , \all_features[2168] ,
    \all_features[2169] , \all_features[2170] , \all_features[2171] ,
    \all_features[2172] , \all_features[2173] , \all_features[2174] ,
    \all_features[2175] , \all_features[2176] , \all_features[2177] ,
    \all_features[2178] , \all_features[2179] , \all_features[2180] ,
    \all_features[2181] , \all_features[2182] , \all_features[2183] ,
    \all_features[2184] , \all_features[2185] , \all_features[2186] ,
    \all_features[2187] , \all_features[2188] , \all_features[2189] ,
    \all_features[2190] , \all_features[2191] , \all_features[2192] ,
    \all_features[2193] , \all_features[2194] , \all_features[2195] ,
    \all_features[2196] , \all_features[2197] , \all_features[2198] ,
    \all_features[2199] , \all_features[2200] , \all_features[2201] ,
    \all_features[2202] , \all_features[2203] , \all_features[2204] ,
    \all_features[2205] , \all_features[2206] , \all_features[2207] ,
    \all_features[2208] , \all_features[2209] , \all_features[2210] ,
    \all_features[2211] , \all_features[2212] , \all_features[2213] ,
    \all_features[2214] , \all_features[2215] , \all_features[2216] ,
    \all_features[2217] , \all_features[2218] , \all_features[2219] ,
    \all_features[2220] , \all_features[2221] , \all_features[2222] ,
    \all_features[2223] , \all_features[2224] , \all_features[2225] ,
    \all_features[2226] , \all_features[2227] , \all_features[2228] ,
    \all_features[2229] , \all_features[2230] , \all_features[2231] ,
    \all_features[2232] , \all_features[2233] , \all_features[2234] ,
    \all_features[2235] , \all_features[2236] , \all_features[2237] ,
    \all_features[2238] , \all_features[2239] , \all_features[2240] ,
    \all_features[2241] , \all_features[2242] , \all_features[2243] ,
    \all_features[2244] , \all_features[2245] , \all_features[2246] ,
    \all_features[2247] , \all_features[2248] , \all_features[2249] ,
    \all_features[2250] , \all_features[2251] , \all_features[2252] ,
    \all_features[2253] , \all_features[2254] , \all_features[2255] ,
    \all_features[2256] , \all_features[2257] , \all_features[2258] ,
    \all_features[2259] , \all_features[2260] , \all_features[2261] ,
    \all_features[2262] , \all_features[2263] , \all_features[2264] ,
    \all_features[2265] , \all_features[2266] , \all_features[2267] ,
    \all_features[2268] , \all_features[2269] , \all_features[2270] ,
    \all_features[2271] , \all_features[2272] , \all_features[2273] ,
    \all_features[2274] , \all_features[2275] , \all_features[2276] ,
    \all_features[2277] , \all_features[2278] , \all_features[2279] ,
    \all_features[2280] , \all_features[2281] , \all_features[2282] ,
    \all_features[2283] , \all_features[2284] , \all_features[2285] ,
    \all_features[2286] , \all_features[2287] , \all_features[2288] ,
    \all_features[2289] , \all_features[2290] , \all_features[2291] ,
    \all_features[2292] , \all_features[2293] , \all_features[2294] ,
    \all_features[2295] , \all_features[2296] , \all_features[2297] ,
    \all_features[2298] , \all_features[2299] , \all_features[2300] ,
    \all_features[2301] , \all_features[2302] , \all_features[2303] ,
    \all_features[2304] , \all_features[2305] , \all_features[2306] ,
    \all_features[2307] , \all_features[2308] , \all_features[2309] ,
    \all_features[2310] , \all_features[2311] , \all_features[2312] ,
    \all_features[2313] , \all_features[2314] , \all_features[2315] ,
    \all_features[2316] , \all_features[2317] , \all_features[2318] ,
    \all_features[2319] , \all_features[2320] , \all_features[2321] ,
    \all_features[2322] , \all_features[2323] , \all_features[2324] ,
    \all_features[2325] , \all_features[2326] , \all_features[2327] ,
    \all_features[2328] , \all_features[2329] , \all_features[2330] ,
    \all_features[2331] , \all_features[2332] , \all_features[2333] ,
    \all_features[2334] , \all_features[2335] , \all_features[2336] ,
    \all_features[2337] , \all_features[2338] , \all_features[2339] ,
    \all_features[2340] , \all_features[2341] , \all_features[2342] ,
    \all_features[2343] , \all_features[2344] , \all_features[2345] ,
    \all_features[2346] , \all_features[2347] , \all_features[2348] ,
    \all_features[2349] , \all_features[2350] , \all_features[2351] ,
    \all_features[2352] , \all_features[2353] , \all_features[2354] ,
    \all_features[2355] , \all_features[2356] , \all_features[2357] ,
    \all_features[2358] , \all_features[2359] , \all_features[2360] ,
    \all_features[2361] , \all_features[2362] , \all_features[2363] ,
    \all_features[2364] , \all_features[2365] , \all_features[2366] ,
    \all_features[2367] , \all_features[2368] , \all_features[2369] ,
    \all_features[2370] , \all_features[2371] , \all_features[2372] ,
    \all_features[2373] , \all_features[2374] , \all_features[2375] ,
    \all_features[2376] , \all_features[2377] , \all_features[2378] ,
    \all_features[2379] , \all_features[2380] , \all_features[2381] ,
    \all_features[2382] , \all_features[2383] , \all_features[2384] ,
    \all_features[2385] , \all_features[2386] , \all_features[2387] ,
    \all_features[2388] , \all_features[2389] , \all_features[2390] ,
    \all_features[2391] , \all_features[2392] , \all_features[2393] ,
    \all_features[2394] , \all_features[2395] , \all_features[2396] ,
    \all_features[2397] , \all_features[2398] , \all_features[2399] ,
    \all_features[2400] , \all_features[2401] , \all_features[2402] ,
    \all_features[2403] , \all_features[2404] , \all_features[2405] ,
    \all_features[2406] , \all_features[2407] , \all_features[2408] ,
    \all_features[2409] , \all_features[2410] , \all_features[2411] ,
    \all_features[2412] , \all_features[2413] , \all_features[2414] ,
    \all_features[2415] , \all_features[2416] , \all_features[2417] ,
    \all_features[2418] , \all_features[2419] , \all_features[2420] ,
    \all_features[2421] , \all_features[2422] , \all_features[2423] ,
    \all_features[2424] , \all_features[2425] , \all_features[2426] ,
    \all_features[2427] , \all_features[2428] , \all_features[2429] ,
    \all_features[2430] , \all_features[2431] , \all_features[2432] ,
    \all_features[2433] , \all_features[2434] , \all_features[2435] ,
    \all_features[2436] , \all_features[2437] , \all_features[2438] ,
    \all_features[2439] , \all_features[2440] , \all_features[2441] ,
    \all_features[2442] , \all_features[2443] , \all_features[2444] ,
    \all_features[2445] , \all_features[2446] , \all_features[2447] ,
    \all_features[2448] , \all_features[2449] , \all_features[2450] ,
    \all_features[2451] , \all_features[2452] , \all_features[2453] ,
    \all_features[2454] , \all_features[2455] , \all_features[2456] ,
    \all_features[2457] , \all_features[2458] , \all_features[2459] ,
    \all_features[2460] , \all_features[2461] , \all_features[2462] ,
    \all_features[2463] , \all_features[2464] , \all_features[2465] ,
    \all_features[2466] , \all_features[2467] , \all_features[2468] ,
    \all_features[2469] , \all_features[2470] , \all_features[2471] ,
    \all_features[2472] , \all_features[2473] , \all_features[2474] ,
    \all_features[2475] , \all_features[2476] , \all_features[2477] ,
    \all_features[2478] , \all_features[2479] , \all_features[2480] ,
    \all_features[2481] , \all_features[2482] , \all_features[2483] ,
    \all_features[2484] , \all_features[2485] , \all_features[2486] ,
    \all_features[2487] , \all_features[2488] , \all_features[2489] ,
    \all_features[2490] , \all_features[2491] , \all_features[2492] ,
    \all_features[2493] , \all_features[2494] , \all_features[2495] ,
    \all_features[2496] , \all_features[2497] , \all_features[2498] ,
    \all_features[2499] , \all_features[2500] , \all_features[2501] ,
    \all_features[2502] , \all_features[2503] , \all_features[2504] ,
    \all_features[2505] , \all_features[2506] , \all_features[2507] ,
    \all_features[2508] , \all_features[2509] , \all_features[2510] ,
    \all_features[2511] , \all_features[2512] , \all_features[2513] ,
    \all_features[2514] , \all_features[2515] , \all_features[2516] ,
    \all_features[2517] , \all_features[2518] , \all_features[2519] ,
    \all_features[2520] , \all_features[2521] , \all_features[2522] ,
    \all_features[2523] , \all_features[2524] , \all_features[2525] ,
    \all_features[2526] , \all_features[2527] , \all_features[2528] ,
    \all_features[2529] , \all_features[2530] , \all_features[2531] ,
    \all_features[2532] , \all_features[2533] , \all_features[2534] ,
    \all_features[2535] , \all_features[2536] , \all_features[2537] ,
    \all_features[2538] , \all_features[2539] , \all_features[2540] ,
    \all_features[2541] , \all_features[2542] , \all_features[2543] ,
    \all_features[2544] , \all_features[2545] , \all_features[2546] ,
    \all_features[2547] , \all_features[2548] , \all_features[2549] ,
    \all_features[2550] , \all_features[2551] , \all_features[2552] ,
    \all_features[2553] , \all_features[2554] , \all_features[2555] ,
    \all_features[2556] , \all_features[2557] , \all_features[2558] ,
    \all_features[2559] , \all_features[2560] , \all_features[2561] ,
    \all_features[2562] , \all_features[2563] , \all_features[2564] ,
    \all_features[2565] , \all_features[2566] , \all_features[2567] ,
    \all_features[2568] , \all_features[2569] , \all_features[2570] ,
    \all_features[2571] , \all_features[2572] , \all_features[2573] ,
    \all_features[2574] , \all_features[2575] , \all_features[2576] ,
    \all_features[2577] , \all_features[2578] , \all_features[2579] ,
    \all_features[2580] , \all_features[2581] , \all_features[2582] ,
    \all_features[2583] , \all_features[2584] , \all_features[2585] ,
    \all_features[2586] , \all_features[2587] , \all_features[2588] ,
    \all_features[2589] , \all_features[2590] , \all_features[2591] ,
    \all_features[2592] , \all_features[2593] , \all_features[2594] ,
    \all_features[2595] , \all_features[2596] , \all_features[2597] ,
    \all_features[2598] , \all_features[2599] , \all_features[2600] ,
    \all_features[2601] , \all_features[2602] , \all_features[2603] ,
    \all_features[2604] , \all_features[2605] , \all_features[2606] ,
    \all_features[2607] , \all_features[2608] , \all_features[2609] ,
    \all_features[2610] , \all_features[2611] , \all_features[2612] ,
    \all_features[2613] , \all_features[2614] , \all_features[2615] ,
    \all_features[2616] , \all_features[2617] , \all_features[2618] ,
    \all_features[2619] , \all_features[2620] , \all_features[2621] ,
    \all_features[2622] , \all_features[2623] , \all_features[2624] ,
    \all_features[2625] , \all_features[2626] , \all_features[2627] ,
    \all_features[2628] , \all_features[2629] , \all_features[2630] ,
    \all_features[2631] , \all_features[2632] , \all_features[2633] ,
    \all_features[2634] , \all_features[2635] , \all_features[2636] ,
    \all_features[2637] , \all_features[2638] , \all_features[2639] ,
    \all_features[2640] , \all_features[2641] , \all_features[2642] ,
    \all_features[2643] , \all_features[2644] , \all_features[2645] ,
    \all_features[2646] , \all_features[2647] , \all_features[2648] ,
    \all_features[2649] , \all_features[2650] , \all_features[2651] ,
    \all_features[2652] , \all_features[2653] , \all_features[2654] ,
    \all_features[2655] , \all_features[2656] , \all_features[2657] ,
    \all_features[2658] , \all_features[2659] , \all_features[2660] ,
    \all_features[2661] , \all_features[2662] , \all_features[2663] ,
    \all_features[2664] , \all_features[2665] , \all_features[2666] ,
    \all_features[2667] , \all_features[2668] , \all_features[2669] ,
    \all_features[2670] , \all_features[2671] , \all_features[2672] ,
    \all_features[2673] , \all_features[2674] , \all_features[2675] ,
    \all_features[2676] , \all_features[2677] , \all_features[2678] ,
    \all_features[2679] , \all_features[2680] , \all_features[2681] ,
    \all_features[2682] , \all_features[2683] , \all_features[2684] ,
    \all_features[2685] , \all_features[2686] , \all_features[2687] ,
    \all_features[2688] , \all_features[2689] , \all_features[2690] ,
    \all_features[2691] , \all_features[2692] , \all_features[2693] ,
    \all_features[2694] , \all_features[2695] , \all_features[2696] ,
    \all_features[2697] , \all_features[2698] , \all_features[2699] ,
    \all_features[2700] , \all_features[2701] , \all_features[2702] ,
    \all_features[2703] , \all_features[2704] , \all_features[2705] ,
    \all_features[2706] , \all_features[2707] , \all_features[2708] ,
    \all_features[2709] , \all_features[2710] , \all_features[2711] ,
    \all_features[2712] , \all_features[2713] , \all_features[2714] ,
    \all_features[2715] , \all_features[2716] , \all_features[2717] ,
    \all_features[2718] , \all_features[2719] , \all_features[2720] ,
    \all_features[2721] , \all_features[2722] , \all_features[2723] ,
    \all_features[2724] , \all_features[2725] , \all_features[2726] ,
    \all_features[2727] , \all_features[2728] , \all_features[2729] ,
    \all_features[2730] , \all_features[2731] , \all_features[2732] ,
    \all_features[2733] , \all_features[2734] , \all_features[2735] ,
    \all_features[2736] , \all_features[2737] , \all_features[2738] ,
    \all_features[2739] , \all_features[2740] , \all_features[2741] ,
    \all_features[2742] , \all_features[2743] , \all_features[2744] ,
    \all_features[2745] , \all_features[2746] , \all_features[2747] ,
    \all_features[2748] , \all_features[2749] , \all_features[2750] ,
    \all_features[2751] , \all_features[2752] , \all_features[2753] ,
    \all_features[2754] , \all_features[2755] , \all_features[2756] ,
    \all_features[2757] , \all_features[2758] , \all_features[2759] ,
    \all_features[2760] , \all_features[2761] , \all_features[2762] ,
    \all_features[2763] , \all_features[2764] , \all_features[2765] ,
    \all_features[2766] , \all_features[2767] , \all_features[2768] ,
    \all_features[2769] , \all_features[2770] , \all_features[2771] ,
    \all_features[2772] , \all_features[2773] , \all_features[2774] ,
    \all_features[2775] , \all_features[2776] , \all_features[2777] ,
    \all_features[2778] , \all_features[2779] , \all_features[2780] ,
    \all_features[2781] , \all_features[2782] , \all_features[2783] ,
    \all_features[2784] , \all_features[2785] , \all_features[2786] ,
    \all_features[2787] , \all_features[2788] , \all_features[2789] ,
    \all_features[2790] , \all_features[2791] , \all_features[2792] ,
    \all_features[2793] , \all_features[2794] , \all_features[2795] ,
    \all_features[2796] , \all_features[2797] , \all_features[2798] ,
    \all_features[2799] , \all_features[2800] , \all_features[2801] ,
    \all_features[2802] , \all_features[2803] , \all_features[2804] ,
    \all_features[2805] , \all_features[2806] , \all_features[2807] ,
    \all_features[2808] , \all_features[2809] , \all_features[2810] ,
    \all_features[2811] , \all_features[2812] , \all_features[2813] ,
    \all_features[2814] , \all_features[2815] , \all_features[2816] ,
    \all_features[2817] , \all_features[2818] , \all_features[2819] ,
    \all_features[2820] , \all_features[2821] , \all_features[2822] ,
    \all_features[2823] , \all_features[2824] , \all_features[2825] ,
    \all_features[2826] , \all_features[2827] , \all_features[2828] ,
    \all_features[2829] , \all_features[2830] , \all_features[2831] ,
    \all_features[2832] , \all_features[2833] , \all_features[2834] ,
    \all_features[2835] , \all_features[2836] , \all_features[2837] ,
    \all_features[2838] , \all_features[2839] , \all_features[2840] ,
    \all_features[2841] , \all_features[2842] , \all_features[2843] ,
    \all_features[2844] , \all_features[2845] , \all_features[2846] ,
    \all_features[2847] , \all_features[2848] , \all_features[2849] ,
    \all_features[2850] , \all_features[2851] , \all_features[2852] ,
    \all_features[2853] , \all_features[2854] , \all_features[2855] ,
    \all_features[2856] , \all_features[2857] , \all_features[2858] ,
    \all_features[2859] , \all_features[2860] , \all_features[2861] ,
    \all_features[2862] , \all_features[2863] , \all_features[2864] ,
    \all_features[2865] , \all_features[2866] , \all_features[2867] ,
    \all_features[2868] , \all_features[2869] , \all_features[2870] ,
    \all_features[2871] , \all_features[2872] , \all_features[2873] ,
    \all_features[2874] , \all_features[2875] , \all_features[2876] ,
    \all_features[2877] , \all_features[2878] , \all_features[2879] ,
    \all_features[2880] , \all_features[2881] , \all_features[2882] ,
    \all_features[2883] , \all_features[2884] , \all_features[2885] ,
    \all_features[2886] , \all_features[2887] , \all_features[2888] ,
    \all_features[2889] , \all_features[2890] , \all_features[2891] ,
    \all_features[2892] , \all_features[2893] , \all_features[2894] ,
    \all_features[2895] , \all_features[2896] , \all_features[2897] ,
    \all_features[2898] , \all_features[2899] , \all_features[2900] ,
    \all_features[2901] , \all_features[2902] , \all_features[2903] ,
    \all_features[2904] , \all_features[2905] , \all_features[2906] ,
    \all_features[2907] , \all_features[2908] , \all_features[2909] ,
    \all_features[2910] , \all_features[2911] , \all_features[2912] ,
    \all_features[2913] , \all_features[2914] , \all_features[2915] ,
    \all_features[2916] , \all_features[2917] , \all_features[2918] ,
    \all_features[2919] , \all_features[2920] , \all_features[2921] ,
    \all_features[2922] , \all_features[2923] , \all_features[2924] ,
    \all_features[2925] , \all_features[2926] , \all_features[2927] ,
    \all_features[2928] , \all_features[2929] , \all_features[2930] ,
    \all_features[2931] , \all_features[2932] , \all_features[2933] ,
    \all_features[2934] , \all_features[2935] , \all_features[2936] ,
    \all_features[2937] , \all_features[2938] , \all_features[2939] ,
    \all_features[2940] , \all_features[2941] , \all_features[2942] ,
    \all_features[2943] , \all_features[2944] , \all_features[2945] ,
    \all_features[2946] , \all_features[2947] , \all_features[2948] ,
    \all_features[2949] , \all_features[2950] , \all_features[2951] ,
    \all_features[2952] , \all_features[2953] , \all_features[2954] ,
    \all_features[2955] , \all_features[2956] , \all_features[2957] ,
    \all_features[2958] , \all_features[2959] , \all_features[2960] ,
    \all_features[2961] , \all_features[2962] , \all_features[2963] ,
    \all_features[2964] , \all_features[2965] , \all_features[2966] ,
    \all_features[2967] , \all_features[2968] , \all_features[2969] ,
    \all_features[2970] , \all_features[2971] , \all_features[2972] ,
    \all_features[2973] , \all_features[2974] , \all_features[2975] ,
    \all_features[2976] , \all_features[2977] , \all_features[2978] ,
    \all_features[2979] , \all_features[2980] , \all_features[2981] ,
    \all_features[2982] , \all_features[2983] , \all_features[2984] ,
    \all_features[2985] , \all_features[2986] , \all_features[2987] ,
    \all_features[2988] , \all_features[2989] , \all_features[2990] ,
    \all_features[2991] , \all_features[2992] , \all_features[2993] ,
    \all_features[2994] , \all_features[2995] , \all_features[2996] ,
    \all_features[2997] , \all_features[2998] , \all_features[2999] ,
    \all_features[3000] , \all_features[3001] , \all_features[3002] ,
    \all_features[3003] , \all_features[3004] , \all_features[3005] ,
    \all_features[3006] , \all_features[3007] , \all_features[3008] ,
    \all_features[3009] , \all_features[3010] , \all_features[3011] ,
    \all_features[3012] , \all_features[3013] , \all_features[3014] ,
    \all_features[3015] , \all_features[3016] , \all_features[3017] ,
    \all_features[3018] , \all_features[3019] , \all_features[3020] ,
    \all_features[3021] , \all_features[3022] , \all_features[3023] ,
    \all_features[3024] , \all_features[3025] , \all_features[3026] ,
    \all_features[3027] , \all_features[3028] , \all_features[3029] ,
    \all_features[3030] , \all_features[3031] , \all_features[3032] ,
    \all_features[3033] , \all_features[3034] , \all_features[3035] ,
    \all_features[3036] , \all_features[3037] , \all_features[3038] ,
    \all_features[3039] , \all_features[3040] , \all_features[3041] ,
    \all_features[3042] , \all_features[3043] , \all_features[3044] ,
    \all_features[3045] , \all_features[3046] , \all_features[3047] ,
    \all_features[3048] , \all_features[3049] , \all_features[3050] ,
    \all_features[3051] , \all_features[3052] , \all_features[3053] ,
    \all_features[3054] , \all_features[3055] , \all_features[3056] ,
    \all_features[3057] , \all_features[3058] , \all_features[3059] ,
    \all_features[3060] , \all_features[3061] , \all_features[3062] ,
    \all_features[3063] , \all_features[3064] , \all_features[3065] ,
    \all_features[3066] , \all_features[3067] , \all_features[3068] ,
    \all_features[3069] , \all_features[3070] , \all_features[3071] ,
    \all_features[3072] , \all_features[3073] , \all_features[3074] ,
    \all_features[3075] , \all_features[3076] , \all_features[3077] ,
    \all_features[3078] , \all_features[3079] , \all_features[3080] ,
    \all_features[3081] , \all_features[3082] , \all_features[3083] ,
    \all_features[3084] , \all_features[3085] , \all_features[3086] ,
    \all_features[3087] , \all_features[3088] , \all_features[3089] ,
    \all_features[3090] , \all_features[3091] , \all_features[3092] ,
    \all_features[3093] , \all_features[3094] , \all_features[3095] ,
    \all_features[3096] , \all_features[3097] , \all_features[3098] ,
    \all_features[3099] , \all_features[3100] , \all_features[3101] ,
    \all_features[3102] , \all_features[3103] , \all_features[3104] ,
    \all_features[3105] , \all_features[3106] , \all_features[3107] ,
    \all_features[3108] , \all_features[3109] , \all_features[3110] ,
    \all_features[3111] , \all_features[3112] , \all_features[3113] ,
    \all_features[3114] , \all_features[3115] , \all_features[3116] ,
    \all_features[3117] , \all_features[3118] , \all_features[3119] ,
    \all_features[3120] , \all_features[3121] , \all_features[3122] ,
    \all_features[3123] , \all_features[3124] , \all_features[3125] ,
    \all_features[3126] , \all_features[3127] , \all_features[3128] ,
    \all_features[3129] , \all_features[3130] , \all_features[3131] ,
    \all_features[3132] , \all_features[3133] , \all_features[3134] ,
    \all_features[3135] , \all_features[3136] , \all_features[3137] ,
    \all_features[3138] , \all_features[3139] , \all_features[3140] ,
    \all_features[3141] , \all_features[3142] , \all_features[3143] ,
    \all_features[3144] , \all_features[3145] , \all_features[3146] ,
    \all_features[3147] , \all_features[3148] , \all_features[3149] ,
    \all_features[3150] , \all_features[3151] , \all_features[3152] ,
    \all_features[3153] , \all_features[3154] , \all_features[3155] ,
    \all_features[3156] , \all_features[3157] , \all_features[3158] ,
    \all_features[3159] , \all_features[3160] , \all_features[3161] ,
    \all_features[3162] , \all_features[3163] , \all_features[3164] ,
    \all_features[3165] , \all_features[3166] , \all_features[3167] ,
    \all_features[3168] , \all_features[3169] , \all_features[3170] ,
    \all_features[3171] , \all_features[3172] , \all_features[3173] ,
    \all_features[3174] , \all_features[3175] , \all_features[3176] ,
    \all_features[3177] , \all_features[3178] , \all_features[3179] ,
    \all_features[3180] , \all_features[3181] , \all_features[3182] ,
    \all_features[3183] , \all_features[3184] , \all_features[3185] ,
    \all_features[3186] , \all_features[3187] , \all_features[3188] ,
    \all_features[3189] , \all_features[3190] , \all_features[3191] ,
    \all_features[3192] , \all_features[3193] , \all_features[3194] ,
    \all_features[3195] , \all_features[3196] , \all_features[3197] ,
    \all_features[3198] , \all_features[3199] , \all_features[3200] ,
    \all_features[3201] , \all_features[3202] , \all_features[3203] ,
    \all_features[3204] , \all_features[3205] , \all_features[3206] ,
    \all_features[3207] , \all_features[3208] , \all_features[3209] ,
    \all_features[3210] , \all_features[3211] , \all_features[3212] ,
    \all_features[3213] , \all_features[3214] , \all_features[3215] ,
    \all_features[3216] , \all_features[3217] , \all_features[3218] ,
    \all_features[3219] , \all_features[3220] , \all_features[3221] ,
    \all_features[3222] , \all_features[3223] , \all_features[3224] ,
    \all_features[3225] , \all_features[3226] , \all_features[3227] ,
    \all_features[3228] , \all_features[3229] , \all_features[3230] ,
    \all_features[3231] , \all_features[3232] , \all_features[3233] ,
    \all_features[3234] , \all_features[3235] , \all_features[3236] ,
    \all_features[3237] , \all_features[3238] , \all_features[3239] ,
    \all_features[3240] , \all_features[3241] , \all_features[3242] ,
    \all_features[3243] , \all_features[3244] , \all_features[3245] ,
    \all_features[3246] , \all_features[3247] , \all_features[3248] ,
    \all_features[3249] , \all_features[3250] , \all_features[3251] ,
    \all_features[3252] , \all_features[3253] , \all_features[3254] ,
    \all_features[3255] , \all_features[3256] , \all_features[3257] ,
    \all_features[3258] , \all_features[3259] , \all_features[3260] ,
    \all_features[3261] , \all_features[3262] , \all_features[3263] ,
    \all_features[3264] , \all_features[3265] , \all_features[3266] ,
    \all_features[3267] , \all_features[3268] , \all_features[3269] ,
    \all_features[3270] , \all_features[3271] , \all_features[3272] ,
    \all_features[3273] , \all_features[3274] , \all_features[3275] ,
    \all_features[3276] , \all_features[3277] , \all_features[3278] ,
    \all_features[3279] , \all_features[3280] , \all_features[3281] ,
    \all_features[3282] , \all_features[3283] , \all_features[3284] ,
    \all_features[3285] , \all_features[3286] , \all_features[3287] ,
    \all_features[3288] , \all_features[3289] , \all_features[3290] ,
    \all_features[3291] , \all_features[3292] , \all_features[3293] ,
    \all_features[3294] , \all_features[3295] , \all_features[3296] ,
    \all_features[3297] , \all_features[3298] , \all_features[3299] ,
    \all_features[3300] , \all_features[3301] , \all_features[3302] ,
    \all_features[3303] , \all_features[3304] , \all_features[3305] ,
    \all_features[3306] , \all_features[3307] , \all_features[3308] ,
    \all_features[3309] , \all_features[3310] , \all_features[3311] ,
    \all_features[3312] , \all_features[3313] , \all_features[3314] ,
    \all_features[3315] , \all_features[3316] , \all_features[3317] ,
    \all_features[3318] , \all_features[3319] , \all_features[3320] ,
    \all_features[3321] , \all_features[3322] , \all_features[3323] ,
    \all_features[3324] , \all_features[3325] , \all_features[3326] ,
    \all_features[3327] , \all_features[3328] , \all_features[3329] ,
    \all_features[3330] , \all_features[3331] , \all_features[3332] ,
    \all_features[3333] , \all_features[3334] , \all_features[3335] ,
    \all_features[3336] , \all_features[3337] , \all_features[3338] ,
    \all_features[3339] , \all_features[3340] , \all_features[3341] ,
    \all_features[3342] , \all_features[3343] , \all_features[3344] ,
    \all_features[3345] , \all_features[3346] , \all_features[3347] ,
    \all_features[3348] , \all_features[3349] , \all_features[3350] ,
    \all_features[3351] , \all_features[3352] , \all_features[3353] ,
    \all_features[3354] , \all_features[3355] , \all_features[3356] ,
    \all_features[3357] , \all_features[3358] , \all_features[3359] ,
    \all_features[3360] , \all_features[3361] , \all_features[3362] ,
    \all_features[3363] , \all_features[3364] , \all_features[3365] ,
    \all_features[3366] , \all_features[3367] , \all_features[3368] ,
    \all_features[3369] , \all_features[3370] , \all_features[3371] ,
    \all_features[3372] , \all_features[3373] , \all_features[3374] ,
    \all_features[3375] , \all_features[3376] , \all_features[3377] ,
    \all_features[3378] , \all_features[3379] , \all_features[3380] ,
    \all_features[3381] , \all_features[3382] , \all_features[3383] ,
    \all_features[3384] , \all_features[3385] , \all_features[3386] ,
    \all_features[3387] , \all_features[3388] , \all_features[3389] ,
    \all_features[3390] , \all_features[3391] , \all_features[3392] ,
    \all_features[3393] , \all_features[3394] , \all_features[3395] ,
    \all_features[3396] , \all_features[3397] , \all_features[3398] ,
    \all_features[3399] , \all_features[3400] , \all_features[3401] ,
    \all_features[3402] , \all_features[3403] , \all_features[3404] ,
    \all_features[3405] , \all_features[3406] , \all_features[3407] ,
    \all_features[3408] , \all_features[3409] , \all_features[3410] ,
    \all_features[3411] , \all_features[3412] , \all_features[3413] ,
    \all_features[3414] , \all_features[3415] , \all_features[3416] ,
    \all_features[3417] , \all_features[3418] , \all_features[3419] ,
    \all_features[3420] , \all_features[3421] , \all_features[3422] ,
    \all_features[3423] , \all_features[3424] , \all_features[3425] ,
    \all_features[3426] , \all_features[3427] , \all_features[3428] ,
    \all_features[3429] , \all_features[3430] , \all_features[3431] ,
    \all_features[3432] , \all_features[3433] , \all_features[3434] ,
    \all_features[3435] , \all_features[3436] , \all_features[3437] ,
    \all_features[3438] , \all_features[3439] , \all_features[3440] ,
    \all_features[3441] , \all_features[3442] , \all_features[3443] ,
    \all_features[3444] , \all_features[3445] , \all_features[3446] ,
    \all_features[3447] , \all_features[3448] , \all_features[3449] ,
    \all_features[3450] , \all_features[3451] , \all_features[3452] ,
    \all_features[3453] , \all_features[3454] , \all_features[3455] ,
    \all_features[3456] , \all_features[3457] , \all_features[3458] ,
    \all_features[3459] , \all_features[3460] , \all_features[3461] ,
    \all_features[3462] , \all_features[3463] , \all_features[3464] ,
    \all_features[3465] , \all_features[3466] , \all_features[3467] ,
    \all_features[3468] , \all_features[3469] , \all_features[3470] ,
    \all_features[3471] , \all_features[3472] , \all_features[3473] ,
    \all_features[3474] , \all_features[3475] , \all_features[3476] ,
    \all_features[3477] , \all_features[3478] , \all_features[3479] ,
    \all_features[3480] , \all_features[3481] , \all_features[3482] ,
    \all_features[3483] , \all_features[3484] , \all_features[3485] ,
    \all_features[3486] , \all_features[3487] , \all_features[3488] ,
    \all_features[3489] , \all_features[3490] , \all_features[3491] ,
    \all_features[3492] , \all_features[3493] , \all_features[3494] ,
    \all_features[3495] , \all_features[3496] , \all_features[3497] ,
    \all_features[3498] , \all_features[3499] , \all_features[3500] ,
    \all_features[3501] , \all_features[3502] , \all_features[3503] ,
    \all_features[3504] , \all_features[3505] , \all_features[3506] ,
    \all_features[3507] , \all_features[3508] , \all_features[3509] ,
    \all_features[3510] , \all_features[3511] , \all_features[3512] ,
    \all_features[3513] , \all_features[3514] , \all_features[3515] ,
    \all_features[3516] , \all_features[3517] , \all_features[3518] ,
    \all_features[3519] , \all_features[3520] , \all_features[3521] ,
    \all_features[3522] , \all_features[3523] , \all_features[3524] ,
    \all_features[3525] , \all_features[3526] , \all_features[3527] ,
    \all_features[3528] , \all_features[3529] , \all_features[3530] ,
    \all_features[3531] , \all_features[3532] , \all_features[3533] ,
    \all_features[3534] , \all_features[3535] , \all_features[3536] ,
    \all_features[3537] , \all_features[3538] , \all_features[3539] ,
    \all_features[3540] , \all_features[3541] , \all_features[3542] ,
    \all_features[3543] , \all_features[3544] , \all_features[3545] ,
    \all_features[3546] , \all_features[3547] , \all_features[3548] ,
    \all_features[3549] , \all_features[3550] , \all_features[3551] ,
    \all_features[3552] , \all_features[3553] , \all_features[3554] ,
    \all_features[3555] , \all_features[3556] , \all_features[3557] ,
    \all_features[3558] , \all_features[3559] , \all_features[3560] ,
    \all_features[3561] , \all_features[3562] , \all_features[3563] ,
    \all_features[3564] , \all_features[3565] , \all_features[3566] ,
    \all_features[3567] , \all_features[3568] , \all_features[3569] ,
    \all_features[3570] , \all_features[3571] , \all_features[3572] ,
    \all_features[3573] , \all_features[3574] , \all_features[3575] ,
    \all_features[3576] , \all_features[3577] , \all_features[3578] ,
    \all_features[3579] , \all_features[3580] , \all_features[3581] ,
    \all_features[3582] , \all_features[3583] , \all_features[3584] ,
    \all_features[3585] , \all_features[3586] , \all_features[3587] ,
    \all_features[3588] , \all_features[3589] , \all_features[3590] ,
    \all_features[3591] , \all_features[3592] , \all_features[3593] ,
    \all_features[3594] , \all_features[3595] , \all_features[3596] ,
    \all_features[3597] , \all_features[3598] , \all_features[3599] ,
    \all_features[3600] , \all_features[3601] , \all_features[3602] ,
    \all_features[3603] , \all_features[3604] , \all_features[3605] ,
    \all_features[3606] , \all_features[3607] , \all_features[3608] ,
    \all_features[3609] , \all_features[3610] , \all_features[3611] ,
    \all_features[3612] , \all_features[3613] , \all_features[3614] ,
    \all_features[3615] , \all_features[3616] , \all_features[3617] ,
    \all_features[3618] , \all_features[3619] , \all_features[3620] ,
    \all_features[3621] , \all_features[3622] , \all_features[3623] ,
    \all_features[3624] , \all_features[3625] , \all_features[3626] ,
    \all_features[3627] , \all_features[3628] , \all_features[3629] ,
    \all_features[3630] , \all_features[3631] , \all_features[3632] ,
    \all_features[3633] , \all_features[3634] , \all_features[3635] ,
    \all_features[3636] , \all_features[3637] , \all_features[3638] ,
    \all_features[3639] , \all_features[3640] , \all_features[3641] ,
    \all_features[3642] , \all_features[3643] , \all_features[3644] ,
    \all_features[3645] , \all_features[3646] , \all_features[3647] ,
    \all_features[3648] , \all_features[3649] , \all_features[3650] ,
    \all_features[3651] , \all_features[3652] , \all_features[3653] ,
    \all_features[3654] , \all_features[3655] , \all_features[3656] ,
    \all_features[3657] , \all_features[3658] , \all_features[3659] ,
    \all_features[3660] , \all_features[3661] , \all_features[3662] ,
    \all_features[3663] , \all_features[3664] , \all_features[3665] ,
    \all_features[3666] , \all_features[3667] , \all_features[3668] ,
    \all_features[3669] , \all_features[3670] , \all_features[3671] ,
    \all_features[3672] , \all_features[3673] , \all_features[3674] ,
    \all_features[3675] , \all_features[3676] , \all_features[3677] ,
    \all_features[3678] , \all_features[3679] , \all_features[3680] ,
    \all_features[3681] , \all_features[3682] , \all_features[3683] ,
    \all_features[3684] , \all_features[3685] , \all_features[3686] ,
    \all_features[3687] , \all_features[3688] , \all_features[3689] ,
    \all_features[3690] , \all_features[3691] , \all_features[3692] ,
    \all_features[3693] , \all_features[3694] , \all_features[3695] ,
    \all_features[3696] , \all_features[3697] , \all_features[3698] ,
    \all_features[3699] , \all_features[3700] , \all_features[3701] ,
    \all_features[3702] , \all_features[3703] , \all_features[3704] ,
    \all_features[3705] , \all_features[3706] , \all_features[3707] ,
    \all_features[3708] , \all_features[3709] , \all_features[3710] ,
    \all_features[3711] , \all_features[3712] , \all_features[3713] ,
    \all_features[3714] , \all_features[3715] , \all_features[3716] ,
    \all_features[3717] , \all_features[3718] , \all_features[3719] ,
    \all_features[3720] , \all_features[3721] , \all_features[3722] ,
    \all_features[3723] , \all_features[3724] , \all_features[3725] ,
    \all_features[3726] , \all_features[3727] , \all_features[3728] ,
    \all_features[3729] , \all_features[3730] , \all_features[3731] ,
    \all_features[3732] , \all_features[3733] , \all_features[3734] ,
    \all_features[3735] , \all_features[3736] , \all_features[3737] ,
    \all_features[3738] , \all_features[3739] , \all_features[3740] ,
    \all_features[3741] , \all_features[3742] , \all_features[3743] ,
    \all_features[3744] , \all_features[3745] , \all_features[3746] ,
    \all_features[3747] , \all_features[3748] , \all_features[3749] ,
    \all_features[3750] , \all_features[3751] , \all_features[3752] ,
    \all_features[3753] , \all_features[3754] , \all_features[3755] ,
    \all_features[3756] , \all_features[3757] , \all_features[3758] ,
    \all_features[3759] , \all_features[3760] , \all_features[3761] ,
    \all_features[3762] , \all_features[3763] , \all_features[3764] ,
    \all_features[3765] , \all_features[3766] , \all_features[3767] ,
    \all_features[3768] , \all_features[3769] , \all_features[3770] ,
    \all_features[3771] , \all_features[3772] , \all_features[3773] ,
    \all_features[3774] , \all_features[3775] , \all_features[3776] ,
    \all_features[3777] , \all_features[3778] , \all_features[3779] ,
    \all_features[3780] , \all_features[3781] , \all_features[3782] ,
    \all_features[3783] , \all_features[3784] , \all_features[3785] ,
    \all_features[3786] , \all_features[3787] , \all_features[3788] ,
    \all_features[3789] , \all_features[3790] , \all_features[3791] ,
    \all_features[3792] , \all_features[3793] , \all_features[3794] ,
    \all_features[3795] , \all_features[3796] , \all_features[3797] ,
    \all_features[3798] , \all_features[3799] , \all_features[3800] ,
    \all_features[3801] , \all_features[3802] , \all_features[3803] ,
    \all_features[3804] , \all_features[3805] , \all_features[3806] ,
    \all_features[3807] , \all_features[3808] , \all_features[3809] ,
    \all_features[3810] , \all_features[3811] , \all_features[3812] ,
    \all_features[3813] , \all_features[3814] , \all_features[3815] ,
    \all_features[3816] , \all_features[3817] , \all_features[3818] ,
    \all_features[3819] , \all_features[3820] , \all_features[3821] ,
    \all_features[3822] , \all_features[3823] , \all_features[3824] ,
    \all_features[3825] , \all_features[3826] , \all_features[3827] ,
    \all_features[3828] , \all_features[3829] , \all_features[3830] ,
    \all_features[3831] , \all_features[3832] , \all_features[3833] ,
    \all_features[3834] , \all_features[3835] , \all_features[3836] ,
    \all_features[3837] , \all_features[3838] , \all_features[3839] ,
    \all_features[3840] , \all_features[3841] , \all_features[3842] ,
    \all_features[3843] , \all_features[3844] , \all_features[3845] ,
    \all_features[3846] , \all_features[3847] , \all_features[3848] ,
    \all_features[3849] , \all_features[3850] , \all_features[3851] ,
    \all_features[3852] , \all_features[3853] , \all_features[3854] ,
    \all_features[3855] , \all_features[3856] , \all_features[3857] ,
    \all_features[3858] , \all_features[3859] , \all_features[3860] ,
    \all_features[3861] , \all_features[3862] , \all_features[3863] ,
    \all_features[3864] , \all_features[3865] , \all_features[3866] ,
    \all_features[3867] , \all_features[3868] , \all_features[3869] ,
    \all_features[3870] , \all_features[3871] , \all_features[3872] ,
    \all_features[3873] , \all_features[3874] , \all_features[3875] ,
    \all_features[3876] , \all_features[3877] , \all_features[3878] ,
    \all_features[3879] , \all_features[3880] , \all_features[3881] ,
    \all_features[3882] , \all_features[3883] , \all_features[3884] ,
    \all_features[3885] , \all_features[3886] , \all_features[3887] ,
    \all_features[3888] , \all_features[3889] , \all_features[3890] ,
    \all_features[3891] , \all_features[3892] , \all_features[3893] ,
    \all_features[3894] , \all_features[3895] , \all_features[3896] ,
    \all_features[3897] , \all_features[3898] , \all_features[3899] ,
    \all_features[3900] , \all_features[3901] , \all_features[3902] ,
    \all_features[3903] , \all_features[3904] , \all_features[3905] ,
    \all_features[3906] , \all_features[3907] , \all_features[3908] ,
    \all_features[3909] , \all_features[3910] , \all_features[3911] ,
    \all_features[3912] , \all_features[3913] , \all_features[3914] ,
    \all_features[3915] , \all_features[3916] , \all_features[3917] ,
    \all_features[3918] , \all_features[3919] , \all_features[3920] ,
    \all_features[3921] , \all_features[3922] , \all_features[3923] ,
    \all_features[3924] , \all_features[3925] , \all_features[3926] ,
    \all_features[3927] , \all_features[3928] , \all_features[3929] ,
    \all_features[3930] , \all_features[3931] , \all_features[3932] ,
    \all_features[3933] , \all_features[3934] , \all_features[3935] ,
    \all_features[3936] , \all_features[3937] , \all_features[3938] ,
    \all_features[3939] , \all_features[3940] , \all_features[3941] ,
    \all_features[3942] , \all_features[3943] , \all_features[3944] ,
    \all_features[3945] , \all_features[3946] , \all_features[3947] ,
    \all_features[3948] , \all_features[3949] , \all_features[3950] ,
    \all_features[3951] , \all_features[3952] , \all_features[3953] ,
    \all_features[3954] , \all_features[3955] , \all_features[3956] ,
    \all_features[3957] , \all_features[3958] , \all_features[3959] ,
    \all_features[3960] , \all_features[3961] , \all_features[3962] ,
    \all_features[3963] , \all_features[3964] , \all_features[3965] ,
    \all_features[3966] , \all_features[3967] , \all_features[3968] ,
    \all_features[3969] , \all_features[3970] , \all_features[3971] ,
    \all_features[3972] , \all_features[3973] , \all_features[3974] ,
    \all_features[3975] , \all_features[3976] , \all_features[3977] ,
    \all_features[3978] , \all_features[3979] , \all_features[3980] ,
    \all_features[3981] , \all_features[3982] , \all_features[3983] ,
    \all_features[3984] , \all_features[3985] , \all_features[3986] ,
    \all_features[3987] , \all_features[3988] , \all_features[3989] ,
    \all_features[3990] , \all_features[3991] , \all_features[3992] ,
    \all_features[3993] , \all_features[3994] , \all_features[3995] ,
    \all_features[3996] , \all_features[3997] , \all_features[3998] ,
    \all_features[3999] , \all_features[4000] , \all_features[4001] ,
    \all_features[4002] , \all_features[4003] , \all_features[4004] ,
    \all_features[4005] , \all_features[4006] , \all_features[4007] ,
    \all_features[4008] , \all_features[4009] , \all_features[4010] ,
    \all_features[4011] , \all_features[4012] , \all_features[4013] ,
    \all_features[4014] , \all_features[4015] , \all_features[4016] ,
    \all_features[4017] , \all_features[4018] , \all_features[4019] ,
    \all_features[4020] , \all_features[4021] , \all_features[4022] ,
    \all_features[4023] , \all_features[4024] , \all_features[4025] ,
    \all_features[4026] , \all_features[4027] , \all_features[4028] ,
    \all_features[4029] , \all_features[4030] , \all_features[4031] ,
    \all_features[4032] , \all_features[4033] , \all_features[4034] ,
    \all_features[4035] , \all_features[4036] , \all_features[4037] ,
    \all_features[4038] , \all_features[4039] , \all_features[4040] ,
    \all_features[4041] , \all_features[4042] , \all_features[4043] ,
    \all_features[4044] , \all_features[4045] , \all_features[4046] ,
    \all_features[4047] , \all_features[4048] , \all_features[4049] ,
    \all_features[4050] , \all_features[4051] , \all_features[4052] ,
    \all_features[4053] , \all_features[4054] , \all_features[4055] ,
    \all_features[4056] , \all_features[4057] , \all_features[4058] ,
    \all_features[4059] , \all_features[4060] , \all_features[4061] ,
    \all_features[4062] , \all_features[4063] , \all_features[4064] ,
    \all_features[4065] , \all_features[4066] , \all_features[4067] ,
    \all_features[4068] , \all_features[4069] , \all_features[4070] ,
    \all_features[4071] , \all_features[4072] , \all_features[4073] ,
    \all_features[4074] , \all_features[4075] , \all_features[4076] ,
    \all_features[4077] , \all_features[4078] , \all_features[4079] ,
    \all_features[4080] , \all_features[4081] , \all_features[4082] ,
    \all_features[4083] , \all_features[4084] , \all_features[4085] ,
    \all_features[4086] , \all_features[4087] , \all_features[4088] ,
    \all_features[4089] , \all_features[4090] , \all_features[4091] ,
    \all_features[4092] , \all_features[4093] , \all_features[4094] ,
    \all_features[4095] , \all_features[4096] , \all_features[4097] ,
    \all_features[4098] , \all_features[4099] , \all_features[4100] ,
    \all_features[4101] , \all_features[4102] , \all_features[4103] ,
    \all_features[4104] , \all_features[4105] , \all_features[4106] ,
    \all_features[4107] , \all_features[4108] , \all_features[4109] ,
    \all_features[4110] , \all_features[4111] , \all_features[4112] ,
    \all_features[4113] , \all_features[4114] , \all_features[4115] ,
    \all_features[4116] , \all_features[4117] , \all_features[4118] ,
    \all_features[4119] , \all_features[4120] , \all_features[4121] ,
    \all_features[4122] , \all_features[4123] , \all_features[4124] ,
    \all_features[4125] , \all_features[4126] , \all_features[4127] ,
    \all_features[4128] , \all_features[4129] , \all_features[4130] ,
    \all_features[4131] , \all_features[4132] , \all_features[4133] ,
    \all_features[4134] , \all_features[4135] , \all_features[4136] ,
    \all_features[4137] , \all_features[4138] , \all_features[4139] ,
    \all_features[4140] , \all_features[4141] , \all_features[4142] ,
    \all_features[4143] , \all_features[4144] , \all_features[4145] ,
    \all_features[4146] , \all_features[4147] , \all_features[4148] ,
    \all_features[4149] , \all_features[4150] , \all_features[4151] ,
    \all_features[4152] , \all_features[4153] , \all_features[4154] ,
    \all_features[4155] , \all_features[4156] , \all_features[4157] ,
    \all_features[4158] , \all_features[4159] , \all_features[4160] ,
    \all_features[4161] , \all_features[4162] , \all_features[4163] ,
    \all_features[4164] , \all_features[4165] , \all_features[4166] ,
    \all_features[4167] , \all_features[4168] , \all_features[4169] ,
    \all_features[4170] , \all_features[4171] , \all_features[4172] ,
    \all_features[4173] , \all_features[4174] , \all_features[4175] ,
    \all_features[4176] , \all_features[4177] , \all_features[4178] ,
    \all_features[4179] , \all_features[4180] , \all_features[4181] ,
    \all_features[4182] , \all_features[4183] , \all_features[4184] ,
    \all_features[4185] , \all_features[4186] , \all_features[4187] ,
    \all_features[4188] , \all_features[4189] , \all_features[4190] ,
    \all_features[4191] , \all_features[4192] , \all_features[4193] ,
    \all_features[4194] , \all_features[4195] , \all_features[4196] ,
    \all_features[4197] , \all_features[4198] , \all_features[4199] ,
    \all_features[4200] , \all_features[4201] , \all_features[4202] ,
    \all_features[4203] , \all_features[4204] , \all_features[4205] ,
    \all_features[4206] , \all_features[4207] , \all_features[4208] ,
    \all_features[4209] , \all_features[4210] , \all_features[4211] ,
    \all_features[4212] , \all_features[4213] , \all_features[4214] ,
    \all_features[4215] , \all_features[4216] , \all_features[4217] ,
    \all_features[4218] , \all_features[4219] , \all_features[4220] ,
    \all_features[4221] , \all_features[4222] , \all_features[4223] ,
    \all_features[4224] , \all_features[4225] , \all_features[4226] ,
    \all_features[4227] , \all_features[4228] , \all_features[4229] ,
    \all_features[4230] , \all_features[4231] , \all_features[4232] ,
    \all_features[4233] , \all_features[4234] , \all_features[4235] ,
    \all_features[4236] , \all_features[4237] , \all_features[4238] ,
    \all_features[4239] , \all_features[4240] , \all_features[4241] ,
    \all_features[4242] , \all_features[4243] , \all_features[4244] ,
    \all_features[4245] , \all_features[4246] , \all_features[4247] ,
    \all_features[4248] , \all_features[4249] , \all_features[4250] ,
    \all_features[4251] , \all_features[4252] , \all_features[4253] ,
    \all_features[4254] , \all_features[4255] , \all_features[4256] ,
    \all_features[4257] , \all_features[4258] , \all_features[4259] ,
    \all_features[4260] , \all_features[4261] , \all_features[4262] ,
    \all_features[4263] , \all_features[4264] , \all_features[4265] ,
    \all_features[4266] , \all_features[4267] , \all_features[4268] ,
    \all_features[4269] , \all_features[4270] , \all_features[4271] ,
    \all_features[4272] , \all_features[4273] , \all_features[4274] ,
    \all_features[4275] , \all_features[4276] , \all_features[4277] ,
    \all_features[4278] , \all_features[4279] , \all_features[4280] ,
    \all_features[4281] , \all_features[4282] , \all_features[4283] ,
    \all_features[4284] , \all_features[4285] , \all_features[4286] ,
    \all_features[4287] , \all_features[4288] , \all_features[4289] ,
    \all_features[4290] , \all_features[4291] , \all_features[4292] ,
    \all_features[4293] , \all_features[4294] , \all_features[4295] ,
    \all_features[4296] , \all_features[4297] , \all_features[4298] ,
    \all_features[4299] , \all_features[4300] , \all_features[4301] ,
    \all_features[4302] , \all_features[4303] , \all_features[4304] ,
    \all_features[4305] , \all_features[4306] , \all_features[4307] ,
    \all_features[4308] , \all_features[4309] , \all_features[4310] ,
    \all_features[4311] , \all_features[4312] , \all_features[4313] ,
    \all_features[4314] , \all_features[4315] , \all_features[4316] ,
    \all_features[4317] , \all_features[4318] , \all_features[4319] ,
    \all_features[4320] , \all_features[4321] , \all_features[4322] ,
    \all_features[4323] , \all_features[4324] , \all_features[4325] ,
    \all_features[4326] , \all_features[4327] , \all_features[4328] ,
    \all_features[4329] , \all_features[4330] , \all_features[4331] ,
    \all_features[4332] , \all_features[4333] , \all_features[4334] ,
    \all_features[4335] , \all_features[4336] , \all_features[4337] ,
    \all_features[4338] , \all_features[4339] , \all_features[4340] ,
    \all_features[4341] , \all_features[4342] , \all_features[4343] ,
    \all_features[4344] , \all_features[4345] , \all_features[4346] ,
    \all_features[4347] , \all_features[4348] , \all_features[4349] ,
    \all_features[4350] , \all_features[4351] , \all_features[4352] ,
    \all_features[4353] , \all_features[4354] , \all_features[4355] ,
    \all_features[4356] , \all_features[4357] , \all_features[4358] ,
    \all_features[4359] , \all_features[4360] , \all_features[4361] ,
    \all_features[4362] , \all_features[4363] , \all_features[4364] ,
    \all_features[4365] , \all_features[4366] , \all_features[4367] ,
    \all_features[4368] , \all_features[4369] , \all_features[4370] ,
    \all_features[4371] , \all_features[4372] , \all_features[4373] ,
    \all_features[4374] , \all_features[4375] , \all_features[4376] ,
    \all_features[4377] , \all_features[4378] , \all_features[4379] ,
    \all_features[4380] , \all_features[4381] , \all_features[4382] ,
    \all_features[4383] , \all_features[4384] , \all_features[4385] ,
    \all_features[4386] , \all_features[4387] , \all_features[4388] ,
    \all_features[4389] , \all_features[4390] , \all_features[4391] ,
    \all_features[4392] , \all_features[4393] , \all_features[4394] ,
    \all_features[4395] , \all_features[4396] , \all_features[4397] ,
    \all_features[4398] , \all_features[4399] , \all_features[4400] ,
    \all_features[4401] , \all_features[4402] , \all_features[4403] ,
    \all_features[4404] , \all_features[4405] , \all_features[4406] ,
    \all_features[4407] , \all_features[4408] , \all_features[4409] ,
    \all_features[4410] , \all_features[4411] , \all_features[4412] ,
    \all_features[4413] , \all_features[4414] , \all_features[4415] ,
    \all_features[4416] , \all_features[4417] , \all_features[4418] ,
    \all_features[4419] , \all_features[4420] , \all_features[4421] ,
    \all_features[4422] , \all_features[4423] , \all_features[4424] ,
    \all_features[4425] , \all_features[4426] , \all_features[4427] ,
    \all_features[4428] , \all_features[4429] , \all_features[4430] ,
    \all_features[4431] , \all_features[4432] , \all_features[4433] ,
    \all_features[4434] , \all_features[4435] , \all_features[4436] ,
    \all_features[4437] , \all_features[4438] , \all_features[4439] ,
    \all_features[4440] , \all_features[4441] , \all_features[4442] ,
    \all_features[4443] , \all_features[4444] , \all_features[4445] ,
    \all_features[4446] , \all_features[4447] , \all_features[4448] ,
    \all_features[4449] , \all_features[4450] , \all_features[4451] ,
    \all_features[4452] , \all_features[4453] , \all_features[4454] ,
    \all_features[4455] , \all_features[4456] , \all_features[4457] ,
    \all_features[4458] , \all_features[4459] , \all_features[4460] ,
    \all_features[4461] , \all_features[4462] , \all_features[4463] ,
    \all_features[4464] , \all_features[4465] , \all_features[4466] ,
    \all_features[4467] , \all_features[4468] , \all_features[4469] ,
    \all_features[4470] , \all_features[4471] , \all_features[4472] ,
    \all_features[4473] , \all_features[4474] , \all_features[4475] ,
    \all_features[4476] , \all_features[4477] , \all_features[4478] ,
    \all_features[4479] , \all_features[4480] , \all_features[4481] ,
    \all_features[4482] , \all_features[4483] , \all_features[4484] ,
    \all_features[4485] , \all_features[4486] , \all_features[4487] ,
    \all_features[4488] , \all_features[4489] , \all_features[4490] ,
    \all_features[4491] , \all_features[4492] , \all_features[4493] ,
    \all_features[4494] , \all_features[4495] , \all_features[4496] ,
    \all_features[4497] , \all_features[4498] , \all_features[4499] ,
    \all_features[4500] , \all_features[4501] , \all_features[4502] ,
    \all_features[4503] , \all_features[4504] , \all_features[4505] ,
    \all_features[4506] , \all_features[4507] , \all_features[4508] ,
    \all_features[4509] , \all_features[4510] , \all_features[4511] ,
    \all_features[4512] , \all_features[4513] , \all_features[4514] ,
    \all_features[4515] , \all_features[4516] , \all_features[4517] ,
    \all_features[4518] , \all_features[4519] , \all_features[4520] ,
    \all_features[4521] , \all_features[4522] , \all_features[4523] ,
    \all_features[4524] , \all_features[4525] , \all_features[4526] ,
    \all_features[4527] , \all_features[4528] , \all_features[4529] ,
    \all_features[4530] , \all_features[4531] , \all_features[4532] ,
    \all_features[4533] , \all_features[4534] , \all_features[4535] ,
    \all_features[4536] , \all_features[4537] , \all_features[4538] ,
    \all_features[4539] , \all_features[4540] , \all_features[4541] ,
    \all_features[4542] , \all_features[4543] , \all_features[4544] ,
    \all_features[4545] , \all_features[4546] , \all_features[4547] ,
    \all_features[4548] , \all_features[4549] , \all_features[4550] ,
    \all_features[4551] , \all_features[4552] , \all_features[4553] ,
    \all_features[4554] , \all_features[4555] , \all_features[4556] ,
    \all_features[4557] , \all_features[4558] , \all_features[4559] ,
    \all_features[4560] , \all_features[4561] , \all_features[4562] ,
    \all_features[4563] , \all_features[4564] , \all_features[4565] ,
    \all_features[4566] , \all_features[4567] , \all_features[4568] ,
    \all_features[4569] , \all_features[4570] , \all_features[4571] ,
    \all_features[4572] , \all_features[4573] , \all_features[4574] ,
    \all_features[4575] , \all_features[4576] , \all_features[4577] ,
    \all_features[4578] , \all_features[4579] , \all_features[4580] ,
    \all_features[4581] , \all_features[4582] , \all_features[4583] ,
    \all_features[4584] , \all_features[4585] , \all_features[4586] ,
    \all_features[4587] , \all_features[4588] , \all_features[4589] ,
    \all_features[4590] , \all_features[4591] , \all_features[4592] ,
    \all_features[4593] , \all_features[4594] , \all_features[4595] ,
    \all_features[4596] , \all_features[4597] , \all_features[4598] ,
    \all_features[4599] , \all_features[4600] , \all_features[4601] ,
    \all_features[4602] , \all_features[4603] , \all_features[4604] ,
    \all_features[4605] , \all_features[4606] , \all_features[4607] ,
    \all_features[4608] , \all_features[4609] , \all_features[4610] ,
    \all_features[4611] , \all_features[4612] , \all_features[4613] ,
    \all_features[4614] , \all_features[4615] , \all_features[4616] ,
    \all_features[4617] , \all_features[4618] , \all_features[4619] ,
    \all_features[4620] , \all_features[4621] , \all_features[4622] ,
    \all_features[4623] , \all_features[4624] , \all_features[4625] ,
    \all_features[4626] , \all_features[4627] , \all_features[4628] ,
    \all_features[4629] , \all_features[4630] , \all_features[4631] ,
    \all_features[4632] , \all_features[4633] , \all_features[4634] ,
    \all_features[4635] , \all_features[4636] , \all_features[4637] ,
    \all_features[4638] , \all_features[4639] , \all_features[4640] ,
    \all_features[4641] , \all_features[4642] , \all_features[4643] ,
    \all_features[4644] , \all_features[4645] , \all_features[4646] ,
    \all_features[4647] , \all_features[4648] , \all_features[4649] ,
    \all_features[4650] , \all_features[4651] , \all_features[4652] ,
    \all_features[4653] , \all_features[4654] , \all_features[4655] ,
    \all_features[4656] , \all_features[4657] , \all_features[4658] ,
    \all_features[4659] , \all_features[4660] , \all_features[4661] ,
    \all_features[4662] , \all_features[4663] , \all_features[4664] ,
    \all_features[4665] , \all_features[4666] , \all_features[4667] ,
    \all_features[4668] , \all_features[4669] , \all_features[4670] ,
    \all_features[4671] , \all_features[4672] , \all_features[4673] ,
    \all_features[4674] , \all_features[4675] , \all_features[4676] ,
    \all_features[4677] , \all_features[4678] , \all_features[4679] ,
    \all_features[4680] , \all_features[4681] , \all_features[4682] ,
    \all_features[4683] , \all_features[4684] , \all_features[4685] ,
    \all_features[4686] , \all_features[4687] , \all_features[4688] ,
    \all_features[4689] , \all_features[4690] , \all_features[4691] ,
    \all_features[4692] , \all_features[4693] , \all_features[4694] ,
    \all_features[4695] , \all_features[4696] , \all_features[4697] ,
    \all_features[4698] , \all_features[4699] , \all_features[4700] ,
    \all_features[4701] , \all_features[4702] , \all_features[4703] ,
    \all_features[4704] , \all_features[4705] , \all_features[4706] ,
    \all_features[4707] , \all_features[4708] , \all_features[4709] ,
    \all_features[4710] , \all_features[4711] , \all_features[4712] ,
    \all_features[4713] , \all_features[4714] , \all_features[4715] ,
    \all_features[4716] , \all_features[4717] , \all_features[4718] ,
    \all_features[4719] , \all_features[4720] , \all_features[4721] ,
    \all_features[4722] , \all_features[4723] , \all_features[4724] ,
    \all_features[4725] , \all_features[4726] , \all_features[4727] ,
    \all_features[4728] , \all_features[4729] , \all_features[4730] ,
    \all_features[4731] , \all_features[4732] , \all_features[4733] ,
    \all_features[4734] , \all_features[4735] , \all_features[4736] ,
    \all_features[4737] , \all_features[4738] , \all_features[4739] ,
    \all_features[4740] , \all_features[4741] , \all_features[4742] ,
    \all_features[4743] , \all_features[4744] , \all_features[4745] ,
    \all_features[4746] , \all_features[4747] , \all_features[4748] ,
    \all_features[4749] , \all_features[4750] , \all_features[4751] ,
    \all_features[4752] , \all_features[4753] , \all_features[4754] ,
    \all_features[4755] , \all_features[4756] , \all_features[4757] ,
    \all_features[4758] , \all_features[4759] , \all_features[4760] ,
    \all_features[4761] , \all_features[4762] , \all_features[4763] ,
    \all_features[4764] , \all_features[4765] , \all_features[4766] ,
    \all_features[4767] , \all_features[4768] , \all_features[4769] ,
    \all_features[4770] , \all_features[4771] , \all_features[4772] ,
    \all_features[4773] , \all_features[4774] , \all_features[4775] ,
    \all_features[4776] , \all_features[4777] , \all_features[4778] ,
    \all_features[4779] , \all_features[4780] , \all_features[4781] ,
    \all_features[4782] , \all_features[4783] , \all_features[4784] ,
    \all_features[4785] , \all_features[4786] , \all_features[4787] ,
    \all_features[4788] , \all_features[4789] , \all_features[4790] ,
    \all_features[4791] , \all_features[4792] , \all_features[4793] ,
    \all_features[4794] , \all_features[4795] , \all_features[4796] ,
    \all_features[4797] , \all_features[4798] , \all_features[4799] ,
    \all_features[4800] , \all_features[4801] , \all_features[4802] ,
    \all_features[4803] , \all_features[4804] , \all_features[4805] ,
    \all_features[4806] , \all_features[4807] , \all_features[4808] ,
    \all_features[4809] , \all_features[4810] , \all_features[4811] ,
    \all_features[4812] , \all_features[4813] , \all_features[4814] ,
    \all_features[4815] , \all_features[4816] , \all_features[4817] ,
    \all_features[4818] , \all_features[4819] , \all_features[4820] ,
    \all_features[4821] , \all_features[4822] , \all_features[4823] ,
    \all_features[4824] , \all_features[4825] , \all_features[4826] ,
    \all_features[4827] , \all_features[4828] , \all_features[4829] ,
    \all_features[4830] , \all_features[4831] , \all_features[4832] ,
    \all_features[4833] , \all_features[4834] , \all_features[4835] ,
    \all_features[4836] , \all_features[4837] , \all_features[4838] ,
    \all_features[4839] , \all_features[4840] , \all_features[4841] ,
    \all_features[4842] , \all_features[4843] , \all_features[4844] ,
    \all_features[4845] , \all_features[4846] , \all_features[4847] ,
    \all_features[4848] , \all_features[4849] , \all_features[4850] ,
    \all_features[4851] , \all_features[4852] , \all_features[4853] ,
    \all_features[4854] , \all_features[4855] , \all_features[4856] ,
    \all_features[4857] , \all_features[4858] , \all_features[4859] ,
    \all_features[4860] , \all_features[4861] , \all_features[4862] ,
    \all_features[4863] , \all_features[4864] , \all_features[4865] ,
    \all_features[4866] , \all_features[4867] , \all_features[4868] ,
    \all_features[4869] , \all_features[4870] , \all_features[4871] ,
    \all_features[4872] , \all_features[4873] , \all_features[4874] ,
    \all_features[4875] , \all_features[4876] , \all_features[4877] ,
    \all_features[4878] , \all_features[4879] , \all_features[4880] ,
    \all_features[4881] , \all_features[4882] , \all_features[4883] ,
    \all_features[4884] , \all_features[4885] , \all_features[4886] ,
    \all_features[4887] , \all_features[4888] , \all_features[4889] ,
    \all_features[4890] , \all_features[4891] , \all_features[4892] ,
    \all_features[4893] , \all_features[4894] , \all_features[4895] ,
    \all_features[4896] , \all_features[4897] , \all_features[4898] ,
    \all_features[4899] , \all_features[4900] , \all_features[4901] ,
    \all_features[4902] , \all_features[4903] , \all_features[4904] ,
    \all_features[4905] , \all_features[4906] , \all_features[4907] ,
    \all_features[4908] , \all_features[4909] , \all_features[4910] ,
    \all_features[4911] , \all_features[4912] , \all_features[4913] ,
    \all_features[4914] , \all_features[4915] , \all_features[4916] ,
    \all_features[4917] , \all_features[4918] , \all_features[4919] ,
    \all_features[4920] , \all_features[4921] , \all_features[4922] ,
    \all_features[4923] , \all_features[4924] , \all_features[4925] ,
    \all_features[4926] , \all_features[4927] , \all_features[4928] ,
    \all_features[4929] , \all_features[4930] , \all_features[4931] ,
    \all_features[4932] , \all_features[4933] , \all_features[4934] ,
    \all_features[4935] , \all_features[4936] , \all_features[4937] ,
    \all_features[4938] , \all_features[4939] , \all_features[4940] ,
    \all_features[4941] , \all_features[4942] , \all_features[4943] ,
    \all_features[4944] , \all_features[4945] , \all_features[4946] ,
    \all_features[4947] , \all_features[4948] , \all_features[4949] ,
    \all_features[4950] , \all_features[4951] , \all_features[4952] ,
    \all_features[4953] , \all_features[4954] , \all_features[4955] ,
    \all_features[4956] , \all_features[4957] , \all_features[4958] ,
    \all_features[4959] , \all_features[4960] , \all_features[4961] ,
    \all_features[4962] , \all_features[4963] , \all_features[4964] ,
    \all_features[4965] , \all_features[4966] , \all_features[4967] ,
    \all_features[4968] , \all_features[4969] , \all_features[4970] ,
    \all_features[4971] , \all_features[4972] , \all_features[4973] ,
    \all_features[4974] , \all_features[4975] , \all_features[4976] ,
    \all_features[4977] , \all_features[4978] , \all_features[4979] ,
    \all_features[4980] , \all_features[4981] , \all_features[4982] ,
    \all_features[4983] , \all_features[4984] , \all_features[4985] ,
    \all_features[4986] , \all_features[4987] , \all_features[4988] ,
    \all_features[4989] , \all_features[4990] , \all_features[4991] ,
    \all_features[4992] , \all_features[4993] , \all_features[4994] ,
    \all_features[4995] , \all_features[4996] , \all_features[4997] ,
    \all_features[4998] , \all_features[4999] , \all_features[5000] ,
    \all_features[5001] , \all_features[5002] , \all_features[5003] ,
    \all_features[5004] , \all_features[5005] , \all_features[5006] ,
    \all_features[5007] , \all_features[5008] , \all_features[5009] ,
    \all_features[5010] , \all_features[5011] , \all_features[5012] ,
    \all_features[5013] , \all_features[5014] , \all_features[5015] ,
    \all_features[5016] , \all_features[5017] , \all_features[5018] ,
    \all_features[5019] , \all_features[5020] , \all_features[5021] ,
    \all_features[5022] , \all_features[5023] , \all_features[5024] ,
    \all_features[5025] , \all_features[5026] , \all_features[5027] ,
    \all_features[5028] , \all_features[5029] , \all_features[5030] ,
    \all_features[5031] , \all_features[5032] , \all_features[5033] ,
    \all_features[5034] , \all_features[5035] , \all_features[5036] ,
    \all_features[5037] , \all_features[5038] , \all_features[5039] ,
    \all_features[5040] , \all_features[5041] , \all_features[5042] ,
    \all_features[5043] , \all_features[5044] , \all_features[5045] ,
    \all_features[5046] , \all_features[5047] , \all_features[5048] ,
    \all_features[5049] , \all_features[5050] , \all_features[5051] ,
    \all_features[5052] , \all_features[5053] , \all_features[5054] ,
    \all_features[5055] , \all_features[5056] , \all_features[5057] ,
    \all_features[5058] , \all_features[5059] , \all_features[5060] ,
    \all_features[5061] , \all_features[5062] , \all_features[5063] ,
    \all_features[5064] , \all_features[5065] , \all_features[5066] ,
    \all_features[5067] , \all_features[5068] , \all_features[5069] ,
    \all_features[5070] , \all_features[5071] , \all_features[5072] ,
    \all_features[5073] , \all_features[5074] , \all_features[5075] ,
    \all_features[5076] , \all_features[5077] , \all_features[5078] ,
    \all_features[5079] , \all_features[5080] , \all_features[5081] ,
    \all_features[5082] , \all_features[5083] , \all_features[5084] ,
    \all_features[5085] , \all_features[5086] , \all_features[5087] ,
    \all_features[5088] , \all_features[5089] , \all_features[5090] ,
    \all_features[5091] , \all_features[5092] , \all_features[5093] ,
    \all_features[5094] , \all_features[5095] , \all_features[5096] ,
    \all_features[5097] , \all_features[5098] , \all_features[5099] ,
    \all_features[5100] , \all_features[5101] , \all_features[5102] ,
    \all_features[5103] , \all_features[5104] , \all_features[5105] ,
    \all_features[5106] , \all_features[5107] , \all_features[5108] ,
    \all_features[5109] , \all_features[5110] , \all_features[5111] ,
    \all_features[5112] , \all_features[5113] , \all_features[5114] ,
    \all_features[5115] , \all_features[5116] , \all_features[5117] ,
    \all_features[5118] , \all_features[5119] , \all_features[5120] ,
    \all_features[5121] , \all_features[5122] , \all_features[5123] ,
    \all_features[5124] , \all_features[5125] , \all_features[5126] ,
    \all_features[5127] , \all_features[5128] , \all_features[5129] ,
    \all_features[5130] , \all_features[5131] , \all_features[5132] ,
    \all_features[5133] , \all_features[5134] , \all_features[5135] ,
    \all_features[5136] , \all_features[5137] , \all_features[5138] ,
    \all_features[5139] , \all_features[5140] , \all_features[5141] ,
    \all_features[5142] , \all_features[5143] , \all_features[5144] ,
    \all_features[5145] , \all_features[5146] , \all_features[5147] ,
    \all_features[5148] , \all_features[5149] , \all_features[5150] ,
    \all_features[5151] , \all_features[5152] , \all_features[5153] ,
    \all_features[5154] , \all_features[5155] , \all_features[5156] ,
    \all_features[5157] , \all_features[5158] , \all_features[5159] ,
    \all_features[5160] , \all_features[5161] , \all_features[5162] ,
    \all_features[5163] , \all_features[5164] , \all_features[5165] ,
    \all_features[5166] , \all_features[5167] , \all_features[5168] ,
    \all_features[5169] , \all_features[5170] , \all_features[5171] ,
    \all_features[5172] , \all_features[5173] , \all_features[5174] ,
    \all_features[5175] , \all_features[5176] , \all_features[5177] ,
    \all_features[5178] , \all_features[5179] , \all_features[5180] ,
    \all_features[5181] , \all_features[5182] , \all_features[5183] ,
    \all_features[5184] , \all_features[5185] , \all_features[5186] ,
    \all_features[5187] , \all_features[5188] , \all_features[5189] ,
    \all_features[5190] , \all_features[5191] , \all_features[5192] ,
    \all_features[5193] , \all_features[5194] , \all_features[5195] ,
    \all_features[5196] , \all_features[5197] , \all_features[5198] ,
    \all_features[5199] , \all_features[5200] , \all_features[5201] ,
    \all_features[5202] , \all_features[5203] , \all_features[5204] ,
    \all_features[5205] , \all_features[5206] , \all_features[5207] ,
    \all_features[5208] , \all_features[5209] , \all_features[5210] ,
    \all_features[5211] , \all_features[5212] , \all_features[5213] ,
    \all_features[5214] , \all_features[5215] , \all_features[5216] ,
    \all_features[5217] , \all_features[5218] , \all_features[5219] ,
    \all_features[5220] , \all_features[5221] , \all_features[5222] ,
    \all_features[5223] , \all_features[5224] , \all_features[5225] ,
    \all_features[5226] , \all_features[5227] , \all_features[5228] ,
    \all_features[5229] , \all_features[5230] , \all_features[5231] ,
    \all_features[5232] , \all_features[5233] , \all_features[5234] ,
    \all_features[5235] , \all_features[5236] , \all_features[5237] ,
    \all_features[5238] , \all_features[5239] , \all_features[5240] ,
    \all_features[5241] , \all_features[5242] , \all_features[5243] ,
    \all_features[5244] , \all_features[5245] , \all_features[5246] ,
    \all_features[5247] , \all_features[5248] , \all_features[5249] ,
    \all_features[5250] , \all_features[5251] , \all_features[5252] ,
    \all_features[5253] , \all_features[5254] , \all_features[5255] ,
    \all_features[5256] , \all_features[5257] , \all_features[5258] ,
    \all_features[5259] , \all_features[5260] , \all_features[5261] ,
    \all_features[5262] , \all_features[5263] , \all_features[5264] ,
    \all_features[5265] , \all_features[5266] , \all_features[5267] ,
    \all_features[5268] , \all_features[5269] , \all_features[5270] ,
    \all_features[5271] , \all_features[5272] , \all_features[5273] ,
    \all_features[5274] , \all_features[5275] , \all_features[5276] ,
    \all_features[5277] , \all_features[5278] , \all_features[5279] ,
    \all_features[5280] , \all_features[5281] , \all_features[5282] ,
    \all_features[5283] , \all_features[5284] , \all_features[5285] ,
    \all_features[5286] , \all_features[5287] , \all_features[5288] ,
    \all_features[5289] , \all_features[5290] , \all_features[5291] ,
    \all_features[5292] , \all_features[5293] , \all_features[5294] ,
    \all_features[5295] , \all_features[5296] , \all_features[5297] ,
    \all_features[5298] , \all_features[5299] , \all_features[5300] ,
    \all_features[5301] , \all_features[5302] , \all_features[5303] ,
    \all_features[5304] , \all_features[5305] , \all_features[5306] ,
    \all_features[5307] , \all_features[5308] , \all_features[5309] ,
    \all_features[5310] , \all_features[5311] , \all_features[5312] ,
    \all_features[5313] , \all_features[5314] , \all_features[5315] ,
    \all_features[5316] , \all_features[5317] , \all_features[5318] ,
    \all_features[5319] , \all_features[5320] , \all_features[5321] ,
    \all_features[5322] , \all_features[5323] , \all_features[5324] ,
    \all_features[5325] , \all_features[5326] , \all_features[5327] ,
    \all_features[5328] , \all_features[5329] , \all_features[5330] ,
    \all_features[5331] , \all_features[5332] , \all_features[5333] ,
    \all_features[5334] , \all_features[5335] , \all_features[5336] ,
    \all_features[5337] , \all_features[5338] , \all_features[5339] ,
    \all_features[5340] , \all_features[5341] , \all_features[5342] ,
    \all_features[5343] , \all_features[5344] , \all_features[5345] ,
    \all_features[5346] , \all_features[5347] , \all_features[5348] ,
    \all_features[5349] , \all_features[5350] , \all_features[5351] ,
    \all_features[5352] , \all_features[5353] , \all_features[5354] ,
    \all_features[5355] , \all_features[5356] , \all_features[5357] ,
    \all_features[5358] , \all_features[5359] , \all_features[5360] ,
    \all_features[5361] , \all_features[5362] , \all_features[5363] ,
    \all_features[5364] , \all_features[5365] , \all_features[5366] ,
    \all_features[5367] , \all_features[5368] , \all_features[5369] ,
    \all_features[5370] , \all_features[5371] , \all_features[5372] ,
    \all_features[5373] , \all_features[5374] , \all_features[5375] ,
    \all_features[5376] , \all_features[5377] , \all_features[5378] ,
    \all_features[5379] , \all_features[5380] , \all_features[5381] ,
    \all_features[5382] , \all_features[5383] , \all_features[5384] ,
    \all_features[5385] , \all_features[5386] , \all_features[5387] ,
    \all_features[5388] , \all_features[5389] , \all_features[5390] ,
    \all_features[5391] , \all_features[5392] , \all_features[5393] ,
    \all_features[5394] , \all_features[5395] , \all_features[5396] ,
    \all_features[5397] , \all_features[5398] , \all_features[5399] ,
    \all_features[5400] , \all_features[5401] , \all_features[5402] ,
    \all_features[5403] , \all_features[5404] , \all_features[5405] ,
    \all_features[5406] , \all_features[5407] , \all_features[5408] ,
    \all_features[5409] , \all_features[5410] , \all_features[5411] ,
    \all_features[5412] , \all_features[5413] , \all_features[5414] ,
    \all_features[5415] , \all_features[5416] , \all_features[5417] ,
    \all_features[5418] , \all_features[5419] , \all_features[5420] ,
    \all_features[5421] , \all_features[5422] , \all_features[5423] ,
    \all_features[5424] , \all_features[5425] , \all_features[5426] ,
    \all_features[5427] , \all_features[5428] , \all_features[5429] ,
    \all_features[5430] , \all_features[5431] , \all_features[5432] ,
    \all_features[5433] , \all_features[5434] , \all_features[5435] ,
    \all_features[5436] , \all_features[5437] , \all_features[5438] ,
    \all_features[5439] , \all_features[5440] , \all_features[5441] ,
    \all_features[5442] , \all_features[5443] , \all_features[5444] ,
    \all_features[5445] , \all_features[5446] , \all_features[5447] ,
    \all_features[5448] , \all_features[5449] , \all_features[5450] ,
    \all_features[5451] , \all_features[5452] , \all_features[5453] ,
    \all_features[5454] , \all_features[5455] , \all_features[5456] ,
    \all_features[5457] , \all_features[5458] , \all_features[5459] ,
    \all_features[5460] , \all_features[5461] , \all_features[5462] ,
    \all_features[5463] , \all_features[5464] , \all_features[5465] ,
    \all_features[5466] , \all_features[5467] , \all_features[5468] ,
    \all_features[5469] , \all_features[5470] , \all_features[5471] ,
    \all_features[5472] , \all_features[5473] , \all_features[5474] ,
    \all_features[5475] , \all_features[5476] , \all_features[5477] ,
    \all_features[5478] , \all_features[5479] , \all_features[5480] ,
    \all_features[5481] , \all_features[5482] , \all_features[5483] ,
    \all_features[5484] , \all_features[5485] , \all_features[5486] ,
    \all_features[5487] , \all_features[5488] , \all_features[5489] ,
    \all_features[5490] , \all_features[5491] , \all_features[5492] ,
    \all_features[5493] , \all_features[5494] , \all_features[5495] ,
    \all_features[5496] , \all_features[5497] , \all_features[5498] ,
    \all_features[5499] , \all_features[5500] , \all_features[5501] ,
    \all_features[5502] , \all_features[5503] , \all_features[5504] ,
    \all_features[5505] , \all_features[5506] , \all_features[5507] ,
    \all_features[5508] , \all_features[5509] , \all_features[5510] ,
    \all_features[5511] , \all_features[5512] , \all_features[5513] ,
    \all_features[5514] , \all_features[5515] , \all_features[5516] ,
    \all_features[5517] , \all_features[5518] , \all_features[5519] ,
    \all_features[5520] , \all_features[5521] , \all_features[5522] ,
    \all_features[5523] , \all_features[5524] , \all_features[5525] ,
    \all_features[5526] , \all_features[5527] , \all_features[5528] ,
    \all_features[5529] , \all_features[5530] , \all_features[5531] ,
    \all_features[5532] , \all_features[5533] , \all_features[5534] ,
    \all_features[5535] , \all_features[5536] , \all_features[5537] ,
    \all_features[5538] , \all_features[5539] , \all_features[5540] ,
    \all_features[5541] , \all_features[5542] , \all_features[5543] ,
    \all_features[5544] , \all_features[5545] , \all_features[5546] ,
    \all_features[5547] , \all_features[5548] , \all_features[5549] ,
    \all_features[5550] , \all_features[5551] , \all_features[5552] ,
    \all_features[5553] , \all_features[5554] , \all_features[5555] ,
    \all_features[5556] , \all_features[5557] , \all_features[5558] ,
    \all_features[5559] , \all_features[5560] , \all_features[5561] ,
    \all_features[5562] , \all_features[5563] , \all_features[5564] ,
    \all_features[5565] , \all_features[5566] , \all_features[5567] ,
    \all_features[5568] , \all_features[5569] , \all_features[5570] ,
    \all_features[5571] , \all_features[5572] , \all_features[5573] ,
    \all_features[5574] , \all_features[5575] , \all_features[5576] ,
    \all_features[5577] , \all_features[5578] , \all_features[5579] ,
    \all_features[5580] , \all_features[5581] , \all_features[5582] ,
    \all_features[5583] , \all_features[5584] , \all_features[5585] ,
    \all_features[5586] , \all_features[5587] , \all_features[5588] ,
    \all_features[5589] , \all_features[5590] , \all_features[5591] ,
    \all_features[5592] , \all_features[5593] , \all_features[5594] ,
    \all_features[5595] , \all_features[5596] , \all_features[5597] ,
    \all_features[5598] , \all_features[5599] , \all_features[5600] ,
    \all_features[5601] , \all_features[5602] , \all_features[5603] ,
    \all_features[5604] , \all_features[5605] , \all_features[5606] ,
    \all_features[5607] , \all_features[5608] , \all_features[5609] ,
    \all_features[5610] , \all_features[5611] , \all_features[5612] ,
    \all_features[5613] , \all_features[5614] , \all_features[5615] ,
    \all_features[5616] , \all_features[5617] , \all_features[5618] ,
    \all_features[5619] , \all_features[5620] , \all_features[5621] ,
    \all_features[5622] , \all_features[5623] , \all_features[5624] ,
    \all_features[5625] , \all_features[5626] , \all_features[5627] ,
    \all_features[5628] , \all_features[5629] , \all_features[5630] ,
    \all_features[5631] , \all_features[5632] , \all_features[5633] ,
    \all_features[5634] , \all_features[5635] , \all_features[5636] ,
    \all_features[5637] , \all_features[5638] , \all_features[5639] ,
    \all_features[5640] , \all_features[5641] , \all_features[5642] ,
    \all_features[5643] , \all_features[5644] , \all_features[5645] ,
    \all_features[5646] , \all_features[5647] , \all_features[5648] ,
    \all_features[5649] , \all_features[5650] , \all_features[5651] ,
    \all_features[5652] , \all_features[5653] , \all_features[5654] ,
    \all_features[5655] , \all_features[5656] , \all_features[5657] ,
    \all_features[5658] , \all_features[5659] , \all_features[5660] ,
    \all_features[5661] , \all_features[5662] , \all_features[5663] ,
    \all_features[5664] , \all_features[5665] , \all_features[5666] ,
    \all_features[5667] , \all_features[5668] , \all_features[5669] ,
    \all_features[5670] , \all_features[5671] , \all_features[5672] ,
    \all_features[5673] , \all_features[5674] , \all_features[5675] ,
    \all_features[5676] , \all_features[5677] , \all_features[5678] ,
    \all_features[5679] , \all_features[5680] , \all_features[5681] ,
    \all_features[5682] , \all_features[5683] , \all_features[5684] ,
    \all_features[5685] , \all_features[5686] , \all_features[5687] ,
    \all_features[5688] , \all_features[5689] , \all_features[5690] ,
    \all_features[5691] , \all_features[5692] , \all_features[5693] ,
    \all_features[5694] , \all_features[5695] , \all_features[5696] ,
    \all_features[5697] , \all_features[5698] , \all_features[5699] ,
    \all_features[5700] , \all_features[5701] , \all_features[5702] ,
    \all_features[5703] , \all_features[5704] , \all_features[5705] ,
    \all_features[5706] , \all_features[5707] , \all_features[5708] ,
    \all_features[5709] , \all_features[5710] , \all_features[5711] ,
    \all_features[5712] , \all_features[5713] , \all_features[5714] ,
    \all_features[5715] , \all_features[5716] , \all_features[5717] ,
    \all_features[5718] , \all_features[5719] , \all_features[5720] ,
    \all_features[5721] , \all_features[5722] , \all_features[5723] ,
    \all_features[5724] , \all_features[5725] , \all_features[5726] ,
    \all_features[5727] , \all_features[5728] , \all_features[5729] ,
    \all_features[5730] , \all_features[5731] , \all_features[5732] ,
    \all_features[5733] , \all_features[5734] , \all_features[5735] ,
    \all_features[5736] , \all_features[5737] , \all_features[5738] ,
    \all_features[5739] , \all_features[5740] , \all_features[5741] ,
    \all_features[5742] , \all_features[5743] , \all_features[5744] ,
    \all_features[5745] , \all_features[5746] , \all_features[5747] ,
    \all_features[5748] , \all_features[5749] , \all_features[5750] ,
    \all_features[5751] , \all_features[5752] , \all_features[5753] ,
    \all_features[5754] , \all_features[5755] , \all_features[5756] ,
    \all_features[5757] , \all_features[5758] , \all_features[5759] ,
    \all_features[5760] , \all_features[5761] , \all_features[5762] ,
    \all_features[5763] , \all_features[5764] , \all_features[5765] ,
    \all_features[5766] , \all_features[5767] , \all_features[5768] ,
    \all_features[5769] , \all_features[5770] , \all_features[5771] ,
    \all_features[5772] , \all_features[5773] , \all_features[5774] ,
    \all_features[5775] , \all_features[5776] , \all_features[5777] ,
    \all_features[5778] , \all_features[5779] , \all_features[5780] ,
    \all_features[5781] , \all_features[5782] , \all_features[5783] ,
    \all_features[5784] , \all_features[5785] , \all_features[5786] ,
    \all_features[5787] , \all_features[5788] , \all_features[5789] ,
    \all_features[5790] , \all_features[5791] , \all_features[5792] ,
    \all_features[5793] , \all_features[5794] , \all_features[5795] ,
    \all_features[5796] , \all_features[5797] , \all_features[5798] ,
    \all_features[5799] , \all_features[5800] , \all_features[5801] ,
    \all_features[5802] , \all_features[5803] , \all_features[5804] ,
    \all_features[5805] , \all_features[5806] , \all_features[5807] ,
    \all_features[5808] , \all_features[5809] , \all_features[5810] ,
    \all_features[5811] , \all_features[5812] , \all_features[5813] ,
    \all_features[5814] , \all_features[5815] , \all_features[5816] ,
    \all_features[5817] , \all_features[5818] , \all_features[5819] ,
    \all_features[5820] , \all_features[5821] , \all_features[5822] ,
    \all_features[5823] , \all_features[5824] , \all_features[5825] ,
    \all_features[5826] , \all_features[5827] , \all_features[5828] ,
    \all_features[5829] , \all_features[5830] , \all_features[5831] ,
    \all_features[5832] , \all_features[5833] , \all_features[5834] ,
    \all_features[5835] , \all_features[5836] , \all_features[5837] ,
    \all_features[5838] , \all_features[5839] , \all_features[5840] ,
    \all_features[5841] , \all_features[5842] , \all_features[5843] ,
    \all_features[5844] , \all_features[5845] , \all_features[5846] ,
    \all_features[5847] , \all_features[5848] , \all_features[5849] ,
    \all_features[5850] , \all_features[5851] , \all_features[5852] ,
    \all_features[5853] , \all_features[5854] , \all_features[5855] ,
    \all_features[5856] , \all_features[5857] , \all_features[5858] ,
    \all_features[5859] , \all_features[5860] , \all_features[5861] ,
    \all_features[5862] , \all_features[5863] , \all_features[5864] ,
    \all_features[5865] , \all_features[5866] , \all_features[5867] ,
    \all_features[5868] , \all_features[5869] , \all_features[5870] ,
    \all_features[5871] , \all_features[5872] , \all_features[5873] ,
    \all_features[5874] , \all_features[5875] , \all_features[5876] ,
    \all_features[5877] , \all_features[5878] , \all_features[5879] ,
    \all_features[5880] , \all_features[5881] , \all_features[5882] ,
    \all_features[5883] , \all_features[5884] , \all_features[5885] ,
    \all_features[5886] , \all_features[5887] , \all_features[5888] ,
    \all_features[5889] , \all_features[5890] , \all_features[5891] ,
    \all_features[5892] , \all_features[5893] , \all_features[5894] ,
    \all_features[5895] , \all_features[5896] , \all_features[5897] ,
    \all_features[5898] , \all_features[5899] , \all_features[5900] ,
    \all_features[5901] , \all_features[5902] , \all_features[5903] ,
    \all_features[5904] , \all_features[5905] , \all_features[5906] ,
    \all_features[5907] , \all_features[5908] , \all_features[5909] ,
    \all_features[5910] , \all_features[5911] , \all_features[5912] ,
    \all_features[5913] , \all_features[5914] , \all_features[5915] ,
    \all_features[5916] , \all_features[5917] , \all_features[5918] ,
    \all_features[5919] , \all_features[5920] , \all_features[5921] ,
    \all_features[5922] , \all_features[5923] , \all_features[5924] ,
    \all_features[5925] , \all_features[5926] , \all_features[5927] ,
    \all_features[5928] , \all_features[5929] , \all_features[5930] ,
    \all_features[5931] , \all_features[5932] , \all_features[5933] ,
    \all_features[5934] , \all_features[5935] , \all_features[5936] ,
    \all_features[5937] , \all_features[5938] , \all_features[5939] ,
    \all_features[5940] , \all_features[5941] , \all_features[5942] ,
    \all_features[5943] , \all_features[5944] , \all_features[5945] ,
    \all_features[5946] , \all_features[5947] , \all_features[5948] ,
    \all_features[5949] , \all_features[5950] , \all_features[5951] ,
    \all_features[5952] , \all_features[5953] , \all_features[5954] ,
    \all_features[5955] , \all_features[5956] , \all_features[5957] ,
    \all_features[5958] , \all_features[5959] , \all_features[5960] ,
    \all_features[5961] , \all_features[5962] , \all_features[5963] ,
    \all_features[5964] , \all_features[5965] , \all_features[5966] ,
    \all_features[5967] , \all_features[5968] , \all_features[5969] ,
    \all_features[5970] , \all_features[5971] , \all_features[5972] ,
    \all_features[5973] , \all_features[5974] , \all_features[5975] ,
    \all_features[5976] , \all_features[5977] , \all_features[5978] ,
    \all_features[5979] , \all_features[5980] , \all_features[5981] ,
    \all_features[5982] , \all_features[5983] , \all_features[5984] ,
    \all_features[5985] , \all_features[5986] , \all_features[5987] ,
    \all_features[5988] , \all_features[5989] , \all_features[5990] ,
    \all_features[5991] , \all_features[5992] , \all_features[5993] ,
    \all_features[5994] , \all_features[5995] , \all_features[5996] ,
    \all_features[5997] , \all_features[5998] , \all_features[5999] ,
    \all_features[6000] , \all_features[6001] , \all_features[6002] ,
    \all_features[6003] , \all_features[6004] , \all_features[6005] ,
    \all_features[6006] , \all_features[6007] , \all_features[6008] ,
    \all_features[6009] , \all_features[6010] , \all_features[6011] ,
    \all_features[6012] , \all_features[6013] , \all_features[6014] ,
    \all_features[6015] , \all_features[6016] , \all_features[6017] ,
    \all_features[6018] , \all_features[6019] , \all_features[6020] ,
    \all_features[6021] , \all_features[6022] , \all_features[6023] ,
    \all_features[6024] , \all_features[6025] , \all_features[6026] ,
    \all_features[6027] , \all_features[6028] , \all_features[6029] ,
    \all_features[6030] , \all_features[6031] , \all_features[6032] ,
    \all_features[6033] , \all_features[6034] , \all_features[6035] ,
    \all_features[6036] , \all_features[6037] , \all_features[6038] ,
    \all_features[6039] , \all_features[6040] , \all_features[6041] ,
    \all_features[6042] , \all_features[6043] , \all_features[6044] ,
    \all_features[6045] , \all_features[6046] , \all_features[6047] ,
    \all_features[6048] , \all_features[6049] , \all_features[6050] ,
    \all_features[6051] , \all_features[6052] , \all_features[6053] ,
    \all_features[6054] , \all_features[6055] , \all_features[6056] ,
    \all_features[6057] , \all_features[6058] , \all_features[6059] ,
    \all_features[6060] , \all_features[6061] , \all_features[6062] ,
    \all_features[6063] , \all_features[6064] , \all_features[6065] ,
    \all_features[6066] , \all_features[6067] , \all_features[6068] ,
    \all_features[6069] , \all_features[6070] , \all_features[6071] ,
    \all_features[6072] , \all_features[6073] , \all_features[6074] ,
    \all_features[6075] , \all_features[6076] , \all_features[6077] ,
    \all_features[6078] , \all_features[6079] , \all_features[6080] ,
    \all_features[6081] , \all_features[6082] , \all_features[6083] ,
    \all_features[6084] , \all_features[6085] , \all_features[6086] ,
    \all_features[6087] , \all_features[6088] , \all_features[6089] ,
    \all_features[6090] , \all_features[6091] , \all_features[6092] ,
    \all_features[6093] , \all_features[6094] , \all_features[6095] ,
    \all_features[6096] , \all_features[6097] , \all_features[6098] ,
    \all_features[6099] , \all_features[6100] , \all_features[6101] ,
    \all_features[6102] , \all_features[6103] , \all_features[6104] ,
    \all_features[6105] , \all_features[6106] , \all_features[6107] ,
    \all_features[6108] , \all_features[6109] , \all_features[6110] ,
    \all_features[6111] , \all_features[6112] , \all_features[6113] ,
    \all_features[6114] , \all_features[6115] , \all_features[6116] ,
    \all_features[6117] , \all_features[6118] , \all_features[6119] ,
    \all_features[6120] , \all_features[6121] , \all_features[6122] ,
    \all_features[6123] , \all_features[6124] , \all_features[6125] ,
    \all_features[6126] , \all_features[6127] , \all_features[6128] ,
    \all_features[6129] , \all_features[6130] , \all_features[6131] ,
    \all_features[6132] , \all_features[6133] , \all_features[6134] ,
    \all_features[6135] , \all_features[6136] , \all_features[6137] ,
    \all_features[6138] , \all_features[6139] , \all_features[6140] ,
    \all_features[6141] , \all_features[6142] , \all_features[6143] ,
    \all_features[6144] , \all_features[6145] , \all_features[6146] ,
    \all_features[6147] , \all_features[6148] , \all_features[6149] ,
    \all_features[6150] , \all_features[6151] , \all_features[6152] ,
    \all_features[6153] , \all_features[6154] , \all_features[6155] ,
    \all_features[6156] , \all_features[6157] , \all_features[6158] ,
    \all_features[6159] , \all_features[6160] , \all_features[6161] ,
    \all_features[6162] , \all_features[6163] , \all_features[6164] ,
    \all_features[6165] , \all_features[6166] , \all_features[6167] ,
    \all_features[6168] , \all_features[6169] , \all_features[6170] ,
    \all_features[6171] , \all_features[6172] , \all_features[6173] ,
    \all_features[6174] , \all_features[6175] , \all_features[6176] ,
    \all_features[6177] , \all_features[6178] , \all_features[6179] ,
    \all_features[6180] , \all_features[6181] , \all_features[6182] ,
    \all_features[6183] , \all_features[6184] , \all_features[6185] ,
    \all_features[6186] , \all_features[6187] , \all_features[6188] ,
    \all_features[6189] , \all_features[6190] , \all_features[6191] ,
    \all_features[6192] , \all_features[6193] , \all_features[6194] ,
    \all_features[6195] , \all_features[6196] , \all_features[6197] ,
    \all_features[6198] , \all_features[6199] , \all_features[6200] ,
    \all_features[6201] , \all_features[6202] , \all_features[6203] ,
    \all_features[6204] , \all_features[6205] , \all_features[6206] ,
    \all_features[6207] , \all_features[6208] , \all_features[6209] ,
    \all_features[6210] , \all_features[6211] , \all_features[6212] ,
    \all_features[6213] , \all_features[6214] , \all_features[6215] ,
    \all_features[6216] , \all_features[6217] , \all_features[6218] ,
    \all_features[6219] , \all_features[6220] , \all_features[6221] ,
    \all_features[6222] , \all_features[6223] , \all_features[6224] ,
    \all_features[6225] , \all_features[6226] , \all_features[6227] ,
    \all_features[6228] , \all_features[6229] , \all_features[6230] ,
    \all_features[6231] , \all_features[6232] , \all_features[6233] ,
    \all_features[6234] , \all_features[6235] , \all_features[6236] ,
    \all_features[6237] , \all_features[6238] , \all_features[6239] ,
    \all_features[6240] , \all_features[6241] , \all_features[6242] ,
    \all_features[6243] , \all_features[6244] , \all_features[6245] ,
    \all_features[6246] , \all_features[6247] , \all_features[6248] ,
    \all_features[6249] , \all_features[6250] , \all_features[6251] ,
    \all_features[6252] , \all_features[6253] , \all_features[6254] ,
    \all_features[6255] , \all_features[6256] , \all_features[6257] ,
    \all_features[6258] , \all_features[6259] , \all_features[6260] ,
    \all_features[6261] , \all_features[6262] , \all_features[6263] ,
    \all_features[6264] , \all_features[6265] , \all_features[6266] ,
    \all_features[6267] , \all_features[6268] , \all_features[6269] ,
    \all_features[6270] , \all_features[6271] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] ,
    \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] ,
    \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] ,
    \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] ,
    \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] ,
    \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] , \o[64] ,
    \o[65] , \o[66] , \o[67] , \o[68] , \o[69]   );
  input  \all_features[0] , \all_features[1] , \all_features[2] ,
    \all_features[3] , \all_features[4] , \all_features[5] ,
    \all_features[6] , \all_features[7] , \all_features[8] ,
    \all_features[9] , \all_features[10] , \all_features[11] ,
    \all_features[12] , \all_features[13] , \all_features[14] ,
    \all_features[15] , \all_features[16] , \all_features[17] ,
    \all_features[18] , \all_features[19] , \all_features[20] ,
    \all_features[21] , \all_features[22] , \all_features[23] ,
    \all_features[24] , \all_features[25] , \all_features[26] ,
    \all_features[27] , \all_features[28] , \all_features[29] ,
    \all_features[30] , \all_features[31] , \all_features[32] ,
    \all_features[33] , \all_features[34] , \all_features[35] ,
    \all_features[36] , \all_features[37] , \all_features[38] ,
    \all_features[39] , \all_features[40] , \all_features[41] ,
    \all_features[42] , \all_features[43] , \all_features[44] ,
    \all_features[45] , \all_features[46] , \all_features[47] ,
    \all_features[48] , \all_features[49] , \all_features[50] ,
    \all_features[51] , \all_features[52] , \all_features[53] ,
    \all_features[54] , \all_features[55] , \all_features[56] ,
    \all_features[57] , \all_features[58] , \all_features[59] ,
    \all_features[60] , \all_features[61] , \all_features[62] ,
    \all_features[63] , \all_features[64] , \all_features[65] ,
    \all_features[66] , \all_features[67] , \all_features[68] ,
    \all_features[69] , \all_features[70] , \all_features[71] ,
    \all_features[72] , \all_features[73] , \all_features[74] ,
    \all_features[75] , \all_features[76] , \all_features[77] ,
    \all_features[78] , \all_features[79] , \all_features[80] ,
    \all_features[81] , \all_features[82] , \all_features[83] ,
    \all_features[84] , \all_features[85] , \all_features[86] ,
    \all_features[87] , \all_features[88] , \all_features[89] ,
    \all_features[90] , \all_features[91] , \all_features[92] ,
    \all_features[93] , \all_features[94] , \all_features[95] ,
    \all_features[96] , \all_features[97] , \all_features[98] ,
    \all_features[99] , \all_features[100] , \all_features[101] ,
    \all_features[102] , \all_features[103] , \all_features[104] ,
    \all_features[105] , \all_features[106] , \all_features[107] ,
    \all_features[108] , \all_features[109] , \all_features[110] ,
    \all_features[111] , \all_features[112] , \all_features[113] ,
    \all_features[114] , \all_features[115] , \all_features[116] ,
    \all_features[117] , \all_features[118] , \all_features[119] ,
    \all_features[120] , \all_features[121] , \all_features[122] ,
    \all_features[123] , \all_features[124] , \all_features[125] ,
    \all_features[126] , \all_features[127] , \all_features[128] ,
    \all_features[129] , \all_features[130] , \all_features[131] ,
    \all_features[132] , \all_features[133] , \all_features[134] ,
    \all_features[135] , \all_features[136] , \all_features[137] ,
    \all_features[138] , \all_features[139] , \all_features[140] ,
    \all_features[141] , \all_features[142] , \all_features[143] ,
    \all_features[144] , \all_features[145] , \all_features[146] ,
    \all_features[147] , \all_features[148] , \all_features[149] ,
    \all_features[150] , \all_features[151] , \all_features[152] ,
    \all_features[153] , \all_features[154] , \all_features[155] ,
    \all_features[156] , \all_features[157] , \all_features[158] ,
    \all_features[159] , \all_features[160] , \all_features[161] ,
    \all_features[162] , \all_features[163] , \all_features[164] ,
    \all_features[165] , \all_features[166] , \all_features[167] ,
    \all_features[168] , \all_features[169] , \all_features[170] ,
    \all_features[171] , \all_features[172] , \all_features[173] ,
    \all_features[174] , \all_features[175] , \all_features[176] ,
    \all_features[177] , \all_features[178] , \all_features[179] ,
    \all_features[180] , \all_features[181] , \all_features[182] ,
    \all_features[183] , \all_features[184] , \all_features[185] ,
    \all_features[186] , \all_features[187] , \all_features[188] ,
    \all_features[189] , \all_features[190] , \all_features[191] ,
    \all_features[192] , \all_features[193] , \all_features[194] ,
    \all_features[195] , \all_features[196] , \all_features[197] ,
    \all_features[198] , \all_features[199] , \all_features[200] ,
    \all_features[201] , \all_features[202] , \all_features[203] ,
    \all_features[204] , \all_features[205] , \all_features[206] ,
    \all_features[207] , \all_features[208] , \all_features[209] ,
    \all_features[210] , \all_features[211] , \all_features[212] ,
    \all_features[213] , \all_features[214] , \all_features[215] ,
    \all_features[216] , \all_features[217] , \all_features[218] ,
    \all_features[219] , \all_features[220] , \all_features[221] ,
    \all_features[222] , \all_features[223] , \all_features[224] ,
    \all_features[225] , \all_features[226] , \all_features[227] ,
    \all_features[228] , \all_features[229] , \all_features[230] ,
    \all_features[231] , \all_features[232] , \all_features[233] ,
    \all_features[234] , \all_features[235] , \all_features[236] ,
    \all_features[237] , \all_features[238] , \all_features[239] ,
    \all_features[240] , \all_features[241] , \all_features[242] ,
    \all_features[243] , \all_features[244] , \all_features[245] ,
    \all_features[246] , \all_features[247] , \all_features[248] ,
    \all_features[249] , \all_features[250] , \all_features[251] ,
    \all_features[252] , \all_features[253] , \all_features[254] ,
    \all_features[255] , \all_features[256] , \all_features[257] ,
    \all_features[258] , \all_features[259] , \all_features[260] ,
    \all_features[261] , \all_features[262] , \all_features[263] ,
    \all_features[264] , \all_features[265] , \all_features[266] ,
    \all_features[267] , \all_features[268] , \all_features[269] ,
    \all_features[270] , \all_features[271] , \all_features[272] ,
    \all_features[273] , \all_features[274] , \all_features[275] ,
    \all_features[276] , \all_features[277] , \all_features[278] ,
    \all_features[279] , \all_features[280] , \all_features[281] ,
    \all_features[282] , \all_features[283] , \all_features[284] ,
    \all_features[285] , \all_features[286] , \all_features[287] ,
    \all_features[288] , \all_features[289] , \all_features[290] ,
    \all_features[291] , \all_features[292] , \all_features[293] ,
    \all_features[294] , \all_features[295] , \all_features[296] ,
    \all_features[297] , \all_features[298] , \all_features[299] ,
    \all_features[300] , \all_features[301] , \all_features[302] ,
    \all_features[303] , \all_features[304] , \all_features[305] ,
    \all_features[306] , \all_features[307] , \all_features[308] ,
    \all_features[309] , \all_features[310] , \all_features[311] ,
    \all_features[312] , \all_features[313] , \all_features[314] ,
    \all_features[315] , \all_features[316] , \all_features[317] ,
    \all_features[318] , \all_features[319] , \all_features[320] ,
    \all_features[321] , \all_features[322] , \all_features[323] ,
    \all_features[324] , \all_features[325] , \all_features[326] ,
    \all_features[327] , \all_features[328] , \all_features[329] ,
    \all_features[330] , \all_features[331] , \all_features[332] ,
    \all_features[333] , \all_features[334] , \all_features[335] ,
    \all_features[336] , \all_features[337] , \all_features[338] ,
    \all_features[339] , \all_features[340] , \all_features[341] ,
    \all_features[342] , \all_features[343] , \all_features[344] ,
    \all_features[345] , \all_features[346] , \all_features[347] ,
    \all_features[348] , \all_features[349] , \all_features[350] ,
    \all_features[351] , \all_features[352] , \all_features[353] ,
    \all_features[354] , \all_features[355] , \all_features[356] ,
    \all_features[357] , \all_features[358] , \all_features[359] ,
    \all_features[360] , \all_features[361] , \all_features[362] ,
    \all_features[363] , \all_features[364] , \all_features[365] ,
    \all_features[366] , \all_features[367] , \all_features[368] ,
    \all_features[369] , \all_features[370] , \all_features[371] ,
    \all_features[372] , \all_features[373] , \all_features[374] ,
    \all_features[375] , \all_features[376] , \all_features[377] ,
    \all_features[378] , \all_features[379] , \all_features[380] ,
    \all_features[381] , \all_features[382] , \all_features[383] ,
    \all_features[384] , \all_features[385] , \all_features[386] ,
    \all_features[387] , \all_features[388] , \all_features[389] ,
    \all_features[390] , \all_features[391] , \all_features[392] ,
    \all_features[393] , \all_features[394] , \all_features[395] ,
    \all_features[396] , \all_features[397] , \all_features[398] ,
    \all_features[399] , \all_features[400] , \all_features[401] ,
    \all_features[402] , \all_features[403] , \all_features[404] ,
    \all_features[405] , \all_features[406] , \all_features[407] ,
    \all_features[408] , \all_features[409] , \all_features[410] ,
    \all_features[411] , \all_features[412] , \all_features[413] ,
    \all_features[414] , \all_features[415] , \all_features[416] ,
    \all_features[417] , \all_features[418] , \all_features[419] ,
    \all_features[420] , \all_features[421] , \all_features[422] ,
    \all_features[423] , \all_features[424] , \all_features[425] ,
    \all_features[426] , \all_features[427] , \all_features[428] ,
    \all_features[429] , \all_features[430] , \all_features[431] ,
    \all_features[432] , \all_features[433] , \all_features[434] ,
    \all_features[435] , \all_features[436] , \all_features[437] ,
    \all_features[438] , \all_features[439] , \all_features[440] ,
    \all_features[441] , \all_features[442] , \all_features[443] ,
    \all_features[444] , \all_features[445] , \all_features[446] ,
    \all_features[447] , \all_features[448] , \all_features[449] ,
    \all_features[450] , \all_features[451] , \all_features[452] ,
    \all_features[453] , \all_features[454] , \all_features[455] ,
    \all_features[456] , \all_features[457] , \all_features[458] ,
    \all_features[459] , \all_features[460] , \all_features[461] ,
    \all_features[462] , \all_features[463] , \all_features[464] ,
    \all_features[465] , \all_features[466] , \all_features[467] ,
    \all_features[468] , \all_features[469] , \all_features[470] ,
    \all_features[471] , \all_features[472] , \all_features[473] ,
    \all_features[474] , \all_features[475] , \all_features[476] ,
    \all_features[477] , \all_features[478] , \all_features[479] ,
    \all_features[480] , \all_features[481] , \all_features[482] ,
    \all_features[483] , \all_features[484] , \all_features[485] ,
    \all_features[486] , \all_features[487] , \all_features[488] ,
    \all_features[489] , \all_features[490] , \all_features[491] ,
    \all_features[492] , \all_features[493] , \all_features[494] ,
    \all_features[495] , \all_features[496] , \all_features[497] ,
    \all_features[498] , \all_features[499] , \all_features[500] ,
    \all_features[501] , \all_features[502] , \all_features[503] ,
    \all_features[504] , \all_features[505] , \all_features[506] ,
    \all_features[507] , \all_features[508] , \all_features[509] ,
    \all_features[510] , \all_features[511] , \all_features[512] ,
    \all_features[513] , \all_features[514] , \all_features[515] ,
    \all_features[516] , \all_features[517] , \all_features[518] ,
    \all_features[519] , \all_features[520] , \all_features[521] ,
    \all_features[522] , \all_features[523] , \all_features[524] ,
    \all_features[525] , \all_features[526] , \all_features[527] ,
    \all_features[528] , \all_features[529] , \all_features[530] ,
    \all_features[531] , \all_features[532] , \all_features[533] ,
    \all_features[534] , \all_features[535] , \all_features[536] ,
    \all_features[537] , \all_features[538] , \all_features[539] ,
    \all_features[540] , \all_features[541] , \all_features[542] ,
    \all_features[543] , \all_features[544] , \all_features[545] ,
    \all_features[546] , \all_features[547] , \all_features[548] ,
    \all_features[549] , \all_features[550] , \all_features[551] ,
    \all_features[552] , \all_features[553] , \all_features[554] ,
    \all_features[555] , \all_features[556] , \all_features[557] ,
    \all_features[558] , \all_features[559] , \all_features[560] ,
    \all_features[561] , \all_features[562] , \all_features[563] ,
    \all_features[564] , \all_features[565] , \all_features[566] ,
    \all_features[567] , \all_features[568] , \all_features[569] ,
    \all_features[570] , \all_features[571] , \all_features[572] ,
    \all_features[573] , \all_features[574] , \all_features[575] ,
    \all_features[576] , \all_features[577] , \all_features[578] ,
    \all_features[579] , \all_features[580] , \all_features[581] ,
    \all_features[582] , \all_features[583] , \all_features[584] ,
    \all_features[585] , \all_features[586] , \all_features[587] ,
    \all_features[588] , \all_features[589] , \all_features[590] ,
    \all_features[591] , \all_features[592] , \all_features[593] ,
    \all_features[594] , \all_features[595] , \all_features[596] ,
    \all_features[597] , \all_features[598] , \all_features[599] ,
    \all_features[600] , \all_features[601] , \all_features[602] ,
    \all_features[603] , \all_features[604] , \all_features[605] ,
    \all_features[606] , \all_features[607] , \all_features[608] ,
    \all_features[609] , \all_features[610] , \all_features[611] ,
    \all_features[612] , \all_features[613] , \all_features[614] ,
    \all_features[615] , \all_features[616] , \all_features[617] ,
    \all_features[618] , \all_features[619] , \all_features[620] ,
    \all_features[621] , \all_features[622] , \all_features[623] ,
    \all_features[624] , \all_features[625] , \all_features[626] ,
    \all_features[627] , \all_features[628] , \all_features[629] ,
    \all_features[630] , \all_features[631] , \all_features[632] ,
    \all_features[633] , \all_features[634] , \all_features[635] ,
    \all_features[636] , \all_features[637] , \all_features[638] ,
    \all_features[639] , \all_features[640] , \all_features[641] ,
    \all_features[642] , \all_features[643] , \all_features[644] ,
    \all_features[645] , \all_features[646] , \all_features[647] ,
    \all_features[648] , \all_features[649] , \all_features[650] ,
    \all_features[651] , \all_features[652] , \all_features[653] ,
    \all_features[654] , \all_features[655] , \all_features[656] ,
    \all_features[657] , \all_features[658] , \all_features[659] ,
    \all_features[660] , \all_features[661] , \all_features[662] ,
    \all_features[663] , \all_features[664] , \all_features[665] ,
    \all_features[666] , \all_features[667] , \all_features[668] ,
    \all_features[669] , \all_features[670] , \all_features[671] ,
    \all_features[672] , \all_features[673] , \all_features[674] ,
    \all_features[675] , \all_features[676] , \all_features[677] ,
    \all_features[678] , \all_features[679] , \all_features[680] ,
    \all_features[681] , \all_features[682] , \all_features[683] ,
    \all_features[684] , \all_features[685] , \all_features[686] ,
    \all_features[687] , \all_features[688] , \all_features[689] ,
    \all_features[690] , \all_features[691] , \all_features[692] ,
    \all_features[693] , \all_features[694] , \all_features[695] ,
    \all_features[696] , \all_features[697] , \all_features[698] ,
    \all_features[699] , \all_features[700] , \all_features[701] ,
    \all_features[702] , \all_features[703] , \all_features[704] ,
    \all_features[705] , \all_features[706] , \all_features[707] ,
    \all_features[708] , \all_features[709] , \all_features[710] ,
    \all_features[711] , \all_features[712] , \all_features[713] ,
    \all_features[714] , \all_features[715] , \all_features[716] ,
    \all_features[717] , \all_features[718] , \all_features[719] ,
    \all_features[720] , \all_features[721] , \all_features[722] ,
    \all_features[723] , \all_features[724] , \all_features[725] ,
    \all_features[726] , \all_features[727] , \all_features[728] ,
    \all_features[729] , \all_features[730] , \all_features[731] ,
    \all_features[732] , \all_features[733] , \all_features[734] ,
    \all_features[735] , \all_features[736] , \all_features[737] ,
    \all_features[738] , \all_features[739] , \all_features[740] ,
    \all_features[741] , \all_features[742] , \all_features[743] ,
    \all_features[744] , \all_features[745] , \all_features[746] ,
    \all_features[747] , \all_features[748] , \all_features[749] ,
    \all_features[750] , \all_features[751] , \all_features[752] ,
    \all_features[753] , \all_features[754] , \all_features[755] ,
    \all_features[756] , \all_features[757] , \all_features[758] ,
    \all_features[759] , \all_features[760] , \all_features[761] ,
    \all_features[762] , \all_features[763] , \all_features[764] ,
    \all_features[765] , \all_features[766] , \all_features[767] ,
    \all_features[768] , \all_features[769] , \all_features[770] ,
    \all_features[771] , \all_features[772] , \all_features[773] ,
    \all_features[774] , \all_features[775] , \all_features[776] ,
    \all_features[777] , \all_features[778] , \all_features[779] ,
    \all_features[780] , \all_features[781] , \all_features[782] ,
    \all_features[783] , \all_features[784] , \all_features[785] ,
    \all_features[786] , \all_features[787] , \all_features[788] ,
    \all_features[789] , \all_features[790] , \all_features[791] ,
    \all_features[792] , \all_features[793] , \all_features[794] ,
    \all_features[795] , \all_features[796] , \all_features[797] ,
    \all_features[798] , \all_features[799] , \all_features[800] ,
    \all_features[801] , \all_features[802] , \all_features[803] ,
    \all_features[804] , \all_features[805] , \all_features[806] ,
    \all_features[807] , \all_features[808] , \all_features[809] ,
    \all_features[810] , \all_features[811] , \all_features[812] ,
    \all_features[813] , \all_features[814] , \all_features[815] ,
    \all_features[816] , \all_features[817] , \all_features[818] ,
    \all_features[819] , \all_features[820] , \all_features[821] ,
    \all_features[822] , \all_features[823] , \all_features[824] ,
    \all_features[825] , \all_features[826] , \all_features[827] ,
    \all_features[828] , \all_features[829] , \all_features[830] ,
    \all_features[831] , \all_features[832] , \all_features[833] ,
    \all_features[834] , \all_features[835] , \all_features[836] ,
    \all_features[837] , \all_features[838] , \all_features[839] ,
    \all_features[840] , \all_features[841] , \all_features[842] ,
    \all_features[843] , \all_features[844] , \all_features[845] ,
    \all_features[846] , \all_features[847] , \all_features[848] ,
    \all_features[849] , \all_features[850] , \all_features[851] ,
    \all_features[852] , \all_features[853] , \all_features[854] ,
    \all_features[855] , \all_features[856] , \all_features[857] ,
    \all_features[858] , \all_features[859] , \all_features[860] ,
    \all_features[861] , \all_features[862] , \all_features[863] ,
    \all_features[864] , \all_features[865] , \all_features[866] ,
    \all_features[867] , \all_features[868] , \all_features[869] ,
    \all_features[870] , \all_features[871] , \all_features[872] ,
    \all_features[873] , \all_features[874] , \all_features[875] ,
    \all_features[876] , \all_features[877] , \all_features[878] ,
    \all_features[879] , \all_features[880] , \all_features[881] ,
    \all_features[882] , \all_features[883] , \all_features[884] ,
    \all_features[885] , \all_features[886] , \all_features[887] ,
    \all_features[888] , \all_features[889] , \all_features[890] ,
    \all_features[891] , \all_features[892] , \all_features[893] ,
    \all_features[894] , \all_features[895] , \all_features[896] ,
    \all_features[897] , \all_features[898] , \all_features[899] ,
    \all_features[900] , \all_features[901] , \all_features[902] ,
    \all_features[903] , \all_features[904] , \all_features[905] ,
    \all_features[906] , \all_features[907] , \all_features[908] ,
    \all_features[909] , \all_features[910] , \all_features[911] ,
    \all_features[912] , \all_features[913] , \all_features[914] ,
    \all_features[915] , \all_features[916] , \all_features[917] ,
    \all_features[918] , \all_features[919] , \all_features[920] ,
    \all_features[921] , \all_features[922] , \all_features[923] ,
    \all_features[924] , \all_features[925] , \all_features[926] ,
    \all_features[927] , \all_features[928] , \all_features[929] ,
    \all_features[930] , \all_features[931] , \all_features[932] ,
    \all_features[933] , \all_features[934] , \all_features[935] ,
    \all_features[936] , \all_features[937] , \all_features[938] ,
    \all_features[939] , \all_features[940] , \all_features[941] ,
    \all_features[942] , \all_features[943] , \all_features[944] ,
    \all_features[945] , \all_features[946] , \all_features[947] ,
    \all_features[948] , \all_features[949] , \all_features[950] ,
    \all_features[951] , \all_features[952] , \all_features[953] ,
    \all_features[954] , \all_features[955] , \all_features[956] ,
    \all_features[957] , \all_features[958] , \all_features[959] ,
    \all_features[960] , \all_features[961] , \all_features[962] ,
    \all_features[963] , \all_features[964] , \all_features[965] ,
    \all_features[966] , \all_features[967] , \all_features[968] ,
    \all_features[969] , \all_features[970] , \all_features[971] ,
    \all_features[972] , \all_features[973] , \all_features[974] ,
    \all_features[975] , \all_features[976] , \all_features[977] ,
    \all_features[978] , \all_features[979] , \all_features[980] ,
    \all_features[981] , \all_features[982] , \all_features[983] ,
    \all_features[984] , \all_features[985] , \all_features[986] ,
    \all_features[987] , \all_features[988] , \all_features[989] ,
    \all_features[990] , \all_features[991] , \all_features[992] ,
    \all_features[993] , \all_features[994] , \all_features[995] ,
    \all_features[996] , \all_features[997] , \all_features[998] ,
    \all_features[999] , \all_features[1000] , \all_features[1001] ,
    \all_features[1002] , \all_features[1003] , \all_features[1004] ,
    \all_features[1005] , \all_features[1006] , \all_features[1007] ,
    \all_features[1008] , \all_features[1009] , \all_features[1010] ,
    \all_features[1011] , \all_features[1012] , \all_features[1013] ,
    \all_features[1014] , \all_features[1015] , \all_features[1016] ,
    \all_features[1017] , \all_features[1018] , \all_features[1019] ,
    \all_features[1020] , \all_features[1021] , \all_features[1022] ,
    \all_features[1023] , \all_features[1024] , \all_features[1025] ,
    \all_features[1026] , \all_features[1027] , \all_features[1028] ,
    \all_features[1029] , \all_features[1030] , \all_features[1031] ,
    \all_features[1032] , \all_features[1033] , \all_features[1034] ,
    \all_features[1035] , \all_features[1036] , \all_features[1037] ,
    \all_features[1038] , \all_features[1039] , \all_features[1040] ,
    \all_features[1041] , \all_features[1042] , \all_features[1043] ,
    \all_features[1044] , \all_features[1045] , \all_features[1046] ,
    \all_features[1047] , \all_features[1048] , \all_features[1049] ,
    \all_features[1050] , \all_features[1051] , \all_features[1052] ,
    \all_features[1053] , \all_features[1054] , \all_features[1055] ,
    \all_features[1056] , \all_features[1057] , \all_features[1058] ,
    \all_features[1059] , \all_features[1060] , \all_features[1061] ,
    \all_features[1062] , \all_features[1063] , \all_features[1064] ,
    \all_features[1065] , \all_features[1066] , \all_features[1067] ,
    \all_features[1068] , \all_features[1069] , \all_features[1070] ,
    \all_features[1071] , \all_features[1072] , \all_features[1073] ,
    \all_features[1074] , \all_features[1075] , \all_features[1076] ,
    \all_features[1077] , \all_features[1078] , \all_features[1079] ,
    \all_features[1080] , \all_features[1081] , \all_features[1082] ,
    \all_features[1083] , \all_features[1084] , \all_features[1085] ,
    \all_features[1086] , \all_features[1087] , \all_features[1088] ,
    \all_features[1089] , \all_features[1090] , \all_features[1091] ,
    \all_features[1092] , \all_features[1093] , \all_features[1094] ,
    \all_features[1095] , \all_features[1096] , \all_features[1097] ,
    \all_features[1098] , \all_features[1099] , \all_features[1100] ,
    \all_features[1101] , \all_features[1102] , \all_features[1103] ,
    \all_features[1104] , \all_features[1105] , \all_features[1106] ,
    \all_features[1107] , \all_features[1108] , \all_features[1109] ,
    \all_features[1110] , \all_features[1111] , \all_features[1112] ,
    \all_features[1113] , \all_features[1114] , \all_features[1115] ,
    \all_features[1116] , \all_features[1117] , \all_features[1118] ,
    \all_features[1119] , \all_features[1120] , \all_features[1121] ,
    \all_features[1122] , \all_features[1123] , \all_features[1124] ,
    \all_features[1125] , \all_features[1126] , \all_features[1127] ,
    \all_features[1128] , \all_features[1129] , \all_features[1130] ,
    \all_features[1131] , \all_features[1132] , \all_features[1133] ,
    \all_features[1134] , \all_features[1135] , \all_features[1136] ,
    \all_features[1137] , \all_features[1138] , \all_features[1139] ,
    \all_features[1140] , \all_features[1141] , \all_features[1142] ,
    \all_features[1143] , \all_features[1144] , \all_features[1145] ,
    \all_features[1146] , \all_features[1147] , \all_features[1148] ,
    \all_features[1149] , \all_features[1150] , \all_features[1151] ,
    \all_features[1152] , \all_features[1153] , \all_features[1154] ,
    \all_features[1155] , \all_features[1156] , \all_features[1157] ,
    \all_features[1158] , \all_features[1159] , \all_features[1160] ,
    \all_features[1161] , \all_features[1162] , \all_features[1163] ,
    \all_features[1164] , \all_features[1165] , \all_features[1166] ,
    \all_features[1167] , \all_features[1168] , \all_features[1169] ,
    \all_features[1170] , \all_features[1171] , \all_features[1172] ,
    \all_features[1173] , \all_features[1174] , \all_features[1175] ,
    \all_features[1176] , \all_features[1177] , \all_features[1178] ,
    \all_features[1179] , \all_features[1180] , \all_features[1181] ,
    \all_features[1182] , \all_features[1183] , \all_features[1184] ,
    \all_features[1185] , \all_features[1186] , \all_features[1187] ,
    \all_features[1188] , \all_features[1189] , \all_features[1190] ,
    \all_features[1191] , \all_features[1192] , \all_features[1193] ,
    \all_features[1194] , \all_features[1195] , \all_features[1196] ,
    \all_features[1197] , \all_features[1198] , \all_features[1199] ,
    \all_features[1200] , \all_features[1201] , \all_features[1202] ,
    \all_features[1203] , \all_features[1204] , \all_features[1205] ,
    \all_features[1206] , \all_features[1207] , \all_features[1208] ,
    \all_features[1209] , \all_features[1210] , \all_features[1211] ,
    \all_features[1212] , \all_features[1213] , \all_features[1214] ,
    \all_features[1215] , \all_features[1216] , \all_features[1217] ,
    \all_features[1218] , \all_features[1219] , \all_features[1220] ,
    \all_features[1221] , \all_features[1222] , \all_features[1223] ,
    \all_features[1224] , \all_features[1225] , \all_features[1226] ,
    \all_features[1227] , \all_features[1228] , \all_features[1229] ,
    \all_features[1230] , \all_features[1231] , \all_features[1232] ,
    \all_features[1233] , \all_features[1234] , \all_features[1235] ,
    \all_features[1236] , \all_features[1237] , \all_features[1238] ,
    \all_features[1239] , \all_features[1240] , \all_features[1241] ,
    \all_features[1242] , \all_features[1243] , \all_features[1244] ,
    \all_features[1245] , \all_features[1246] , \all_features[1247] ,
    \all_features[1248] , \all_features[1249] , \all_features[1250] ,
    \all_features[1251] , \all_features[1252] , \all_features[1253] ,
    \all_features[1254] , \all_features[1255] , \all_features[1256] ,
    \all_features[1257] , \all_features[1258] , \all_features[1259] ,
    \all_features[1260] , \all_features[1261] , \all_features[1262] ,
    \all_features[1263] , \all_features[1264] , \all_features[1265] ,
    \all_features[1266] , \all_features[1267] , \all_features[1268] ,
    \all_features[1269] , \all_features[1270] , \all_features[1271] ,
    \all_features[1272] , \all_features[1273] , \all_features[1274] ,
    \all_features[1275] , \all_features[1276] , \all_features[1277] ,
    \all_features[1278] , \all_features[1279] , \all_features[1280] ,
    \all_features[1281] , \all_features[1282] , \all_features[1283] ,
    \all_features[1284] , \all_features[1285] , \all_features[1286] ,
    \all_features[1287] , \all_features[1288] , \all_features[1289] ,
    \all_features[1290] , \all_features[1291] , \all_features[1292] ,
    \all_features[1293] , \all_features[1294] , \all_features[1295] ,
    \all_features[1296] , \all_features[1297] , \all_features[1298] ,
    \all_features[1299] , \all_features[1300] , \all_features[1301] ,
    \all_features[1302] , \all_features[1303] , \all_features[1304] ,
    \all_features[1305] , \all_features[1306] , \all_features[1307] ,
    \all_features[1308] , \all_features[1309] , \all_features[1310] ,
    \all_features[1311] , \all_features[1312] , \all_features[1313] ,
    \all_features[1314] , \all_features[1315] , \all_features[1316] ,
    \all_features[1317] , \all_features[1318] , \all_features[1319] ,
    \all_features[1320] , \all_features[1321] , \all_features[1322] ,
    \all_features[1323] , \all_features[1324] , \all_features[1325] ,
    \all_features[1326] , \all_features[1327] , \all_features[1328] ,
    \all_features[1329] , \all_features[1330] , \all_features[1331] ,
    \all_features[1332] , \all_features[1333] , \all_features[1334] ,
    \all_features[1335] , \all_features[1336] , \all_features[1337] ,
    \all_features[1338] , \all_features[1339] , \all_features[1340] ,
    \all_features[1341] , \all_features[1342] , \all_features[1343] ,
    \all_features[1344] , \all_features[1345] , \all_features[1346] ,
    \all_features[1347] , \all_features[1348] , \all_features[1349] ,
    \all_features[1350] , \all_features[1351] , \all_features[1352] ,
    \all_features[1353] , \all_features[1354] , \all_features[1355] ,
    \all_features[1356] , \all_features[1357] , \all_features[1358] ,
    \all_features[1359] , \all_features[1360] , \all_features[1361] ,
    \all_features[1362] , \all_features[1363] , \all_features[1364] ,
    \all_features[1365] , \all_features[1366] , \all_features[1367] ,
    \all_features[1368] , \all_features[1369] , \all_features[1370] ,
    \all_features[1371] , \all_features[1372] , \all_features[1373] ,
    \all_features[1374] , \all_features[1375] , \all_features[1376] ,
    \all_features[1377] , \all_features[1378] , \all_features[1379] ,
    \all_features[1380] , \all_features[1381] , \all_features[1382] ,
    \all_features[1383] , \all_features[1384] , \all_features[1385] ,
    \all_features[1386] , \all_features[1387] , \all_features[1388] ,
    \all_features[1389] , \all_features[1390] , \all_features[1391] ,
    \all_features[1392] , \all_features[1393] , \all_features[1394] ,
    \all_features[1395] , \all_features[1396] , \all_features[1397] ,
    \all_features[1398] , \all_features[1399] , \all_features[1400] ,
    \all_features[1401] , \all_features[1402] , \all_features[1403] ,
    \all_features[1404] , \all_features[1405] , \all_features[1406] ,
    \all_features[1407] , \all_features[1408] , \all_features[1409] ,
    \all_features[1410] , \all_features[1411] , \all_features[1412] ,
    \all_features[1413] , \all_features[1414] , \all_features[1415] ,
    \all_features[1416] , \all_features[1417] , \all_features[1418] ,
    \all_features[1419] , \all_features[1420] , \all_features[1421] ,
    \all_features[1422] , \all_features[1423] , \all_features[1424] ,
    \all_features[1425] , \all_features[1426] , \all_features[1427] ,
    \all_features[1428] , \all_features[1429] , \all_features[1430] ,
    \all_features[1431] , \all_features[1432] , \all_features[1433] ,
    \all_features[1434] , \all_features[1435] , \all_features[1436] ,
    \all_features[1437] , \all_features[1438] , \all_features[1439] ,
    \all_features[1440] , \all_features[1441] , \all_features[1442] ,
    \all_features[1443] , \all_features[1444] , \all_features[1445] ,
    \all_features[1446] , \all_features[1447] , \all_features[1448] ,
    \all_features[1449] , \all_features[1450] , \all_features[1451] ,
    \all_features[1452] , \all_features[1453] , \all_features[1454] ,
    \all_features[1455] , \all_features[1456] , \all_features[1457] ,
    \all_features[1458] , \all_features[1459] , \all_features[1460] ,
    \all_features[1461] , \all_features[1462] , \all_features[1463] ,
    \all_features[1464] , \all_features[1465] , \all_features[1466] ,
    \all_features[1467] , \all_features[1468] , \all_features[1469] ,
    \all_features[1470] , \all_features[1471] , \all_features[1472] ,
    \all_features[1473] , \all_features[1474] , \all_features[1475] ,
    \all_features[1476] , \all_features[1477] , \all_features[1478] ,
    \all_features[1479] , \all_features[1480] , \all_features[1481] ,
    \all_features[1482] , \all_features[1483] , \all_features[1484] ,
    \all_features[1485] , \all_features[1486] , \all_features[1487] ,
    \all_features[1488] , \all_features[1489] , \all_features[1490] ,
    \all_features[1491] , \all_features[1492] , \all_features[1493] ,
    \all_features[1494] , \all_features[1495] , \all_features[1496] ,
    \all_features[1497] , \all_features[1498] , \all_features[1499] ,
    \all_features[1500] , \all_features[1501] , \all_features[1502] ,
    \all_features[1503] , \all_features[1504] , \all_features[1505] ,
    \all_features[1506] , \all_features[1507] , \all_features[1508] ,
    \all_features[1509] , \all_features[1510] , \all_features[1511] ,
    \all_features[1512] , \all_features[1513] , \all_features[1514] ,
    \all_features[1515] , \all_features[1516] , \all_features[1517] ,
    \all_features[1518] , \all_features[1519] , \all_features[1520] ,
    \all_features[1521] , \all_features[1522] , \all_features[1523] ,
    \all_features[1524] , \all_features[1525] , \all_features[1526] ,
    \all_features[1527] , \all_features[1528] , \all_features[1529] ,
    \all_features[1530] , \all_features[1531] , \all_features[1532] ,
    \all_features[1533] , \all_features[1534] , \all_features[1535] ,
    \all_features[1536] , \all_features[1537] , \all_features[1538] ,
    \all_features[1539] , \all_features[1540] , \all_features[1541] ,
    \all_features[1542] , \all_features[1543] , \all_features[1544] ,
    \all_features[1545] , \all_features[1546] , \all_features[1547] ,
    \all_features[1548] , \all_features[1549] , \all_features[1550] ,
    \all_features[1551] , \all_features[1552] , \all_features[1553] ,
    \all_features[1554] , \all_features[1555] , \all_features[1556] ,
    \all_features[1557] , \all_features[1558] , \all_features[1559] ,
    \all_features[1560] , \all_features[1561] , \all_features[1562] ,
    \all_features[1563] , \all_features[1564] , \all_features[1565] ,
    \all_features[1566] , \all_features[1567] , \all_features[1568] ,
    \all_features[1569] , \all_features[1570] , \all_features[1571] ,
    \all_features[1572] , \all_features[1573] , \all_features[1574] ,
    \all_features[1575] , \all_features[1576] , \all_features[1577] ,
    \all_features[1578] , \all_features[1579] , \all_features[1580] ,
    \all_features[1581] , \all_features[1582] , \all_features[1583] ,
    \all_features[1584] , \all_features[1585] , \all_features[1586] ,
    \all_features[1587] , \all_features[1588] , \all_features[1589] ,
    \all_features[1590] , \all_features[1591] , \all_features[1592] ,
    \all_features[1593] , \all_features[1594] , \all_features[1595] ,
    \all_features[1596] , \all_features[1597] , \all_features[1598] ,
    \all_features[1599] , \all_features[1600] , \all_features[1601] ,
    \all_features[1602] , \all_features[1603] , \all_features[1604] ,
    \all_features[1605] , \all_features[1606] , \all_features[1607] ,
    \all_features[1608] , \all_features[1609] , \all_features[1610] ,
    \all_features[1611] , \all_features[1612] , \all_features[1613] ,
    \all_features[1614] , \all_features[1615] , \all_features[1616] ,
    \all_features[1617] , \all_features[1618] , \all_features[1619] ,
    \all_features[1620] , \all_features[1621] , \all_features[1622] ,
    \all_features[1623] , \all_features[1624] , \all_features[1625] ,
    \all_features[1626] , \all_features[1627] , \all_features[1628] ,
    \all_features[1629] , \all_features[1630] , \all_features[1631] ,
    \all_features[1632] , \all_features[1633] , \all_features[1634] ,
    \all_features[1635] , \all_features[1636] , \all_features[1637] ,
    \all_features[1638] , \all_features[1639] , \all_features[1640] ,
    \all_features[1641] , \all_features[1642] , \all_features[1643] ,
    \all_features[1644] , \all_features[1645] , \all_features[1646] ,
    \all_features[1647] , \all_features[1648] , \all_features[1649] ,
    \all_features[1650] , \all_features[1651] , \all_features[1652] ,
    \all_features[1653] , \all_features[1654] , \all_features[1655] ,
    \all_features[1656] , \all_features[1657] , \all_features[1658] ,
    \all_features[1659] , \all_features[1660] , \all_features[1661] ,
    \all_features[1662] , \all_features[1663] , \all_features[1664] ,
    \all_features[1665] , \all_features[1666] , \all_features[1667] ,
    \all_features[1668] , \all_features[1669] , \all_features[1670] ,
    \all_features[1671] , \all_features[1672] , \all_features[1673] ,
    \all_features[1674] , \all_features[1675] , \all_features[1676] ,
    \all_features[1677] , \all_features[1678] , \all_features[1679] ,
    \all_features[1680] , \all_features[1681] , \all_features[1682] ,
    \all_features[1683] , \all_features[1684] , \all_features[1685] ,
    \all_features[1686] , \all_features[1687] , \all_features[1688] ,
    \all_features[1689] , \all_features[1690] , \all_features[1691] ,
    \all_features[1692] , \all_features[1693] , \all_features[1694] ,
    \all_features[1695] , \all_features[1696] , \all_features[1697] ,
    \all_features[1698] , \all_features[1699] , \all_features[1700] ,
    \all_features[1701] , \all_features[1702] , \all_features[1703] ,
    \all_features[1704] , \all_features[1705] , \all_features[1706] ,
    \all_features[1707] , \all_features[1708] , \all_features[1709] ,
    \all_features[1710] , \all_features[1711] , \all_features[1712] ,
    \all_features[1713] , \all_features[1714] , \all_features[1715] ,
    \all_features[1716] , \all_features[1717] , \all_features[1718] ,
    \all_features[1719] , \all_features[1720] , \all_features[1721] ,
    \all_features[1722] , \all_features[1723] , \all_features[1724] ,
    \all_features[1725] , \all_features[1726] , \all_features[1727] ,
    \all_features[1728] , \all_features[1729] , \all_features[1730] ,
    \all_features[1731] , \all_features[1732] , \all_features[1733] ,
    \all_features[1734] , \all_features[1735] , \all_features[1736] ,
    \all_features[1737] , \all_features[1738] , \all_features[1739] ,
    \all_features[1740] , \all_features[1741] , \all_features[1742] ,
    \all_features[1743] , \all_features[1744] , \all_features[1745] ,
    \all_features[1746] , \all_features[1747] , \all_features[1748] ,
    \all_features[1749] , \all_features[1750] , \all_features[1751] ,
    \all_features[1752] , \all_features[1753] , \all_features[1754] ,
    \all_features[1755] , \all_features[1756] , \all_features[1757] ,
    \all_features[1758] , \all_features[1759] , \all_features[1760] ,
    \all_features[1761] , \all_features[1762] , \all_features[1763] ,
    \all_features[1764] , \all_features[1765] , \all_features[1766] ,
    \all_features[1767] , \all_features[1768] , \all_features[1769] ,
    \all_features[1770] , \all_features[1771] , \all_features[1772] ,
    \all_features[1773] , \all_features[1774] , \all_features[1775] ,
    \all_features[1776] , \all_features[1777] , \all_features[1778] ,
    \all_features[1779] , \all_features[1780] , \all_features[1781] ,
    \all_features[1782] , \all_features[1783] , \all_features[1784] ,
    \all_features[1785] , \all_features[1786] , \all_features[1787] ,
    \all_features[1788] , \all_features[1789] , \all_features[1790] ,
    \all_features[1791] , \all_features[1792] , \all_features[1793] ,
    \all_features[1794] , \all_features[1795] , \all_features[1796] ,
    \all_features[1797] , \all_features[1798] , \all_features[1799] ,
    \all_features[1800] , \all_features[1801] , \all_features[1802] ,
    \all_features[1803] , \all_features[1804] , \all_features[1805] ,
    \all_features[1806] , \all_features[1807] , \all_features[1808] ,
    \all_features[1809] , \all_features[1810] , \all_features[1811] ,
    \all_features[1812] , \all_features[1813] , \all_features[1814] ,
    \all_features[1815] , \all_features[1816] , \all_features[1817] ,
    \all_features[1818] , \all_features[1819] , \all_features[1820] ,
    \all_features[1821] , \all_features[1822] , \all_features[1823] ,
    \all_features[1824] , \all_features[1825] , \all_features[1826] ,
    \all_features[1827] , \all_features[1828] , \all_features[1829] ,
    \all_features[1830] , \all_features[1831] , \all_features[1832] ,
    \all_features[1833] , \all_features[1834] , \all_features[1835] ,
    \all_features[1836] , \all_features[1837] , \all_features[1838] ,
    \all_features[1839] , \all_features[1840] , \all_features[1841] ,
    \all_features[1842] , \all_features[1843] , \all_features[1844] ,
    \all_features[1845] , \all_features[1846] , \all_features[1847] ,
    \all_features[1848] , \all_features[1849] , \all_features[1850] ,
    \all_features[1851] , \all_features[1852] , \all_features[1853] ,
    \all_features[1854] , \all_features[1855] , \all_features[1856] ,
    \all_features[1857] , \all_features[1858] , \all_features[1859] ,
    \all_features[1860] , \all_features[1861] , \all_features[1862] ,
    \all_features[1863] , \all_features[1864] , \all_features[1865] ,
    \all_features[1866] , \all_features[1867] , \all_features[1868] ,
    \all_features[1869] , \all_features[1870] , \all_features[1871] ,
    \all_features[1872] , \all_features[1873] , \all_features[1874] ,
    \all_features[1875] , \all_features[1876] , \all_features[1877] ,
    \all_features[1878] , \all_features[1879] , \all_features[1880] ,
    \all_features[1881] , \all_features[1882] , \all_features[1883] ,
    \all_features[1884] , \all_features[1885] , \all_features[1886] ,
    \all_features[1887] , \all_features[1888] , \all_features[1889] ,
    \all_features[1890] , \all_features[1891] , \all_features[1892] ,
    \all_features[1893] , \all_features[1894] , \all_features[1895] ,
    \all_features[1896] , \all_features[1897] , \all_features[1898] ,
    \all_features[1899] , \all_features[1900] , \all_features[1901] ,
    \all_features[1902] , \all_features[1903] , \all_features[1904] ,
    \all_features[1905] , \all_features[1906] , \all_features[1907] ,
    \all_features[1908] , \all_features[1909] , \all_features[1910] ,
    \all_features[1911] , \all_features[1912] , \all_features[1913] ,
    \all_features[1914] , \all_features[1915] , \all_features[1916] ,
    \all_features[1917] , \all_features[1918] , \all_features[1919] ,
    \all_features[1920] , \all_features[1921] , \all_features[1922] ,
    \all_features[1923] , \all_features[1924] , \all_features[1925] ,
    \all_features[1926] , \all_features[1927] , \all_features[1928] ,
    \all_features[1929] , \all_features[1930] , \all_features[1931] ,
    \all_features[1932] , \all_features[1933] , \all_features[1934] ,
    \all_features[1935] , \all_features[1936] , \all_features[1937] ,
    \all_features[1938] , \all_features[1939] , \all_features[1940] ,
    \all_features[1941] , \all_features[1942] , \all_features[1943] ,
    \all_features[1944] , \all_features[1945] , \all_features[1946] ,
    \all_features[1947] , \all_features[1948] , \all_features[1949] ,
    \all_features[1950] , \all_features[1951] , \all_features[1952] ,
    \all_features[1953] , \all_features[1954] , \all_features[1955] ,
    \all_features[1956] , \all_features[1957] , \all_features[1958] ,
    \all_features[1959] , \all_features[1960] , \all_features[1961] ,
    \all_features[1962] , \all_features[1963] , \all_features[1964] ,
    \all_features[1965] , \all_features[1966] , \all_features[1967] ,
    \all_features[1968] , \all_features[1969] , \all_features[1970] ,
    \all_features[1971] , \all_features[1972] , \all_features[1973] ,
    \all_features[1974] , \all_features[1975] , \all_features[1976] ,
    \all_features[1977] , \all_features[1978] , \all_features[1979] ,
    \all_features[1980] , \all_features[1981] , \all_features[1982] ,
    \all_features[1983] , \all_features[1984] , \all_features[1985] ,
    \all_features[1986] , \all_features[1987] , \all_features[1988] ,
    \all_features[1989] , \all_features[1990] , \all_features[1991] ,
    \all_features[1992] , \all_features[1993] , \all_features[1994] ,
    \all_features[1995] , \all_features[1996] , \all_features[1997] ,
    \all_features[1998] , \all_features[1999] , \all_features[2000] ,
    \all_features[2001] , \all_features[2002] , \all_features[2003] ,
    \all_features[2004] , \all_features[2005] , \all_features[2006] ,
    \all_features[2007] , \all_features[2008] , \all_features[2009] ,
    \all_features[2010] , \all_features[2011] , \all_features[2012] ,
    \all_features[2013] , \all_features[2014] , \all_features[2015] ,
    \all_features[2016] , \all_features[2017] , \all_features[2018] ,
    \all_features[2019] , \all_features[2020] , \all_features[2021] ,
    \all_features[2022] , \all_features[2023] , \all_features[2024] ,
    \all_features[2025] , \all_features[2026] , \all_features[2027] ,
    \all_features[2028] , \all_features[2029] , \all_features[2030] ,
    \all_features[2031] , \all_features[2032] , \all_features[2033] ,
    \all_features[2034] , \all_features[2035] , \all_features[2036] ,
    \all_features[2037] , \all_features[2038] , \all_features[2039] ,
    \all_features[2040] , \all_features[2041] , \all_features[2042] ,
    \all_features[2043] , \all_features[2044] , \all_features[2045] ,
    \all_features[2046] , \all_features[2047] , \all_features[2048] ,
    \all_features[2049] , \all_features[2050] , \all_features[2051] ,
    \all_features[2052] , \all_features[2053] , \all_features[2054] ,
    \all_features[2055] , \all_features[2056] , \all_features[2057] ,
    \all_features[2058] , \all_features[2059] , \all_features[2060] ,
    \all_features[2061] , \all_features[2062] , \all_features[2063] ,
    \all_features[2064] , \all_features[2065] , \all_features[2066] ,
    \all_features[2067] , \all_features[2068] , \all_features[2069] ,
    \all_features[2070] , \all_features[2071] , \all_features[2072] ,
    \all_features[2073] , \all_features[2074] , \all_features[2075] ,
    \all_features[2076] , \all_features[2077] , \all_features[2078] ,
    \all_features[2079] , \all_features[2080] , \all_features[2081] ,
    \all_features[2082] , \all_features[2083] , \all_features[2084] ,
    \all_features[2085] , \all_features[2086] , \all_features[2087] ,
    \all_features[2088] , \all_features[2089] , \all_features[2090] ,
    \all_features[2091] , \all_features[2092] , \all_features[2093] ,
    \all_features[2094] , \all_features[2095] , \all_features[2096] ,
    \all_features[2097] , \all_features[2098] , \all_features[2099] ,
    \all_features[2100] , \all_features[2101] , \all_features[2102] ,
    \all_features[2103] , \all_features[2104] , \all_features[2105] ,
    \all_features[2106] , \all_features[2107] , \all_features[2108] ,
    \all_features[2109] , \all_features[2110] , \all_features[2111] ,
    \all_features[2112] , \all_features[2113] , \all_features[2114] ,
    \all_features[2115] , \all_features[2116] , \all_features[2117] ,
    \all_features[2118] , \all_features[2119] , \all_features[2120] ,
    \all_features[2121] , \all_features[2122] , \all_features[2123] ,
    \all_features[2124] , \all_features[2125] , \all_features[2126] ,
    \all_features[2127] , \all_features[2128] , \all_features[2129] ,
    \all_features[2130] , \all_features[2131] , \all_features[2132] ,
    \all_features[2133] , \all_features[2134] , \all_features[2135] ,
    \all_features[2136] , \all_features[2137] , \all_features[2138] ,
    \all_features[2139] , \all_features[2140] , \all_features[2141] ,
    \all_features[2142] , \all_features[2143] , \all_features[2144] ,
    \all_features[2145] , \all_features[2146] , \all_features[2147] ,
    \all_features[2148] , \all_features[2149] , \all_features[2150] ,
    \all_features[2151] , \all_features[2152] , \all_features[2153] ,
    \all_features[2154] , \all_features[2155] , \all_features[2156] ,
    \all_features[2157] , \all_features[2158] , \all_features[2159] ,
    \all_features[2160] , \all_features[2161] , \all_features[2162] ,
    \all_features[2163] , \all_features[2164] , \all_features[2165] ,
    \all_features[2166] , \all_features[2167] , \all_features[2168] ,
    \all_features[2169] , \all_features[2170] , \all_features[2171] ,
    \all_features[2172] , \all_features[2173] , \all_features[2174] ,
    \all_features[2175] , \all_features[2176] , \all_features[2177] ,
    \all_features[2178] , \all_features[2179] , \all_features[2180] ,
    \all_features[2181] , \all_features[2182] , \all_features[2183] ,
    \all_features[2184] , \all_features[2185] , \all_features[2186] ,
    \all_features[2187] , \all_features[2188] , \all_features[2189] ,
    \all_features[2190] , \all_features[2191] , \all_features[2192] ,
    \all_features[2193] , \all_features[2194] , \all_features[2195] ,
    \all_features[2196] , \all_features[2197] , \all_features[2198] ,
    \all_features[2199] , \all_features[2200] , \all_features[2201] ,
    \all_features[2202] , \all_features[2203] , \all_features[2204] ,
    \all_features[2205] , \all_features[2206] , \all_features[2207] ,
    \all_features[2208] , \all_features[2209] , \all_features[2210] ,
    \all_features[2211] , \all_features[2212] , \all_features[2213] ,
    \all_features[2214] , \all_features[2215] , \all_features[2216] ,
    \all_features[2217] , \all_features[2218] , \all_features[2219] ,
    \all_features[2220] , \all_features[2221] , \all_features[2222] ,
    \all_features[2223] , \all_features[2224] , \all_features[2225] ,
    \all_features[2226] , \all_features[2227] , \all_features[2228] ,
    \all_features[2229] , \all_features[2230] , \all_features[2231] ,
    \all_features[2232] , \all_features[2233] , \all_features[2234] ,
    \all_features[2235] , \all_features[2236] , \all_features[2237] ,
    \all_features[2238] , \all_features[2239] , \all_features[2240] ,
    \all_features[2241] , \all_features[2242] , \all_features[2243] ,
    \all_features[2244] , \all_features[2245] , \all_features[2246] ,
    \all_features[2247] , \all_features[2248] , \all_features[2249] ,
    \all_features[2250] , \all_features[2251] , \all_features[2252] ,
    \all_features[2253] , \all_features[2254] , \all_features[2255] ,
    \all_features[2256] , \all_features[2257] , \all_features[2258] ,
    \all_features[2259] , \all_features[2260] , \all_features[2261] ,
    \all_features[2262] , \all_features[2263] , \all_features[2264] ,
    \all_features[2265] , \all_features[2266] , \all_features[2267] ,
    \all_features[2268] , \all_features[2269] , \all_features[2270] ,
    \all_features[2271] , \all_features[2272] , \all_features[2273] ,
    \all_features[2274] , \all_features[2275] , \all_features[2276] ,
    \all_features[2277] , \all_features[2278] , \all_features[2279] ,
    \all_features[2280] , \all_features[2281] , \all_features[2282] ,
    \all_features[2283] , \all_features[2284] , \all_features[2285] ,
    \all_features[2286] , \all_features[2287] , \all_features[2288] ,
    \all_features[2289] , \all_features[2290] , \all_features[2291] ,
    \all_features[2292] , \all_features[2293] , \all_features[2294] ,
    \all_features[2295] , \all_features[2296] , \all_features[2297] ,
    \all_features[2298] , \all_features[2299] , \all_features[2300] ,
    \all_features[2301] , \all_features[2302] , \all_features[2303] ,
    \all_features[2304] , \all_features[2305] , \all_features[2306] ,
    \all_features[2307] , \all_features[2308] , \all_features[2309] ,
    \all_features[2310] , \all_features[2311] , \all_features[2312] ,
    \all_features[2313] , \all_features[2314] , \all_features[2315] ,
    \all_features[2316] , \all_features[2317] , \all_features[2318] ,
    \all_features[2319] , \all_features[2320] , \all_features[2321] ,
    \all_features[2322] , \all_features[2323] , \all_features[2324] ,
    \all_features[2325] , \all_features[2326] , \all_features[2327] ,
    \all_features[2328] , \all_features[2329] , \all_features[2330] ,
    \all_features[2331] , \all_features[2332] , \all_features[2333] ,
    \all_features[2334] , \all_features[2335] , \all_features[2336] ,
    \all_features[2337] , \all_features[2338] , \all_features[2339] ,
    \all_features[2340] , \all_features[2341] , \all_features[2342] ,
    \all_features[2343] , \all_features[2344] , \all_features[2345] ,
    \all_features[2346] , \all_features[2347] , \all_features[2348] ,
    \all_features[2349] , \all_features[2350] , \all_features[2351] ,
    \all_features[2352] , \all_features[2353] , \all_features[2354] ,
    \all_features[2355] , \all_features[2356] , \all_features[2357] ,
    \all_features[2358] , \all_features[2359] , \all_features[2360] ,
    \all_features[2361] , \all_features[2362] , \all_features[2363] ,
    \all_features[2364] , \all_features[2365] , \all_features[2366] ,
    \all_features[2367] , \all_features[2368] , \all_features[2369] ,
    \all_features[2370] , \all_features[2371] , \all_features[2372] ,
    \all_features[2373] , \all_features[2374] , \all_features[2375] ,
    \all_features[2376] , \all_features[2377] , \all_features[2378] ,
    \all_features[2379] , \all_features[2380] , \all_features[2381] ,
    \all_features[2382] , \all_features[2383] , \all_features[2384] ,
    \all_features[2385] , \all_features[2386] , \all_features[2387] ,
    \all_features[2388] , \all_features[2389] , \all_features[2390] ,
    \all_features[2391] , \all_features[2392] , \all_features[2393] ,
    \all_features[2394] , \all_features[2395] , \all_features[2396] ,
    \all_features[2397] , \all_features[2398] , \all_features[2399] ,
    \all_features[2400] , \all_features[2401] , \all_features[2402] ,
    \all_features[2403] , \all_features[2404] , \all_features[2405] ,
    \all_features[2406] , \all_features[2407] , \all_features[2408] ,
    \all_features[2409] , \all_features[2410] , \all_features[2411] ,
    \all_features[2412] , \all_features[2413] , \all_features[2414] ,
    \all_features[2415] , \all_features[2416] , \all_features[2417] ,
    \all_features[2418] , \all_features[2419] , \all_features[2420] ,
    \all_features[2421] , \all_features[2422] , \all_features[2423] ,
    \all_features[2424] , \all_features[2425] , \all_features[2426] ,
    \all_features[2427] , \all_features[2428] , \all_features[2429] ,
    \all_features[2430] , \all_features[2431] , \all_features[2432] ,
    \all_features[2433] , \all_features[2434] , \all_features[2435] ,
    \all_features[2436] , \all_features[2437] , \all_features[2438] ,
    \all_features[2439] , \all_features[2440] , \all_features[2441] ,
    \all_features[2442] , \all_features[2443] , \all_features[2444] ,
    \all_features[2445] , \all_features[2446] , \all_features[2447] ,
    \all_features[2448] , \all_features[2449] , \all_features[2450] ,
    \all_features[2451] , \all_features[2452] , \all_features[2453] ,
    \all_features[2454] , \all_features[2455] , \all_features[2456] ,
    \all_features[2457] , \all_features[2458] , \all_features[2459] ,
    \all_features[2460] , \all_features[2461] , \all_features[2462] ,
    \all_features[2463] , \all_features[2464] , \all_features[2465] ,
    \all_features[2466] , \all_features[2467] , \all_features[2468] ,
    \all_features[2469] , \all_features[2470] , \all_features[2471] ,
    \all_features[2472] , \all_features[2473] , \all_features[2474] ,
    \all_features[2475] , \all_features[2476] , \all_features[2477] ,
    \all_features[2478] , \all_features[2479] , \all_features[2480] ,
    \all_features[2481] , \all_features[2482] , \all_features[2483] ,
    \all_features[2484] , \all_features[2485] , \all_features[2486] ,
    \all_features[2487] , \all_features[2488] , \all_features[2489] ,
    \all_features[2490] , \all_features[2491] , \all_features[2492] ,
    \all_features[2493] , \all_features[2494] , \all_features[2495] ,
    \all_features[2496] , \all_features[2497] , \all_features[2498] ,
    \all_features[2499] , \all_features[2500] , \all_features[2501] ,
    \all_features[2502] , \all_features[2503] , \all_features[2504] ,
    \all_features[2505] , \all_features[2506] , \all_features[2507] ,
    \all_features[2508] , \all_features[2509] , \all_features[2510] ,
    \all_features[2511] , \all_features[2512] , \all_features[2513] ,
    \all_features[2514] , \all_features[2515] , \all_features[2516] ,
    \all_features[2517] , \all_features[2518] , \all_features[2519] ,
    \all_features[2520] , \all_features[2521] , \all_features[2522] ,
    \all_features[2523] , \all_features[2524] , \all_features[2525] ,
    \all_features[2526] , \all_features[2527] , \all_features[2528] ,
    \all_features[2529] , \all_features[2530] , \all_features[2531] ,
    \all_features[2532] , \all_features[2533] , \all_features[2534] ,
    \all_features[2535] , \all_features[2536] , \all_features[2537] ,
    \all_features[2538] , \all_features[2539] , \all_features[2540] ,
    \all_features[2541] , \all_features[2542] , \all_features[2543] ,
    \all_features[2544] , \all_features[2545] , \all_features[2546] ,
    \all_features[2547] , \all_features[2548] , \all_features[2549] ,
    \all_features[2550] , \all_features[2551] , \all_features[2552] ,
    \all_features[2553] , \all_features[2554] , \all_features[2555] ,
    \all_features[2556] , \all_features[2557] , \all_features[2558] ,
    \all_features[2559] , \all_features[2560] , \all_features[2561] ,
    \all_features[2562] , \all_features[2563] , \all_features[2564] ,
    \all_features[2565] , \all_features[2566] , \all_features[2567] ,
    \all_features[2568] , \all_features[2569] , \all_features[2570] ,
    \all_features[2571] , \all_features[2572] , \all_features[2573] ,
    \all_features[2574] , \all_features[2575] , \all_features[2576] ,
    \all_features[2577] , \all_features[2578] , \all_features[2579] ,
    \all_features[2580] , \all_features[2581] , \all_features[2582] ,
    \all_features[2583] , \all_features[2584] , \all_features[2585] ,
    \all_features[2586] , \all_features[2587] , \all_features[2588] ,
    \all_features[2589] , \all_features[2590] , \all_features[2591] ,
    \all_features[2592] , \all_features[2593] , \all_features[2594] ,
    \all_features[2595] , \all_features[2596] , \all_features[2597] ,
    \all_features[2598] , \all_features[2599] , \all_features[2600] ,
    \all_features[2601] , \all_features[2602] , \all_features[2603] ,
    \all_features[2604] , \all_features[2605] , \all_features[2606] ,
    \all_features[2607] , \all_features[2608] , \all_features[2609] ,
    \all_features[2610] , \all_features[2611] , \all_features[2612] ,
    \all_features[2613] , \all_features[2614] , \all_features[2615] ,
    \all_features[2616] , \all_features[2617] , \all_features[2618] ,
    \all_features[2619] , \all_features[2620] , \all_features[2621] ,
    \all_features[2622] , \all_features[2623] , \all_features[2624] ,
    \all_features[2625] , \all_features[2626] , \all_features[2627] ,
    \all_features[2628] , \all_features[2629] , \all_features[2630] ,
    \all_features[2631] , \all_features[2632] , \all_features[2633] ,
    \all_features[2634] , \all_features[2635] , \all_features[2636] ,
    \all_features[2637] , \all_features[2638] , \all_features[2639] ,
    \all_features[2640] , \all_features[2641] , \all_features[2642] ,
    \all_features[2643] , \all_features[2644] , \all_features[2645] ,
    \all_features[2646] , \all_features[2647] , \all_features[2648] ,
    \all_features[2649] , \all_features[2650] , \all_features[2651] ,
    \all_features[2652] , \all_features[2653] , \all_features[2654] ,
    \all_features[2655] , \all_features[2656] , \all_features[2657] ,
    \all_features[2658] , \all_features[2659] , \all_features[2660] ,
    \all_features[2661] , \all_features[2662] , \all_features[2663] ,
    \all_features[2664] , \all_features[2665] , \all_features[2666] ,
    \all_features[2667] , \all_features[2668] , \all_features[2669] ,
    \all_features[2670] , \all_features[2671] , \all_features[2672] ,
    \all_features[2673] , \all_features[2674] , \all_features[2675] ,
    \all_features[2676] , \all_features[2677] , \all_features[2678] ,
    \all_features[2679] , \all_features[2680] , \all_features[2681] ,
    \all_features[2682] , \all_features[2683] , \all_features[2684] ,
    \all_features[2685] , \all_features[2686] , \all_features[2687] ,
    \all_features[2688] , \all_features[2689] , \all_features[2690] ,
    \all_features[2691] , \all_features[2692] , \all_features[2693] ,
    \all_features[2694] , \all_features[2695] , \all_features[2696] ,
    \all_features[2697] , \all_features[2698] , \all_features[2699] ,
    \all_features[2700] , \all_features[2701] , \all_features[2702] ,
    \all_features[2703] , \all_features[2704] , \all_features[2705] ,
    \all_features[2706] , \all_features[2707] , \all_features[2708] ,
    \all_features[2709] , \all_features[2710] , \all_features[2711] ,
    \all_features[2712] , \all_features[2713] , \all_features[2714] ,
    \all_features[2715] , \all_features[2716] , \all_features[2717] ,
    \all_features[2718] , \all_features[2719] , \all_features[2720] ,
    \all_features[2721] , \all_features[2722] , \all_features[2723] ,
    \all_features[2724] , \all_features[2725] , \all_features[2726] ,
    \all_features[2727] , \all_features[2728] , \all_features[2729] ,
    \all_features[2730] , \all_features[2731] , \all_features[2732] ,
    \all_features[2733] , \all_features[2734] , \all_features[2735] ,
    \all_features[2736] , \all_features[2737] , \all_features[2738] ,
    \all_features[2739] , \all_features[2740] , \all_features[2741] ,
    \all_features[2742] , \all_features[2743] , \all_features[2744] ,
    \all_features[2745] , \all_features[2746] , \all_features[2747] ,
    \all_features[2748] , \all_features[2749] , \all_features[2750] ,
    \all_features[2751] , \all_features[2752] , \all_features[2753] ,
    \all_features[2754] , \all_features[2755] , \all_features[2756] ,
    \all_features[2757] , \all_features[2758] , \all_features[2759] ,
    \all_features[2760] , \all_features[2761] , \all_features[2762] ,
    \all_features[2763] , \all_features[2764] , \all_features[2765] ,
    \all_features[2766] , \all_features[2767] , \all_features[2768] ,
    \all_features[2769] , \all_features[2770] , \all_features[2771] ,
    \all_features[2772] , \all_features[2773] , \all_features[2774] ,
    \all_features[2775] , \all_features[2776] , \all_features[2777] ,
    \all_features[2778] , \all_features[2779] , \all_features[2780] ,
    \all_features[2781] , \all_features[2782] , \all_features[2783] ,
    \all_features[2784] , \all_features[2785] , \all_features[2786] ,
    \all_features[2787] , \all_features[2788] , \all_features[2789] ,
    \all_features[2790] , \all_features[2791] , \all_features[2792] ,
    \all_features[2793] , \all_features[2794] , \all_features[2795] ,
    \all_features[2796] , \all_features[2797] , \all_features[2798] ,
    \all_features[2799] , \all_features[2800] , \all_features[2801] ,
    \all_features[2802] , \all_features[2803] , \all_features[2804] ,
    \all_features[2805] , \all_features[2806] , \all_features[2807] ,
    \all_features[2808] , \all_features[2809] , \all_features[2810] ,
    \all_features[2811] , \all_features[2812] , \all_features[2813] ,
    \all_features[2814] , \all_features[2815] , \all_features[2816] ,
    \all_features[2817] , \all_features[2818] , \all_features[2819] ,
    \all_features[2820] , \all_features[2821] , \all_features[2822] ,
    \all_features[2823] , \all_features[2824] , \all_features[2825] ,
    \all_features[2826] , \all_features[2827] , \all_features[2828] ,
    \all_features[2829] , \all_features[2830] , \all_features[2831] ,
    \all_features[2832] , \all_features[2833] , \all_features[2834] ,
    \all_features[2835] , \all_features[2836] , \all_features[2837] ,
    \all_features[2838] , \all_features[2839] , \all_features[2840] ,
    \all_features[2841] , \all_features[2842] , \all_features[2843] ,
    \all_features[2844] , \all_features[2845] , \all_features[2846] ,
    \all_features[2847] , \all_features[2848] , \all_features[2849] ,
    \all_features[2850] , \all_features[2851] , \all_features[2852] ,
    \all_features[2853] , \all_features[2854] , \all_features[2855] ,
    \all_features[2856] , \all_features[2857] , \all_features[2858] ,
    \all_features[2859] , \all_features[2860] , \all_features[2861] ,
    \all_features[2862] , \all_features[2863] , \all_features[2864] ,
    \all_features[2865] , \all_features[2866] , \all_features[2867] ,
    \all_features[2868] , \all_features[2869] , \all_features[2870] ,
    \all_features[2871] , \all_features[2872] , \all_features[2873] ,
    \all_features[2874] , \all_features[2875] , \all_features[2876] ,
    \all_features[2877] , \all_features[2878] , \all_features[2879] ,
    \all_features[2880] , \all_features[2881] , \all_features[2882] ,
    \all_features[2883] , \all_features[2884] , \all_features[2885] ,
    \all_features[2886] , \all_features[2887] , \all_features[2888] ,
    \all_features[2889] , \all_features[2890] , \all_features[2891] ,
    \all_features[2892] , \all_features[2893] , \all_features[2894] ,
    \all_features[2895] , \all_features[2896] , \all_features[2897] ,
    \all_features[2898] , \all_features[2899] , \all_features[2900] ,
    \all_features[2901] , \all_features[2902] , \all_features[2903] ,
    \all_features[2904] , \all_features[2905] , \all_features[2906] ,
    \all_features[2907] , \all_features[2908] , \all_features[2909] ,
    \all_features[2910] , \all_features[2911] , \all_features[2912] ,
    \all_features[2913] , \all_features[2914] , \all_features[2915] ,
    \all_features[2916] , \all_features[2917] , \all_features[2918] ,
    \all_features[2919] , \all_features[2920] , \all_features[2921] ,
    \all_features[2922] , \all_features[2923] , \all_features[2924] ,
    \all_features[2925] , \all_features[2926] , \all_features[2927] ,
    \all_features[2928] , \all_features[2929] , \all_features[2930] ,
    \all_features[2931] , \all_features[2932] , \all_features[2933] ,
    \all_features[2934] , \all_features[2935] , \all_features[2936] ,
    \all_features[2937] , \all_features[2938] , \all_features[2939] ,
    \all_features[2940] , \all_features[2941] , \all_features[2942] ,
    \all_features[2943] , \all_features[2944] , \all_features[2945] ,
    \all_features[2946] , \all_features[2947] , \all_features[2948] ,
    \all_features[2949] , \all_features[2950] , \all_features[2951] ,
    \all_features[2952] , \all_features[2953] , \all_features[2954] ,
    \all_features[2955] , \all_features[2956] , \all_features[2957] ,
    \all_features[2958] , \all_features[2959] , \all_features[2960] ,
    \all_features[2961] , \all_features[2962] , \all_features[2963] ,
    \all_features[2964] , \all_features[2965] , \all_features[2966] ,
    \all_features[2967] , \all_features[2968] , \all_features[2969] ,
    \all_features[2970] , \all_features[2971] , \all_features[2972] ,
    \all_features[2973] , \all_features[2974] , \all_features[2975] ,
    \all_features[2976] , \all_features[2977] , \all_features[2978] ,
    \all_features[2979] , \all_features[2980] , \all_features[2981] ,
    \all_features[2982] , \all_features[2983] , \all_features[2984] ,
    \all_features[2985] , \all_features[2986] , \all_features[2987] ,
    \all_features[2988] , \all_features[2989] , \all_features[2990] ,
    \all_features[2991] , \all_features[2992] , \all_features[2993] ,
    \all_features[2994] , \all_features[2995] , \all_features[2996] ,
    \all_features[2997] , \all_features[2998] , \all_features[2999] ,
    \all_features[3000] , \all_features[3001] , \all_features[3002] ,
    \all_features[3003] , \all_features[3004] , \all_features[3005] ,
    \all_features[3006] , \all_features[3007] , \all_features[3008] ,
    \all_features[3009] , \all_features[3010] , \all_features[3011] ,
    \all_features[3012] , \all_features[3013] , \all_features[3014] ,
    \all_features[3015] , \all_features[3016] , \all_features[3017] ,
    \all_features[3018] , \all_features[3019] , \all_features[3020] ,
    \all_features[3021] , \all_features[3022] , \all_features[3023] ,
    \all_features[3024] , \all_features[3025] , \all_features[3026] ,
    \all_features[3027] , \all_features[3028] , \all_features[3029] ,
    \all_features[3030] , \all_features[3031] , \all_features[3032] ,
    \all_features[3033] , \all_features[3034] , \all_features[3035] ,
    \all_features[3036] , \all_features[3037] , \all_features[3038] ,
    \all_features[3039] , \all_features[3040] , \all_features[3041] ,
    \all_features[3042] , \all_features[3043] , \all_features[3044] ,
    \all_features[3045] , \all_features[3046] , \all_features[3047] ,
    \all_features[3048] , \all_features[3049] , \all_features[3050] ,
    \all_features[3051] , \all_features[3052] , \all_features[3053] ,
    \all_features[3054] , \all_features[3055] , \all_features[3056] ,
    \all_features[3057] , \all_features[3058] , \all_features[3059] ,
    \all_features[3060] , \all_features[3061] , \all_features[3062] ,
    \all_features[3063] , \all_features[3064] , \all_features[3065] ,
    \all_features[3066] , \all_features[3067] , \all_features[3068] ,
    \all_features[3069] , \all_features[3070] , \all_features[3071] ,
    \all_features[3072] , \all_features[3073] , \all_features[3074] ,
    \all_features[3075] , \all_features[3076] , \all_features[3077] ,
    \all_features[3078] , \all_features[3079] , \all_features[3080] ,
    \all_features[3081] , \all_features[3082] , \all_features[3083] ,
    \all_features[3084] , \all_features[3085] , \all_features[3086] ,
    \all_features[3087] , \all_features[3088] , \all_features[3089] ,
    \all_features[3090] , \all_features[3091] , \all_features[3092] ,
    \all_features[3093] , \all_features[3094] , \all_features[3095] ,
    \all_features[3096] , \all_features[3097] , \all_features[3098] ,
    \all_features[3099] , \all_features[3100] , \all_features[3101] ,
    \all_features[3102] , \all_features[3103] , \all_features[3104] ,
    \all_features[3105] , \all_features[3106] , \all_features[3107] ,
    \all_features[3108] , \all_features[3109] , \all_features[3110] ,
    \all_features[3111] , \all_features[3112] , \all_features[3113] ,
    \all_features[3114] , \all_features[3115] , \all_features[3116] ,
    \all_features[3117] , \all_features[3118] , \all_features[3119] ,
    \all_features[3120] , \all_features[3121] , \all_features[3122] ,
    \all_features[3123] , \all_features[3124] , \all_features[3125] ,
    \all_features[3126] , \all_features[3127] , \all_features[3128] ,
    \all_features[3129] , \all_features[3130] , \all_features[3131] ,
    \all_features[3132] , \all_features[3133] , \all_features[3134] ,
    \all_features[3135] , \all_features[3136] , \all_features[3137] ,
    \all_features[3138] , \all_features[3139] , \all_features[3140] ,
    \all_features[3141] , \all_features[3142] , \all_features[3143] ,
    \all_features[3144] , \all_features[3145] , \all_features[3146] ,
    \all_features[3147] , \all_features[3148] , \all_features[3149] ,
    \all_features[3150] , \all_features[3151] , \all_features[3152] ,
    \all_features[3153] , \all_features[3154] , \all_features[3155] ,
    \all_features[3156] , \all_features[3157] , \all_features[3158] ,
    \all_features[3159] , \all_features[3160] , \all_features[3161] ,
    \all_features[3162] , \all_features[3163] , \all_features[3164] ,
    \all_features[3165] , \all_features[3166] , \all_features[3167] ,
    \all_features[3168] , \all_features[3169] , \all_features[3170] ,
    \all_features[3171] , \all_features[3172] , \all_features[3173] ,
    \all_features[3174] , \all_features[3175] , \all_features[3176] ,
    \all_features[3177] , \all_features[3178] , \all_features[3179] ,
    \all_features[3180] , \all_features[3181] , \all_features[3182] ,
    \all_features[3183] , \all_features[3184] , \all_features[3185] ,
    \all_features[3186] , \all_features[3187] , \all_features[3188] ,
    \all_features[3189] , \all_features[3190] , \all_features[3191] ,
    \all_features[3192] , \all_features[3193] , \all_features[3194] ,
    \all_features[3195] , \all_features[3196] , \all_features[3197] ,
    \all_features[3198] , \all_features[3199] , \all_features[3200] ,
    \all_features[3201] , \all_features[3202] , \all_features[3203] ,
    \all_features[3204] , \all_features[3205] , \all_features[3206] ,
    \all_features[3207] , \all_features[3208] , \all_features[3209] ,
    \all_features[3210] , \all_features[3211] , \all_features[3212] ,
    \all_features[3213] , \all_features[3214] , \all_features[3215] ,
    \all_features[3216] , \all_features[3217] , \all_features[3218] ,
    \all_features[3219] , \all_features[3220] , \all_features[3221] ,
    \all_features[3222] , \all_features[3223] , \all_features[3224] ,
    \all_features[3225] , \all_features[3226] , \all_features[3227] ,
    \all_features[3228] , \all_features[3229] , \all_features[3230] ,
    \all_features[3231] , \all_features[3232] , \all_features[3233] ,
    \all_features[3234] , \all_features[3235] , \all_features[3236] ,
    \all_features[3237] , \all_features[3238] , \all_features[3239] ,
    \all_features[3240] , \all_features[3241] , \all_features[3242] ,
    \all_features[3243] , \all_features[3244] , \all_features[3245] ,
    \all_features[3246] , \all_features[3247] , \all_features[3248] ,
    \all_features[3249] , \all_features[3250] , \all_features[3251] ,
    \all_features[3252] , \all_features[3253] , \all_features[3254] ,
    \all_features[3255] , \all_features[3256] , \all_features[3257] ,
    \all_features[3258] , \all_features[3259] , \all_features[3260] ,
    \all_features[3261] , \all_features[3262] , \all_features[3263] ,
    \all_features[3264] , \all_features[3265] , \all_features[3266] ,
    \all_features[3267] , \all_features[3268] , \all_features[3269] ,
    \all_features[3270] , \all_features[3271] , \all_features[3272] ,
    \all_features[3273] , \all_features[3274] , \all_features[3275] ,
    \all_features[3276] , \all_features[3277] , \all_features[3278] ,
    \all_features[3279] , \all_features[3280] , \all_features[3281] ,
    \all_features[3282] , \all_features[3283] , \all_features[3284] ,
    \all_features[3285] , \all_features[3286] , \all_features[3287] ,
    \all_features[3288] , \all_features[3289] , \all_features[3290] ,
    \all_features[3291] , \all_features[3292] , \all_features[3293] ,
    \all_features[3294] , \all_features[3295] , \all_features[3296] ,
    \all_features[3297] , \all_features[3298] , \all_features[3299] ,
    \all_features[3300] , \all_features[3301] , \all_features[3302] ,
    \all_features[3303] , \all_features[3304] , \all_features[3305] ,
    \all_features[3306] , \all_features[3307] , \all_features[3308] ,
    \all_features[3309] , \all_features[3310] , \all_features[3311] ,
    \all_features[3312] , \all_features[3313] , \all_features[3314] ,
    \all_features[3315] , \all_features[3316] , \all_features[3317] ,
    \all_features[3318] , \all_features[3319] , \all_features[3320] ,
    \all_features[3321] , \all_features[3322] , \all_features[3323] ,
    \all_features[3324] , \all_features[3325] , \all_features[3326] ,
    \all_features[3327] , \all_features[3328] , \all_features[3329] ,
    \all_features[3330] , \all_features[3331] , \all_features[3332] ,
    \all_features[3333] , \all_features[3334] , \all_features[3335] ,
    \all_features[3336] , \all_features[3337] , \all_features[3338] ,
    \all_features[3339] , \all_features[3340] , \all_features[3341] ,
    \all_features[3342] , \all_features[3343] , \all_features[3344] ,
    \all_features[3345] , \all_features[3346] , \all_features[3347] ,
    \all_features[3348] , \all_features[3349] , \all_features[3350] ,
    \all_features[3351] , \all_features[3352] , \all_features[3353] ,
    \all_features[3354] , \all_features[3355] , \all_features[3356] ,
    \all_features[3357] , \all_features[3358] , \all_features[3359] ,
    \all_features[3360] , \all_features[3361] , \all_features[3362] ,
    \all_features[3363] , \all_features[3364] , \all_features[3365] ,
    \all_features[3366] , \all_features[3367] , \all_features[3368] ,
    \all_features[3369] , \all_features[3370] , \all_features[3371] ,
    \all_features[3372] , \all_features[3373] , \all_features[3374] ,
    \all_features[3375] , \all_features[3376] , \all_features[3377] ,
    \all_features[3378] , \all_features[3379] , \all_features[3380] ,
    \all_features[3381] , \all_features[3382] , \all_features[3383] ,
    \all_features[3384] , \all_features[3385] , \all_features[3386] ,
    \all_features[3387] , \all_features[3388] , \all_features[3389] ,
    \all_features[3390] , \all_features[3391] , \all_features[3392] ,
    \all_features[3393] , \all_features[3394] , \all_features[3395] ,
    \all_features[3396] , \all_features[3397] , \all_features[3398] ,
    \all_features[3399] , \all_features[3400] , \all_features[3401] ,
    \all_features[3402] , \all_features[3403] , \all_features[3404] ,
    \all_features[3405] , \all_features[3406] , \all_features[3407] ,
    \all_features[3408] , \all_features[3409] , \all_features[3410] ,
    \all_features[3411] , \all_features[3412] , \all_features[3413] ,
    \all_features[3414] , \all_features[3415] , \all_features[3416] ,
    \all_features[3417] , \all_features[3418] , \all_features[3419] ,
    \all_features[3420] , \all_features[3421] , \all_features[3422] ,
    \all_features[3423] , \all_features[3424] , \all_features[3425] ,
    \all_features[3426] , \all_features[3427] , \all_features[3428] ,
    \all_features[3429] , \all_features[3430] , \all_features[3431] ,
    \all_features[3432] , \all_features[3433] , \all_features[3434] ,
    \all_features[3435] , \all_features[3436] , \all_features[3437] ,
    \all_features[3438] , \all_features[3439] , \all_features[3440] ,
    \all_features[3441] , \all_features[3442] , \all_features[3443] ,
    \all_features[3444] , \all_features[3445] , \all_features[3446] ,
    \all_features[3447] , \all_features[3448] , \all_features[3449] ,
    \all_features[3450] , \all_features[3451] , \all_features[3452] ,
    \all_features[3453] , \all_features[3454] , \all_features[3455] ,
    \all_features[3456] , \all_features[3457] , \all_features[3458] ,
    \all_features[3459] , \all_features[3460] , \all_features[3461] ,
    \all_features[3462] , \all_features[3463] , \all_features[3464] ,
    \all_features[3465] , \all_features[3466] , \all_features[3467] ,
    \all_features[3468] , \all_features[3469] , \all_features[3470] ,
    \all_features[3471] , \all_features[3472] , \all_features[3473] ,
    \all_features[3474] , \all_features[3475] , \all_features[3476] ,
    \all_features[3477] , \all_features[3478] , \all_features[3479] ,
    \all_features[3480] , \all_features[3481] , \all_features[3482] ,
    \all_features[3483] , \all_features[3484] , \all_features[3485] ,
    \all_features[3486] , \all_features[3487] , \all_features[3488] ,
    \all_features[3489] , \all_features[3490] , \all_features[3491] ,
    \all_features[3492] , \all_features[3493] , \all_features[3494] ,
    \all_features[3495] , \all_features[3496] , \all_features[3497] ,
    \all_features[3498] , \all_features[3499] , \all_features[3500] ,
    \all_features[3501] , \all_features[3502] , \all_features[3503] ,
    \all_features[3504] , \all_features[3505] , \all_features[3506] ,
    \all_features[3507] , \all_features[3508] , \all_features[3509] ,
    \all_features[3510] , \all_features[3511] , \all_features[3512] ,
    \all_features[3513] , \all_features[3514] , \all_features[3515] ,
    \all_features[3516] , \all_features[3517] , \all_features[3518] ,
    \all_features[3519] , \all_features[3520] , \all_features[3521] ,
    \all_features[3522] , \all_features[3523] , \all_features[3524] ,
    \all_features[3525] , \all_features[3526] , \all_features[3527] ,
    \all_features[3528] , \all_features[3529] , \all_features[3530] ,
    \all_features[3531] , \all_features[3532] , \all_features[3533] ,
    \all_features[3534] , \all_features[3535] , \all_features[3536] ,
    \all_features[3537] , \all_features[3538] , \all_features[3539] ,
    \all_features[3540] , \all_features[3541] , \all_features[3542] ,
    \all_features[3543] , \all_features[3544] , \all_features[3545] ,
    \all_features[3546] , \all_features[3547] , \all_features[3548] ,
    \all_features[3549] , \all_features[3550] , \all_features[3551] ,
    \all_features[3552] , \all_features[3553] , \all_features[3554] ,
    \all_features[3555] , \all_features[3556] , \all_features[3557] ,
    \all_features[3558] , \all_features[3559] , \all_features[3560] ,
    \all_features[3561] , \all_features[3562] , \all_features[3563] ,
    \all_features[3564] , \all_features[3565] , \all_features[3566] ,
    \all_features[3567] , \all_features[3568] , \all_features[3569] ,
    \all_features[3570] , \all_features[3571] , \all_features[3572] ,
    \all_features[3573] , \all_features[3574] , \all_features[3575] ,
    \all_features[3576] , \all_features[3577] , \all_features[3578] ,
    \all_features[3579] , \all_features[3580] , \all_features[3581] ,
    \all_features[3582] , \all_features[3583] , \all_features[3584] ,
    \all_features[3585] , \all_features[3586] , \all_features[3587] ,
    \all_features[3588] , \all_features[3589] , \all_features[3590] ,
    \all_features[3591] , \all_features[3592] , \all_features[3593] ,
    \all_features[3594] , \all_features[3595] , \all_features[3596] ,
    \all_features[3597] , \all_features[3598] , \all_features[3599] ,
    \all_features[3600] , \all_features[3601] , \all_features[3602] ,
    \all_features[3603] , \all_features[3604] , \all_features[3605] ,
    \all_features[3606] , \all_features[3607] , \all_features[3608] ,
    \all_features[3609] , \all_features[3610] , \all_features[3611] ,
    \all_features[3612] , \all_features[3613] , \all_features[3614] ,
    \all_features[3615] , \all_features[3616] , \all_features[3617] ,
    \all_features[3618] , \all_features[3619] , \all_features[3620] ,
    \all_features[3621] , \all_features[3622] , \all_features[3623] ,
    \all_features[3624] , \all_features[3625] , \all_features[3626] ,
    \all_features[3627] , \all_features[3628] , \all_features[3629] ,
    \all_features[3630] , \all_features[3631] , \all_features[3632] ,
    \all_features[3633] , \all_features[3634] , \all_features[3635] ,
    \all_features[3636] , \all_features[3637] , \all_features[3638] ,
    \all_features[3639] , \all_features[3640] , \all_features[3641] ,
    \all_features[3642] , \all_features[3643] , \all_features[3644] ,
    \all_features[3645] , \all_features[3646] , \all_features[3647] ,
    \all_features[3648] , \all_features[3649] , \all_features[3650] ,
    \all_features[3651] , \all_features[3652] , \all_features[3653] ,
    \all_features[3654] , \all_features[3655] , \all_features[3656] ,
    \all_features[3657] , \all_features[3658] , \all_features[3659] ,
    \all_features[3660] , \all_features[3661] , \all_features[3662] ,
    \all_features[3663] , \all_features[3664] , \all_features[3665] ,
    \all_features[3666] , \all_features[3667] , \all_features[3668] ,
    \all_features[3669] , \all_features[3670] , \all_features[3671] ,
    \all_features[3672] , \all_features[3673] , \all_features[3674] ,
    \all_features[3675] , \all_features[3676] , \all_features[3677] ,
    \all_features[3678] , \all_features[3679] , \all_features[3680] ,
    \all_features[3681] , \all_features[3682] , \all_features[3683] ,
    \all_features[3684] , \all_features[3685] , \all_features[3686] ,
    \all_features[3687] , \all_features[3688] , \all_features[3689] ,
    \all_features[3690] , \all_features[3691] , \all_features[3692] ,
    \all_features[3693] , \all_features[3694] , \all_features[3695] ,
    \all_features[3696] , \all_features[3697] , \all_features[3698] ,
    \all_features[3699] , \all_features[3700] , \all_features[3701] ,
    \all_features[3702] , \all_features[3703] , \all_features[3704] ,
    \all_features[3705] , \all_features[3706] , \all_features[3707] ,
    \all_features[3708] , \all_features[3709] , \all_features[3710] ,
    \all_features[3711] , \all_features[3712] , \all_features[3713] ,
    \all_features[3714] , \all_features[3715] , \all_features[3716] ,
    \all_features[3717] , \all_features[3718] , \all_features[3719] ,
    \all_features[3720] , \all_features[3721] , \all_features[3722] ,
    \all_features[3723] , \all_features[3724] , \all_features[3725] ,
    \all_features[3726] , \all_features[3727] , \all_features[3728] ,
    \all_features[3729] , \all_features[3730] , \all_features[3731] ,
    \all_features[3732] , \all_features[3733] , \all_features[3734] ,
    \all_features[3735] , \all_features[3736] , \all_features[3737] ,
    \all_features[3738] , \all_features[3739] , \all_features[3740] ,
    \all_features[3741] , \all_features[3742] , \all_features[3743] ,
    \all_features[3744] , \all_features[3745] , \all_features[3746] ,
    \all_features[3747] , \all_features[3748] , \all_features[3749] ,
    \all_features[3750] , \all_features[3751] , \all_features[3752] ,
    \all_features[3753] , \all_features[3754] , \all_features[3755] ,
    \all_features[3756] , \all_features[3757] , \all_features[3758] ,
    \all_features[3759] , \all_features[3760] , \all_features[3761] ,
    \all_features[3762] , \all_features[3763] , \all_features[3764] ,
    \all_features[3765] , \all_features[3766] , \all_features[3767] ,
    \all_features[3768] , \all_features[3769] , \all_features[3770] ,
    \all_features[3771] , \all_features[3772] , \all_features[3773] ,
    \all_features[3774] , \all_features[3775] , \all_features[3776] ,
    \all_features[3777] , \all_features[3778] , \all_features[3779] ,
    \all_features[3780] , \all_features[3781] , \all_features[3782] ,
    \all_features[3783] , \all_features[3784] , \all_features[3785] ,
    \all_features[3786] , \all_features[3787] , \all_features[3788] ,
    \all_features[3789] , \all_features[3790] , \all_features[3791] ,
    \all_features[3792] , \all_features[3793] , \all_features[3794] ,
    \all_features[3795] , \all_features[3796] , \all_features[3797] ,
    \all_features[3798] , \all_features[3799] , \all_features[3800] ,
    \all_features[3801] , \all_features[3802] , \all_features[3803] ,
    \all_features[3804] , \all_features[3805] , \all_features[3806] ,
    \all_features[3807] , \all_features[3808] , \all_features[3809] ,
    \all_features[3810] , \all_features[3811] , \all_features[3812] ,
    \all_features[3813] , \all_features[3814] , \all_features[3815] ,
    \all_features[3816] , \all_features[3817] , \all_features[3818] ,
    \all_features[3819] , \all_features[3820] , \all_features[3821] ,
    \all_features[3822] , \all_features[3823] , \all_features[3824] ,
    \all_features[3825] , \all_features[3826] , \all_features[3827] ,
    \all_features[3828] , \all_features[3829] , \all_features[3830] ,
    \all_features[3831] , \all_features[3832] , \all_features[3833] ,
    \all_features[3834] , \all_features[3835] , \all_features[3836] ,
    \all_features[3837] , \all_features[3838] , \all_features[3839] ,
    \all_features[3840] , \all_features[3841] , \all_features[3842] ,
    \all_features[3843] , \all_features[3844] , \all_features[3845] ,
    \all_features[3846] , \all_features[3847] , \all_features[3848] ,
    \all_features[3849] , \all_features[3850] , \all_features[3851] ,
    \all_features[3852] , \all_features[3853] , \all_features[3854] ,
    \all_features[3855] , \all_features[3856] , \all_features[3857] ,
    \all_features[3858] , \all_features[3859] , \all_features[3860] ,
    \all_features[3861] , \all_features[3862] , \all_features[3863] ,
    \all_features[3864] , \all_features[3865] , \all_features[3866] ,
    \all_features[3867] , \all_features[3868] , \all_features[3869] ,
    \all_features[3870] , \all_features[3871] , \all_features[3872] ,
    \all_features[3873] , \all_features[3874] , \all_features[3875] ,
    \all_features[3876] , \all_features[3877] , \all_features[3878] ,
    \all_features[3879] , \all_features[3880] , \all_features[3881] ,
    \all_features[3882] , \all_features[3883] , \all_features[3884] ,
    \all_features[3885] , \all_features[3886] , \all_features[3887] ,
    \all_features[3888] , \all_features[3889] , \all_features[3890] ,
    \all_features[3891] , \all_features[3892] , \all_features[3893] ,
    \all_features[3894] , \all_features[3895] , \all_features[3896] ,
    \all_features[3897] , \all_features[3898] , \all_features[3899] ,
    \all_features[3900] , \all_features[3901] , \all_features[3902] ,
    \all_features[3903] , \all_features[3904] , \all_features[3905] ,
    \all_features[3906] , \all_features[3907] , \all_features[3908] ,
    \all_features[3909] , \all_features[3910] , \all_features[3911] ,
    \all_features[3912] , \all_features[3913] , \all_features[3914] ,
    \all_features[3915] , \all_features[3916] , \all_features[3917] ,
    \all_features[3918] , \all_features[3919] , \all_features[3920] ,
    \all_features[3921] , \all_features[3922] , \all_features[3923] ,
    \all_features[3924] , \all_features[3925] , \all_features[3926] ,
    \all_features[3927] , \all_features[3928] , \all_features[3929] ,
    \all_features[3930] , \all_features[3931] , \all_features[3932] ,
    \all_features[3933] , \all_features[3934] , \all_features[3935] ,
    \all_features[3936] , \all_features[3937] , \all_features[3938] ,
    \all_features[3939] , \all_features[3940] , \all_features[3941] ,
    \all_features[3942] , \all_features[3943] , \all_features[3944] ,
    \all_features[3945] , \all_features[3946] , \all_features[3947] ,
    \all_features[3948] , \all_features[3949] , \all_features[3950] ,
    \all_features[3951] , \all_features[3952] , \all_features[3953] ,
    \all_features[3954] , \all_features[3955] , \all_features[3956] ,
    \all_features[3957] , \all_features[3958] , \all_features[3959] ,
    \all_features[3960] , \all_features[3961] , \all_features[3962] ,
    \all_features[3963] , \all_features[3964] , \all_features[3965] ,
    \all_features[3966] , \all_features[3967] , \all_features[3968] ,
    \all_features[3969] , \all_features[3970] , \all_features[3971] ,
    \all_features[3972] , \all_features[3973] , \all_features[3974] ,
    \all_features[3975] , \all_features[3976] , \all_features[3977] ,
    \all_features[3978] , \all_features[3979] , \all_features[3980] ,
    \all_features[3981] , \all_features[3982] , \all_features[3983] ,
    \all_features[3984] , \all_features[3985] , \all_features[3986] ,
    \all_features[3987] , \all_features[3988] , \all_features[3989] ,
    \all_features[3990] , \all_features[3991] , \all_features[3992] ,
    \all_features[3993] , \all_features[3994] , \all_features[3995] ,
    \all_features[3996] , \all_features[3997] , \all_features[3998] ,
    \all_features[3999] , \all_features[4000] , \all_features[4001] ,
    \all_features[4002] , \all_features[4003] , \all_features[4004] ,
    \all_features[4005] , \all_features[4006] , \all_features[4007] ,
    \all_features[4008] , \all_features[4009] , \all_features[4010] ,
    \all_features[4011] , \all_features[4012] , \all_features[4013] ,
    \all_features[4014] , \all_features[4015] , \all_features[4016] ,
    \all_features[4017] , \all_features[4018] , \all_features[4019] ,
    \all_features[4020] , \all_features[4021] , \all_features[4022] ,
    \all_features[4023] , \all_features[4024] , \all_features[4025] ,
    \all_features[4026] , \all_features[4027] , \all_features[4028] ,
    \all_features[4029] , \all_features[4030] , \all_features[4031] ,
    \all_features[4032] , \all_features[4033] , \all_features[4034] ,
    \all_features[4035] , \all_features[4036] , \all_features[4037] ,
    \all_features[4038] , \all_features[4039] , \all_features[4040] ,
    \all_features[4041] , \all_features[4042] , \all_features[4043] ,
    \all_features[4044] , \all_features[4045] , \all_features[4046] ,
    \all_features[4047] , \all_features[4048] , \all_features[4049] ,
    \all_features[4050] , \all_features[4051] , \all_features[4052] ,
    \all_features[4053] , \all_features[4054] , \all_features[4055] ,
    \all_features[4056] , \all_features[4057] , \all_features[4058] ,
    \all_features[4059] , \all_features[4060] , \all_features[4061] ,
    \all_features[4062] , \all_features[4063] , \all_features[4064] ,
    \all_features[4065] , \all_features[4066] , \all_features[4067] ,
    \all_features[4068] , \all_features[4069] , \all_features[4070] ,
    \all_features[4071] , \all_features[4072] , \all_features[4073] ,
    \all_features[4074] , \all_features[4075] , \all_features[4076] ,
    \all_features[4077] , \all_features[4078] , \all_features[4079] ,
    \all_features[4080] , \all_features[4081] , \all_features[4082] ,
    \all_features[4083] , \all_features[4084] , \all_features[4085] ,
    \all_features[4086] , \all_features[4087] , \all_features[4088] ,
    \all_features[4089] , \all_features[4090] , \all_features[4091] ,
    \all_features[4092] , \all_features[4093] , \all_features[4094] ,
    \all_features[4095] , \all_features[4096] , \all_features[4097] ,
    \all_features[4098] , \all_features[4099] , \all_features[4100] ,
    \all_features[4101] , \all_features[4102] , \all_features[4103] ,
    \all_features[4104] , \all_features[4105] , \all_features[4106] ,
    \all_features[4107] , \all_features[4108] , \all_features[4109] ,
    \all_features[4110] , \all_features[4111] , \all_features[4112] ,
    \all_features[4113] , \all_features[4114] , \all_features[4115] ,
    \all_features[4116] , \all_features[4117] , \all_features[4118] ,
    \all_features[4119] , \all_features[4120] , \all_features[4121] ,
    \all_features[4122] , \all_features[4123] , \all_features[4124] ,
    \all_features[4125] , \all_features[4126] , \all_features[4127] ,
    \all_features[4128] , \all_features[4129] , \all_features[4130] ,
    \all_features[4131] , \all_features[4132] , \all_features[4133] ,
    \all_features[4134] , \all_features[4135] , \all_features[4136] ,
    \all_features[4137] , \all_features[4138] , \all_features[4139] ,
    \all_features[4140] , \all_features[4141] , \all_features[4142] ,
    \all_features[4143] , \all_features[4144] , \all_features[4145] ,
    \all_features[4146] , \all_features[4147] , \all_features[4148] ,
    \all_features[4149] , \all_features[4150] , \all_features[4151] ,
    \all_features[4152] , \all_features[4153] , \all_features[4154] ,
    \all_features[4155] , \all_features[4156] , \all_features[4157] ,
    \all_features[4158] , \all_features[4159] , \all_features[4160] ,
    \all_features[4161] , \all_features[4162] , \all_features[4163] ,
    \all_features[4164] , \all_features[4165] , \all_features[4166] ,
    \all_features[4167] , \all_features[4168] , \all_features[4169] ,
    \all_features[4170] , \all_features[4171] , \all_features[4172] ,
    \all_features[4173] , \all_features[4174] , \all_features[4175] ,
    \all_features[4176] , \all_features[4177] , \all_features[4178] ,
    \all_features[4179] , \all_features[4180] , \all_features[4181] ,
    \all_features[4182] , \all_features[4183] , \all_features[4184] ,
    \all_features[4185] , \all_features[4186] , \all_features[4187] ,
    \all_features[4188] , \all_features[4189] , \all_features[4190] ,
    \all_features[4191] , \all_features[4192] , \all_features[4193] ,
    \all_features[4194] , \all_features[4195] , \all_features[4196] ,
    \all_features[4197] , \all_features[4198] , \all_features[4199] ,
    \all_features[4200] , \all_features[4201] , \all_features[4202] ,
    \all_features[4203] , \all_features[4204] , \all_features[4205] ,
    \all_features[4206] , \all_features[4207] , \all_features[4208] ,
    \all_features[4209] , \all_features[4210] , \all_features[4211] ,
    \all_features[4212] , \all_features[4213] , \all_features[4214] ,
    \all_features[4215] , \all_features[4216] , \all_features[4217] ,
    \all_features[4218] , \all_features[4219] , \all_features[4220] ,
    \all_features[4221] , \all_features[4222] , \all_features[4223] ,
    \all_features[4224] , \all_features[4225] , \all_features[4226] ,
    \all_features[4227] , \all_features[4228] , \all_features[4229] ,
    \all_features[4230] , \all_features[4231] , \all_features[4232] ,
    \all_features[4233] , \all_features[4234] , \all_features[4235] ,
    \all_features[4236] , \all_features[4237] , \all_features[4238] ,
    \all_features[4239] , \all_features[4240] , \all_features[4241] ,
    \all_features[4242] , \all_features[4243] , \all_features[4244] ,
    \all_features[4245] , \all_features[4246] , \all_features[4247] ,
    \all_features[4248] , \all_features[4249] , \all_features[4250] ,
    \all_features[4251] , \all_features[4252] , \all_features[4253] ,
    \all_features[4254] , \all_features[4255] , \all_features[4256] ,
    \all_features[4257] , \all_features[4258] , \all_features[4259] ,
    \all_features[4260] , \all_features[4261] , \all_features[4262] ,
    \all_features[4263] , \all_features[4264] , \all_features[4265] ,
    \all_features[4266] , \all_features[4267] , \all_features[4268] ,
    \all_features[4269] , \all_features[4270] , \all_features[4271] ,
    \all_features[4272] , \all_features[4273] , \all_features[4274] ,
    \all_features[4275] , \all_features[4276] , \all_features[4277] ,
    \all_features[4278] , \all_features[4279] , \all_features[4280] ,
    \all_features[4281] , \all_features[4282] , \all_features[4283] ,
    \all_features[4284] , \all_features[4285] , \all_features[4286] ,
    \all_features[4287] , \all_features[4288] , \all_features[4289] ,
    \all_features[4290] , \all_features[4291] , \all_features[4292] ,
    \all_features[4293] , \all_features[4294] , \all_features[4295] ,
    \all_features[4296] , \all_features[4297] , \all_features[4298] ,
    \all_features[4299] , \all_features[4300] , \all_features[4301] ,
    \all_features[4302] , \all_features[4303] , \all_features[4304] ,
    \all_features[4305] , \all_features[4306] , \all_features[4307] ,
    \all_features[4308] , \all_features[4309] , \all_features[4310] ,
    \all_features[4311] , \all_features[4312] , \all_features[4313] ,
    \all_features[4314] , \all_features[4315] , \all_features[4316] ,
    \all_features[4317] , \all_features[4318] , \all_features[4319] ,
    \all_features[4320] , \all_features[4321] , \all_features[4322] ,
    \all_features[4323] , \all_features[4324] , \all_features[4325] ,
    \all_features[4326] , \all_features[4327] , \all_features[4328] ,
    \all_features[4329] , \all_features[4330] , \all_features[4331] ,
    \all_features[4332] , \all_features[4333] , \all_features[4334] ,
    \all_features[4335] , \all_features[4336] , \all_features[4337] ,
    \all_features[4338] , \all_features[4339] , \all_features[4340] ,
    \all_features[4341] , \all_features[4342] , \all_features[4343] ,
    \all_features[4344] , \all_features[4345] , \all_features[4346] ,
    \all_features[4347] , \all_features[4348] , \all_features[4349] ,
    \all_features[4350] , \all_features[4351] , \all_features[4352] ,
    \all_features[4353] , \all_features[4354] , \all_features[4355] ,
    \all_features[4356] , \all_features[4357] , \all_features[4358] ,
    \all_features[4359] , \all_features[4360] , \all_features[4361] ,
    \all_features[4362] , \all_features[4363] , \all_features[4364] ,
    \all_features[4365] , \all_features[4366] , \all_features[4367] ,
    \all_features[4368] , \all_features[4369] , \all_features[4370] ,
    \all_features[4371] , \all_features[4372] , \all_features[4373] ,
    \all_features[4374] , \all_features[4375] , \all_features[4376] ,
    \all_features[4377] , \all_features[4378] , \all_features[4379] ,
    \all_features[4380] , \all_features[4381] , \all_features[4382] ,
    \all_features[4383] , \all_features[4384] , \all_features[4385] ,
    \all_features[4386] , \all_features[4387] , \all_features[4388] ,
    \all_features[4389] , \all_features[4390] , \all_features[4391] ,
    \all_features[4392] , \all_features[4393] , \all_features[4394] ,
    \all_features[4395] , \all_features[4396] , \all_features[4397] ,
    \all_features[4398] , \all_features[4399] , \all_features[4400] ,
    \all_features[4401] , \all_features[4402] , \all_features[4403] ,
    \all_features[4404] , \all_features[4405] , \all_features[4406] ,
    \all_features[4407] , \all_features[4408] , \all_features[4409] ,
    \all_features[4410] , \all_features[4411] , \all_features[4412] ,
    \all_features[4413] , \all_features[4414] , \all_features[4415] ,
    \all_features[4416] , \all_features[4417] , \all_features[4418] ,
    \all_features[4419] , \all_features[4420] , \all_features[4421] ,
    \all_features[4422] , \all_features[4423] , \all_features[4424] ,
    \all_features[4425] , \all_features[4426] , \all_features[4427] ,
    \all_features[4428] , \all_features[4429] , \all_features[4430] ,
    \all_features[4431] , \all_features[4432] , \all_features[4433] ,
    \all_features[4434] , \all_features[4435] , \all_features[4436] ,
    \all_features[4437] , \all_features[4438] , \all_features[4439] ,
    \all_features[4440] , \all_features[4441] , \all_features[4442] ,
    \all_features[4443] , \all_features[4444] , \all_features[4445] ,
    \all_features[4446] , \all_features[4447] , \all_features[4448] ,
    \all_features[4449] , \all_features[4450] , \all_features[4451] ,
    \all_features[4452] , \all_features[4453] , \all_features[4454] ,
    \all_features[4455] , \all_features[4456] , \all_features[4457] ,
    \all_features[4458] , \all_features[4459] , \all_features[4460] ,
    \all_features[4461] , \all_features[4462] , \all_features[4463] ,
    \all_features[4464] , \all_features[4465] , \all_features[4466] ,
    \all_features[4467] , \all_features[4468] , \all_features[4469] ,
    \all_features[4470] , \all_features[4471] , \all_features[4472] ,
    \all_features[4473] , \all_features[4474] , \all_features[4475] ,
    \all_features[4476] , \all_features[4477] , \all_features[4478] ,
    \all_features[4479] , \all_features[4480] , \all_features[4481] ,
    \all_features[4482] , \all_features[4483] , \all_features[4484] ,
    \all_features[4485] , \all_features[4486] , \all_features[4487] ,
    \all_features[4488] , \all_features[4489] , \all_features[4490] ,
    \all_features[4491] , \all_features[4492] , \all_features[4493] ,
    \all_features[4494] , \all_features[4495] , \all_features[4496] ,
    \all_features[4497] , \all_features[4498] , \all_features[4499] ,
    \all_features[4500] , \all_features[4501] , \all_features[4502] ,
    \all_features[4503] , \all_features[4504] , \all_features[4505] ,
    \all_features[4506] , \all_features[4507] , \all_features[4508] ,
    \all_features[4509] , \all_features[4510] , \all_features[4511] ,
    \all_features[4512] , \all_features[4513] , \all_features[4514] ,
    \all_features[4515] , \all_features[4516] , \all_features[4517] ,
    \all_features[4518] , \all_features[4519] , \all_features[4520] ,
    \all_features[4521] , \all_features[4522] , \all_features[4523] ,
    \all_features[4524] , \all_features[4525] , \all_features[4526] ,
    \all_features[4527] , \all_features[4528] , \all_features[4529] ,
    \all_features[4530] , \all_features[4531] , \all_features[4532] ,
    \all_features[4533] , \all_features[4534] , \all_features[4535] ,
    \all_features[4536] , \all_features[4537] , \all_features[4538] ,
    \all_features[4539] , \all_features[4540] , \all_features[4541] ,
    \all_features[4542] , \all_features[4543] , \all_features[4544] ,
    \all_features[4545] , \all_features[4546] , \all_features[4547] ,
    \all_features[4548] , \all_features[4549] , \all_features[4550] ,
    \all_features[4551] , \all_features[4552] , \all_features[4553] ,
    \all_features[4554] , \all_features[4555] , \all_features[4556] ,
    \all_features[4557] , \all_features[4558] , \all_features[4559] ,
    \all_features[4560] , \all_features[4561] , \all_features[4562] ,
    \all_features[4563] , \all_features[4564] , \all_features[4565] ,
    \all_features[4566] , \all_features[4567] , \all_features[4568] ,
    \all_features[4569] , \all_features[4570] , \all_features[4571] ,
    \all_features[4572] , \all_features[4573] , \all_features[4574] ,
    \all_features[4575] , \all_features[4576] , \all_features[4577] ,
    \all_features[4578] , \all_features[4579] , \all_features[4580] ,
    \all_features[4581] , \all_features[4582] , \all_features[4583] ,
    \all_features[4584] , \all_features[4585] , \all_features[4586] ,
    \all_features[4587] , \all_features[4588] , \all_features[4589] ,
    \all_features[4590] , \all_features[4591] , \all_features[4592] ,
    \all_features[4593] , \all_features[4594] , \all_features[4595] ,
    \all_features[4596] , \all_features[4597] , \all_features[4598] ,
    \all_features[4599] , \all_features[4600] , \all_features[4601] ,
    \all_features[4602] , \all_features[4603] , \all_features[4604] ,
    \all_features[4605] , \all_features[4606] , \all_features[4607] ,
    \all_features[4608] , \all_features[4609] , \all_features[4610] ,
    \all_features[4611] , \all_features[4612] , \all_features[4613] ,
    \all_features[4614] , \all_features[4615] , \all_features[4616] ,
    \all_features[4617] , \all_features[4618] , \all_features[4619] ,
    \all_features[4620] , \all_features[4621] , \all_features[4622] ,
    \all_features[4623] , \all_features[4624] , \all_features[4625] ,
    \all_features[4626] , \all_features[4627] , \all_features[4628] ,
    \all_features[4629] , \all_features[4630] , \all_features[4631] ,
    \all_features[4632] , \all_features[4633] , \all_features[4634] ,
    \all_features[4635] , \all_features[4636] , \all_features[4637] ,
    \all_features[4638] , \all_features[4639] , \all_features[4640] ,
    \all_features[4641] , \all_features[4642] , \all_features[4643] ,
    \all_features[4644] , \all_features[4645] , \all_features[4646] ,
    \all_features[4647] , \all_features[4648] , \all_features[4649] ,
    \all_features[4650] , \all_features[4651] , \all_features[4652] ,
    \all_features[4653] , \all_features[4654] , \all_features[4655] ,
    \all_features[4656] , \all_features[4657] , \all_features[4658] ,
    \all_features[4659] , \all_features[4660] , \all_features[4661] ,
    \all_features[4662] , \all_features[4663] , \all_features[4664] ,
    \all_features[4665] , \all_features[4666] , \all_features[4667] ,
    \all_features[4668] , \all_features[4669] , \all_features[4670] ,
    \all_features[4671] , \all_features[4672] , \all_features[4673] ,
    \all_features[4674] , \all_features[4675] , \all_features[4676] ,
    \all_features[4677] , \all_features[4678] , \all_features[4679] ,
    \all_features[4680] , \all_features[4681] , \all_features[4682] ,
    \all_features[4683] , \all_features[4684] , \all_features[4685] ,
    \all_features[4686] , \all_features[4687] , \all_features[4688] ,
    \all_features[4689] , \all_features[4690] , \all_features[4691] ,
    \all_features[4692] , \all_features[4693] , \all_features[4694] ,
    \all_features[4695] , \all_features[4696] , \all_features[4697] ,
    \all_features[4698] , \all_features[4699] , \all_features[4700] ,
    \all_features[4701] , \all_features[4702] , \all_features[4703] ,
    \all_features[4704] , \all_features[4705] , \all_features[4706] ,
    \all_features[4707] , \all_features[4708] , \all_features[4709] ,
    \all_features[4710] , \all_features[4711] , \all_features[4712] ,
    \all_features[4713] , \all_features[4714] , \all_features[4715] ,
    \all_features[4716] , \all_features[4717] , \all_features[4718] ,
    \all_features[4719] , \all_features[4720] , \all_features[4721] ,
    \all_features[4722] , \all_features[4723] , \all_features[4724] ,
    \all_features[4725] , \all_features[4726] , \all_features[4727] ,
    \all_features[4728] , \all_features[4729] , \all_features[4730] ,
    \all_features[4731] , \all_features[4732] , \all_features[4733] ,
    \all_features[4734] , \all_features[4735] , \all_features[4736] ,
    \all_features[4737] , \all_features[4738] , \all_features[4739] ,
    \all_features[4740] , \all_features[4741] , \all_features[4742] ,
    \all_features[4743] , \all_features[4744] , \all_features[4745] ,
    \all_features[4746] , \all_features[4747] , \all_features[4748] ,
    \all_features[4749] , \all_features[4750] , \all_features[4751] ,
    \all_features[4752] , \all_features[4753] , \all_features[4754] ,
    \all_features[4755] , \all_features[4756] , \all_features[4757] ,
    \all_features[4758] , \all_features[4759] , \all_features[4760] ,
    \all_features[4761] , \all_features[4762] , \all_features[4763] ,
    \all_features[4764] , \all_features[4765] , \all_features[4766] ,
    \all_features[4767] , \all_features[4768] , \all_features[4769] ,
    \all_features[4770] , \all_features[4771] , \all_features[4772] ,
    \all_features[4773] , \all_features[4774] , \all_features[4775] ,
    \all_features[4776] , \all_features[4777] , \all_features[4778] ,
    \all_features[4779] , \all_features[4780] , \all_features[4781] ,
    \all_features[4782] , \all_features[4783] , \all_features[4784] ,
    \all_features[4785] , \all_features[4786] , \all_features[4787] ,
    \all_features[4788] , \all_features[4789] , \all_features[4790] ,
    \all_features[4791] , \all_features[4792] , \all_features[4793] ,
    \all_features[4794] , \all_features[4795] , \all_features[4796] ,
    \all_features[4797] , \all_features[4798] , \all_features[4799] ,
    \all_features[4800] , \all_features[4801] , \all_features[4802] ,
    \all_features[4803] , \all_features[4804] , \all_features[4805] ,
    \all_features[4806] , \all_features[4807] , \all_features[4808] ,
    \all_features[4809] , \all_features[4810] , \all_features[4811] ,
    \all_features[4812] , \all_features[4813] , \all_features[4814] ,
    \all_features[4815] , \all_features[4816] , \all_features[4817] ,
    \all_features[4818] , \all_features[4819] , \all_features[4820] ,
    \all_features[4821] , \all_features[4822] , \all_features[4823] ,
    \all_features[4824] , \all_features[4825] , \all_features[4826] ,
    \all_features[4827] , \all_features[4828] , \all_features[4829] ,
    \all_features[4830] , \all_features[4831] , \all_features[4832] ,
    \all_features[4833] , \all_features[4834] , \all_features[4835] ,
    \all_features[4836] , \all_features[4837] , \all_features[4838] ,
    \all_features[4839] , \all_features[4840] , \all_features[4841] ,
    \all_features[4842] , \all_features[4843] , \all_features[4844] ,
    \all_features[4845] , \all_features[4846] , \all_features[4847] ,
    \all_features[4848] , \all_features[4849] , \all_features[4850] ,
    \all_features[4851] , \all_features[4852] , \all_features[4853] ,
    \all_features[4854] , \all_features[4855] , \all_features[4856] ,
    \all_features[4857] , \all_features[4858] , \all_features[4859] ,
    \all_features[4860] , \all_features[4861] , \all_features[4862] ,
    \all_features[4863] , \all_features[4864] , \all_features[4865] ,
    \all_features[4866] , \all_features[4867] , \all_features[4868] ,
    \all_features[4869] , \all_features[4870] , \all_features[4871] ,
    \all_features[4872] , \all_features[4873] , \all_features[4874] ,
    \all_features[4875] , \all_features[4876] , \all_features[4877] ,
    \all_features[4878] , \all_features[4879] , \all_features[4880] ,
    \all_features[4881] , \all_features[4882] , \all_features[4883] ,
    \all_features[4884] , \all_features[4885] , \all_features[4886] ,
    \all_features[4887] , \all_features[4888] , \all_features[4889] ,
    \all_features[4890] , \all_features[4891] , \all_features[4892] ,
    \all_features[4893] , \all_features[4894] , \all_features[4895] ,
    \all_features[4896] , \all_features[4897] , \all_features[4898] ,
    \all_features[4899] , \all_features[4900] , \all_features[4901] ,
    \all_features[4902] , \all_features[4903] , \all_features[4904] ,
    \all_features[4905] , \all_features[4906] , \all_features[4907] ,
    \all_features[4908] , \all_features[4909] , \all_features[4910] ,
    \all_features[4911] , \all_features[4912] , \all_features[4913] ,
    \all_features[4914] , \all_features[4915] , \all_features[4916] ,
    \all_features[4917] , \all_features[4918] , \all_features[4919] ,
    \all_features[4920] , \all_features[4921] , \all_features[4922] ,
    \all_features[4923] , \all_features[4924] , \all_features[4925] ,
    \all_features[4926] , \all_features[4927] , \all_features[4928] ,
    \all_features[4929] , \all_features[4930] , \all_features[4931] ,
    \all_features[4932] , \all_features[4933] , \all_features[4934] ,
    \all_features[4935] , \all_features[4936] , \all_features[4937] ,
    \all_features[4938] , \all_features[4939] , \all_features[4940] ,
    \all_features[4941] , \all_features[4942] , \all_features[4943] ,
    \all_features[4944] , \all_features[4945] , \all_features[4946] ,
    \all_features[4947] , \all_features[4948] , \all_features[4949] ,
    \all_features[4950] , \all_features[4951] , \all_features[4952] ,
    \all_features[4953] , \all_features[4954] , \all_features[4955] ,
    \all_features[4956] , \all_features[4957] , \all_features[4958] ,
    \all_features[4959] , \all_features[4960] , \all_features[4961] ,
    \all_features[4962] , \all_features[4963] , \all_features[4964] ,
    \all_features[4965] , \all_features[4966] , \all_features[4967] ,
    \all_features[4968] , \all_features[4969] , \all_features[4970] ,
    \all_features[4971] , \all_features[4972] , \all_features[4973] ,
    \all_features[4974] , \all_features[4975] , \all_features[4976] ,
    \all_features[4977] , \all_features[4978] , \all_features[4979] ,
    \all_features[4980] , \all_features[4981] , \all_features[4982] ,
    \all_features[4983] , \all_features[4984] , \all_features[4985] ,
    \all_features[4986] , \all_features[4987] , \all_features[4988] ,
    \all_features[4989] , \all_features[4990] , \all_features[4991] ,
    \all_features[4992] , \all_features[4993] , \all_features[4994] ,
    \all_features[4995] , \all_features[4996] , \all_features[4997] ,
    \all_features[4998] , \all_features[4999] , \all_features[5000] ,
    \all_features[5001] , \all_features[5002] , \all_features[5003] ,
    \all_features[5004] , \all_features[5005] , \all_features[5006] ,
    \all_features[5007] , \all_features[5008] , \all_features[5009] ,
    \all_features[5010] , \all_features[5011] , \all_features[5012] ,
    \all_features[5013] , \all_features[5014] , \all_features[5015] ,
    \all_features[5016] , \all_features[5017] , \all_features[5018] ,
    \all_features[5019] , \all_features[5020] , \all_features[5021] ,
    \all_features[5022] , \all_features[5023] , \all_features[5024] ,
    \all_features[5025] , \all_features[5026] , \all_features[5027] ,
    \all_features[5028] , \all_features[5029] , \all_features[5030] ,
    \all_features[5031] , \all_features[5032] , \all_features[5033] ,
    \all_features[5034] , \all_features[5035] , \all_features[5036] ,
    \all_features[5037] , \all_features[5038] , \all_features[5039] ,
    \all_features[5040] , \all_features[5041] , \all_features[5042] ,
    \all_features[5043] , \all_features[5044] , \all_features[5045] ,
    \all_features[5046] , \all_features[5047] , \all_features[5048] ,
    \all_features[5049] , \all_features[5050] , \all_features[5051] ,
    \all_features[5052] , \all_features[5053] , \all_features[5054] ,
    \all_features[5055] , \all_features[5056] , \all_features[5057] ,
    \all_features[5058] , \all_features[5059] , \all_features[5060] ,
    \all_features[5061] , \all_features[5062] , \all_features[5063] ,
    \all_features[5064] , \all_features[5065] , \all_features[5066] ,
    \all_features[5067] , \all_features[5068] , \all_features[5069] ,
    \all_features[5070] , \all_features[5071] , \all_features[5072] ,
    \all_features[5073] , \all_features[5074] , \all_features[5075] ,
    \all_features[5076] , \all_features[5077] , \all_features[5078] ,
    \all_features[5079] , \all_features[5080] , \all_features[5081] ,
    \all_features[5082] , \all_features[5083] , \all_features[5084] ,
    \all_features[5085] , \all_features[5086] , \all_features[5087] ,
    \all_features[5088] , \all_features[5089] , \all_features[5090] ,
    \all_features[5091] , \all_features[5092] , \all_features[5093] ,
    \all_features[5094] , \all_features[5095] , \all_features[5096] ,
    \all_features[5097] , \all_features[5098] , \all_features[5099] ,
    \all_features[5100] , \all_features[5101] , \all_features[5102] ,
    \all_features[5103] , \all_features[5104] , \all_features[5105] ,
    \all_features[5106] , \all_features[5107] , \all_features[5108] ,
    \all_features[5109] , \all_features[5110] , \all_features[5111] ,
    \all_features[5112] , \all_features[5113] , \all_features[5114] ,
    \all_features[5115] , \all_features[5116] , \all_features[5117] ,
    \all_features[5118] , \all_features[5119] , \all_features[5120] ,
    \all_features[5121] , \all_features[5122] , \all_features[5123] ,
    \all_features[5124] , \all_features[5125] , \all_features[5126] ,
    \all_features[5127] , \all_features[5128] , \all_features[5129] ,
    \all_features[5130] , \all_features[5131] , \all_features[5132] ,
    \all_features[5133] , \all_features[5134] , \all_features[5135] ,
    \all_features[5136] , \all_features[5137] , \all_features[5138] ,
    \all_features[5139] , \all_features[5140] , \all_features[5141] ,
    \all_features[5142] , \all_features[5143] , \all_features[5144] ,
    \all_features[5145] , \all_features[5146] , \all_features[5147] ,
    \all_features[5148] , \all_features[5149] , \all_features[5150] ,
    \all_features[5151] , \all_features[5152] , \all_features[5153] ,
    \all_features[5154] , \all_features[5155] , \all_features[5156] ,
    \all_features[5157] , \all_features[5158] , \all_features[5159] ,
    \all_features[5160] , \all_features[5161] , \all_features[5162] ,
    \all_features[5163] , \all_features[5164] , \all_features[5165] ,
    \all_features[5166] , \all_features[5167] , \all_features[5168] ,
    \all_features[5169] , \all_features[5170] , \all_features[5171] ,
    \all_features[5172] , \all_features[5173] , \all_features[5174] ,
    \all_features[5175] , \all_features[5176] , \all_features[5177] ,
    \all_features[5178] , \all_features[5179] , \all_features[5180] ,
    \all_features[5181] , \all_features[5182] , \all_features[5183] ,
    \all_features[5184] , \all_features[5185] , \all_features[5186] ,
    \all_features[5187] , \all_features[5188] , \all_features[5189] ,
    \all_features[5190] , \all_features[5191] , \all_features[5192] ,
    \all_features[5193] , \all_features[5194] , \all_features[5195] ,
    \all_features[5196] , \all_features[5197] , \all_features[5198] ,
    \all_features[5199] , \all_features[5200] , \all_features[5201] ,
    \all_features[5202] , \all_features[5203] , \all_features[5204] ,
    \all_features[5205] , \all_features[5206] , \all_features[5207] ,
    \all_features[5208] , \all_features[5209] , \all_features[5210] ,
    \all_features[5211] , \all_features[5212] , \all_features[5213] ,
    \all_features[5214] , \all_features[5215] , \all_features[5216] ,
    \all_features[5217] , \all_features[5218] , \all_features[5219] ,
    \all_features[5220] , \all_features[5221] , \all_features[5222] ,
    \all_features[5223] , \all_features[5224] , \all_features[5225] ,
    \all_features[5226] , \all_features[5227] , \all_features[5228] ,
    \all_features[5229] , \all_features[5230] , \all_features[5231] ,
    \all_features[5232] , \all_features[5233] , \all_features[5234] ,
    \all_features[5235] , \all_features[5236] , \all_features[5237] ,
    \all_features[5238] , \all_features[5239] , \all_features[5240] ,
    \all_features[5241] , \all_features[5242] , \all_features[5243] ,
    \all_features[5244] , \all_features[5245] , \all_features[5246] ,
    \all_features[5247] , \all_features[5248] , \all_features[5249] ,
    \all_features[5250] , \all_features[5251] , \all_features[5252] ,
    \all_features[5253] , \all_features[5254] , \all_features[5255] ,
    \all_features[5256] , \all_features[5257] , \all_features[5258] ,
    \all_features[5259] , \all_features[5260] , \all_features[5261] ,
    \all_features[5262] , \all_features[5263] , \all_features[5264] ,
    \all_features[5265] , \all_features[5266] , \all_features[5267] ,
    \all_features[5268] , \all_features[5269] , \all_features[5270] ,
    \all_features[5271] , \all_features[5272] , \all_features[5273] ,
    \all_features[5274] , \all_features[5275] , \all_features[5276] ,
    \all_features[5277] , \all_features[5278] , \all_features[5279] ,
    \all_features[5280] , \all_features[5281] , \all_features[5282] ,
    \all_features[5283] , \all_features[5284] , \all_features[5285] ,
    \all_features[5286] , \all_features[5287] , \all_features[5288] ,
    \all_features[5289] , \all_features[5290] , \all_features[5291] ,
    \all_features[5292] , \all_features[5293] , \all_features[5294] ,
    \all_features[5295] , \all_features[5296] , \all_features[5297] ,
    \all_features[5298] , \all_features[5299] , \all_features[5300] ,
    \all_features[5301] , \all_features[5302] , \all_features[5303] ,
    \all_features[5304] , \all_features[5305] , \all_features[5306] ,
    \all_features[5307] , \all_features[5308] , \all_features[5309] ,
    \all_features[5310] , \all_features[5311] , \all_features[5312] ,
    \all_features[5313] , \all_features[5314] , \all_features[5315] ,
    \all_features[5316] , \all_features[5317] , \all_features[5318] ,
    \all_features[5319] , \all_features[5320] , \all_features[5321] ,
    \all_features[5322] , \all_features[5323] , \all_features[5324] ,
    \all_features[5325] , \all_features[5326] , \all_features[5327] ,
    \all_features[5328] , \all_features[5329] , \all_features[5330] ,
    \all_features[5331] , \all_features[5332] , \all_features[5333] ,
    \all_features[5334] , \all_features[5335] , \all_features[5336] ,
    \all_features[5337] , \all_features[5338] , \all_features[5339] ,
    \all_features[5340] , \all_features[5341] , \all_features[5342] ,
    \all_features[5343] , \all_features[5344] , \all_features[5345] ,
    \all_features[5346] , \all_features[5347] , \all_features[5348] ,
    \all_features[5349] , \all_features[5350] , \all_features[5351] ,
    \all_features[5352] , \all_features[5353] , \all_features[5354] ,
    \all_features[5355] , \all_features[5356] , \all_features[5357] ,
    \all_features[5358] , \all_features[5359] , \all_features[5360] ,
    \all_features[5361] , \all_features[5362] , \all_features[5363] ,
    \all_features[5364] , \all_features[5365] , \all_features[5366] ,
    \all_features[5367] , \all_features[5368] , \all_features[5369] ,
    \all_features[5370] , \all_features[5371] , \all_features[5372] ,
    \all_features[5373] , \all_features[5374] , \all_features[5375] ,
    \all_features[5376] , \all_features[5377] , \all_features[5378] ,
    \all_features[5379] , \all_features[5380] , \all_features[5381] ,
    \all_features[5382] , \all_features[5383] , \all_features[5384] ,
    \all_features[5385] , \all_features[5386] , \all_features[5387] ,
    \all_features[5388] , \all_features[5389] , \all_features[5390] ,
    \all_features[5391] , \all_features[5392] , \all_features[5393] ,
    \all_features[5394] , \all_features[5395] , \all_features[5396] ,
    \all_features[5397] , \all_features[5398] , \all_features[5399] ,
    \all_features[5400] , \all_features[5401] , \all_features[5402] ,
    \all_features[5403] , \all_features[5404] , \all_features[5405] ,
    \all_features[5406] , \all_features[5407] , \all_features[5408] ,
    \all_features[5409] , \all_features[5410] , \all_features[5411] ,
    \all_features[5412] , \all_features[5413] , \all_features[5414] ,
    \all_features[5415] , \all_features[5416] , \all_features[5417] ,
    \all_features[5418] , \all_features[5419] , \all_features[5420] ,
    \all_features[5421] , \all_features[5422] , \all_features[5423] ,
    \all_features[5424] , \all_features[5425] , \all_features[5426] ,
    \all_features[5427] , \all_features[5428] , \all_features[5429] ,
    \all_features[5430] , \all_features[5431] , \all_features[5432] ,
    \all_features[5433] , \all_features[5434] , \all_features[5435] ,
    \all_features[5436] , \all_features[5437] , \all_features[5438] ,
    \all_features[5439] , \all_features[5440] , \all_features[5441] ,
    \all_features[5442] , \all_features[5443] , \all_features[5444] ,
    \all_features[5445] , \all_features[5446] , \all_features[5447] ,
    \all_features[5448] , \all_features[5449] , \all_features[5450] ,
    \all_features[5451] , \all_features[5452] , \all_features[5453] ,
    \all_features[5454] , \all_features[5455] , \all_features[5456] ,
    \all_features[5457] , \all_features[5458] , \all_features[5459] ,
    \all_features[5460] , \all_features[5461] , \all_features[5462] ,
    \all_features[5463] , \all_features[5464] , \all_features[5465] ,
    \all_features[5466] , \all_features[5467] , \all_features[5468] ,
    \all_features[5469] , \all_features[5470] , \all_features[5471] ,
    \all_features[5472] , \all_features[5473] , \all_features[5474] ,
    \all_features[5475] , \all_features[5476] , \all_features[5477] ,
    \all_features[5478] , \all_features[5479] , \all_features[5480] ,
    \all_features[5481] , \all_features[5482] , \all_features[5483] ,
    \all_features[5484] , \all_features[5485] , \all_features[5486] ,
    \all_features[5487] , \all_features[5488] , \all_features[5489] ,
    \all_features[5490] , \all_features[5491] , \all_features[5492] ,
    \all_features[5493] , \all_features[5494] , \all_features[5495] ,
    \all_features[5496] , \all_features[5497] , \all_features[5498] ,
    \all_features[5499] , \all_features[5500] , \all_features[5501] ,
    \all_features[5502] , \all_features[5503] , \all_features[5504] ,
    \all_features[5505] , \all_features[5506] , \all_features[5507] ,
    \all_features[5508] , \all_features[5509] , \all_features[5510] ,
    \all_features[5511] , \all_features[5512] , \all_features[5513] ,
    \all_features[5514] , \all_features[5515] , \all_features[5516] ,
    \all_features[5517] , \all_features[5518] , \all_features[5519] ,
    \all_features[5520] , \all_features[5521] , \all_features[5522] ,
    \all_features[5523] , \all_features[5524] , \all_features[5525] ,
    \all_features[5526] , \all_features[5527] , \all_features[5528] ,
    \all_features[5529] , \all_features[5530] , \all_features[5531] ,
    \all_features[5532] , \all_features[5533] , \all_features[5534] ,
    \all_features[5535] , \all_features[5536] , \all_features[5537] ,
    \all_features[5538] , \all_features[5539] , \all_features[5540] ,
    \all_features[5541] , \all_features[5542] , \all_features[5543] ,
    \all_features[5544] , \all_features[5545] , \all_features[5546] ,
    \all_features[5547] , \all_features[5548] , \all_features[5549] ,
    \all_features[5550] , \all_features[5551] , \all_features[5552] ,
    \all_features[5553] , \all_features[5554] , \all_features[5555] ,
    \all_features[5556] , \all_features[5557] , \all_features[5558] ,
    \all_features[5559] , \all_features[5560] , \all_features[5561] ,
    \all_features[5562] , \all_features[5563] , \all_features[5564] ,
    \all_features[5565] , \all_features[5566] , \all_features[5567] ,
    \all_features[5568] , \all_features[5569] , \all_features[5570] ,
    \all_features[5571] , \all_features[5572] , \all_features[5573] ,
    \all_features[5574] , \all_features[5575] , \all_features[5576] ,
    \all_features[5577] , \all_features[5578] , \all_features[5579] ,
    \all_features[5580] , \all_features[5581] , \all_features[5582] ,
    \all_features[5583] , \all_features[5584] , \all_features[5585] ,
    \all_features[5586] , \all_features[5587] , \all_features[5588] ,
    \all_features[5589] , \all_features[5590] , \all_features[5591] ,
    \all_features[5592] , \all_features[5593] , \all_features[5594] ,
    \all_features[5595] , \all_features[5596] , \all_features[5597] ,
    \all_features[5598] , \all_features[5599] , \all_features[5600] ,
    \all_features[5601] , \all_features[5602] , \all_features[5603] ,
    \all_features[5604] , \all_features[5605] , \all_features[5606] ,
    \all_features[5607] , \all_features[5608] , \all_features[5609] ,
    \all_features[5610] , \all_features[5611] , \all_features[5612] ,
    \all_features[5613] , \all_features[5614] , \all_features[5615] ,
    \all_features[5616] , \all_features[5617] , \all_features[5618] ,
    \all_features[5619] , \all_features[5620] , \all_features[5621] ,
    \all_features[5622] , \all_features[5623] , \all_features[5624] ,
    \all_features[5625] , \all_features[5626] , \all_features[5627] ,
    \all_features[5628] , \all_features[5629] , \all_features[5630] ,
    \all_features[5631] , \all_features[5632] , \all_features[5633] ,
    \all_features[5634] , \all_features[5635] , \all_features[5636] ,
    \all_features[5637] , \all_features[5638] , \all_features[5639] ,
    \all_features[5640] , \all_features[5641] , \all_features[5642] ,
    \all_features[5643] , \all_features[5644] , \all_features[5645] ,
    \all_features[5646] , \all_features[5647] , \all_features[5648] ,
    \all_features[5649] , \all_features[5650] , \all_features[5651] ,
    \all_features[5652] , \all_features[5653] , \all_features[5654] ,
    \all_features[5655] , \all_features[5656] , \all_features[5657] ,
    \all_features[5658] , \all_features[5659] , \all_features[5660] ,
    \all_features[5661] , \all_features[5662] , \all_features[5663] ,
    \all_features[5664] , \all_features[5665] , \all_features[5666] ,
    \all_features[5667] , \all_features[5668] , \all_features[5669] ,
    \all_features[5670] , \all_features[5671] , \all_features[5672] ,
    \all_features[5673] , \all_features[5674] , \all_features[5675] ,
    \all_features[5676] , \all_features[5677] , \all_features[5678] ,
    \all_features[5679] , \all_features[5680] , \all_features[5681] ,
    \all_features[5682] , \all_features[5683] , \all_features[5684] ,
    \all_features[5685] , \all_features[5686] , \all_features[5687] ,
    \all_features[5688] , \all_features[5689] , \all_features[5690] ,
    \all_features[5691] , \all_features[5692] , \all_features[5693] ,
    \all_features[5694] , \all_features[5695] , \all_features[5696] ,
    \all_features[5697] , \all_features[5698] , \all_features[5699] ,
    \all_features[5700] , \all_features[5701] , \all_features[5702] ,
    \all_features[5703] , \all_features[5704] , \all_features[5705] ,
    \all_features[5706] , \all_features[5707] , \all_features[5708] ,
    \all_features[5709] , \all_features[5710] , \all_features[5711] ,
    \all_features[5712] , \all_features[5713] , \all_features[5714] ,
    \all_features[5715] , \all_features[5716] , \all_features[5717] ,
    \all_features[5718] , \all_features[5719] , \all_features[5720] ,
    \all_features[5721] , \all_features[5722] , \all_features[5723] ,
    \all_features[5724] , \all_features[5725] , \all_features[5726] ,
    \all_features[5727] , \all_features[5728] , \all_features[5729] ,
    \all_features[5730] , \all_features[5731] , \all_features[5732] ,
    \all_features[5733] , \all_features[5734] , \all_features[5735] ,
    \all_features[5736] , \all_features[5737] , \all_features[5738] ,
    \all_features[5739] , \all_features[5740] , \all_features[5741] ,
    \all_features[5742] , \all_features[5743] , \all_features[5744] ,
    \all_features[5745] , \all_features[5746] , \all_features[5747] ,
    \all_features[5748] , \all_features[5749] , \all_features[5750] ,
    \all_features[5751] , \all_features[5752] , \all_features[5753] ,
    \all_features[5754] , \all_features[5755] , \all_features[5756] ,
    \all_features[5757] , \all_features[5758] , \all_features[5759] ,
    \all_features[5760] , \all_features[5761] , \all_features[5762] ,
    \all_features[5763] , \all_features[5764] , \all_features[5765] ,
    \all_features[5766] , \all_features[5767] , \all_features[5768] ,
    \all_features[5769] , \all_features[5770] , \all_features[5771] ,
    \all_features[5772] , \all_features[5773] , \all_features[5774] ,
    \all_features[5775] , \all_features[5776] , \all_features[5777] ,
    \all_features[5778] , \all_features[5779] , \all_features[5780] ,
    \all_features[5781] , \all_features[5782] , \all_features[5783] ,
    \all_features[5784] , \all_features[5785] , \all_features[5786] ,
    \all_features[5787] , \all_features[5788] , \all_features[5789] ,
    \all_features[5790] , \all_features[5791] , \all_features[5792] ,
    \all_features[5793] , \all_features[5794] , \all_features[5795] ,
    \all_features[5796] , \all_features[5797] , \all_features[5798] ,
    \all_features[5799] , \all_features[5800] , \all_features[5801] ,
    \all_features[5802] , \all_features[5803] , \all_features[5804] ,
    \all_features[5805] , \all_features[5806] , \all_features[5807] ,
    \all_features[5808] , \all_features[5809] , \all_features[5810] ,
    \all_features[5811] , \all_features[5812] , \all_features[5813] ,
    \all_features[5814] , \all_features[5815] , \all_features[5816] ,
    \all_features[5817] , \all_features[5818] , \all_features[5819] ,
    \all_features[5820] , \all_features[5821] , \all_features[5822] ,
    \all_features[5823] , \all_features[5824] , \all_features[5825] ,
    \all_features[5826] , \all_features[5827] , \all_features[5828] ,
    \all_features[5829] , \all_features[5830] , \all_features[5831] ,
    \all_features[5832] , \all_features[5833] , \all_features[5834] ,
    \all_features[5835] , \all_features[5836] , \all_features[5837] ,
    \all_features[5838] , \all_features[5839] , \all_features[5840] ,
    \all_features[5841] , \all_features[5842] , \all_features[5843] ,
    \all_features[5844] , \all_features[5845] , \all_features[5846] ,
    \all_features[5847] , \all_features[5848] , \all_features[5849] ,
    \all_features[5850] , \all_features[5851] , \all_features[5852] ,
    \all_features[5853] , \all_features[5854] , \all_features[5855] ,
    \all_features[5856] , \all_features[5857] , \all_features[5858] ,
    \all_features[5859] , \all_features[5860] , \all_features[5861] ,
    \all_features[5862] , \all_features[5863] , \all_features[5864] ,
    \all_features[5865] , \all_features[5866] , \all_features[5867] ,
    \all_features[5868] , \all_features[5869] , \all_features[5870] ,
    \all_features[5871] , \all_features[5872] , \all_features[5873] ,
    \all_features[5874] , \all_features[5875] , \all_features[5876] ,
    \all_features[5877] , \all_features[5878] , \all_features[5879] ,
    \all_features[5880] , \all_features[5881] , \all_features[5882] ,
    \all_features[5883] , \all_features[5884] , \all_features[5885] ,
    \all_features[5886] , \all_features[5887] , \all_features[5888] ,
    \all_features[5889] , \all_features[5890] , \all_features[5891] ,
    \all_features[5892] , \all_features[5893] , \all_features[5894] ,
    \all_features[5895] , \all_features[5896] , \all_features[5897] ,
    \all_features[5898] , \all_features[5899] , \all_features[5900] ,
    \all_features[5901] , \all_features[5902] , \all_features[5903] ,
    \all_features[5904] , \all_features[5905] , \all_features[5906] ,
    \all_features[5907] , \all_features[5908] , \all_features[5909] ,
    \all_features[5910] , \all_features[5911] , \all_features[5912] ,
    \all_features[5913] , \all_features[5914] , \all_features[5915] ,
    \all_features[5916] , \all_features[5917] , \all_features[5918] ,
    \all_features[5919] , \all_features[5920] , \all_features[5921] ,
    \all_features[5922] , \all_features[5923] , \all_features[5924] ,
    \all_features[5925] , \all_features[5926] , \all_features[5927] ,
    \all_features[5928] , \all_features[5929] , \all_features[5930] ,
    \all_features[5931] , \all_features[5932] , \all_features[5933] ,
    \all_features[5934] , \all_features[5935] , \all_features[5936] ,
    \all_features[5937] , \all_features[5938] , \all_features[5939] ,
    \all_features[5940] , \all_features[5941] , \all_features[5942] ,
    \all_features[5943] , \all_features[5944] , \all_features[5945] ,
    \all_features[5946] , \all_features[5947] , \all_features[5948] ,
    \all_features[5949] , \all_features[5950] , \all_features[5951] ,
    \all_features[5952] , \all_features[5953] , \all_features[5954] ,
    \all_features[5955] , \all_features[5956] , \all_features[5957] ,
    \all_features[5958] , \all_features[5959] , \all_features[5960] ,
    \all_features[5961] , \all_features[5962] , \all_features[5963] ,
    \all_features[5964] , \all_features[5965] , \all_features[5966] ,
    \all_features[5967] , \all_features[5968] , \all_features[5969] ,
    \all_features[5970] , \all_features[5971] , \all_features[5972] ,
    \all_features[5973] , \all_features[5974] , \all_features[5975] ,
    \all_features[5976] , \all_features[5977] , \all_features[5978] ,
    \all_features[5979] , \all_features[5980] , \all_features[5981] ,
    \all_features[5982] , \all_features[5983] , \all_features[5984] ,
    \all_features[5985] , \all_features[5986] , \all_features[5987] ,
    \all_features[5988] , \all_features[5989] , \all_features[5990] ,
    \all_features[5991] , \all_features[5992] , \all_features[5993] ,
    \all_features[5994] , \all_features[5995] , \all_features[5996] ,
    \all_features[5997] , \all_features[5998] , \all_features[5999] ,
    \all_features[6000] , \all_features[6001] , \all_features[6002] ,
    \all_features[6003] , \all_features[6004] , \all_features[6005] ,
    \all_features[6006] , \all_features[6007] , \all_features[6008] ,
    \all_features[6009] , \all_features[6010] , \all_features[6011] ,
    \all_features[6012] , \all_features[6013] , \all_features[6014] ,
    \all_features[6015] , \all_features[6016] , \all_features[6017] ,
    \all_features[6018] , \all_features[6019] , \all_features[6020] ,
    \all_features[6021] , \all_features[6022] , \all_features[6023] ,
    \all_features[6024] , \all_features[6025] , \all_features[6026] ,
    \all_features[6027] , \all_features[6028] , \all_features[6029] ,
    \all_features[6030] , \all_features[6031] , \all_features[6032] ,
    \all_features[6033] , \all_features[6034] , \all_features[6035] ,
    \all_features[6036] , \all_features[6037] , \all_features[6038] ,
    \all_features[6039] , \all_features[6040] , \all_features[6041] ,
    \all_features[6042] , \all_features[6043] , \all_features[6044] ,
    \all_features[6045] , \all_features[6046] , \all_features[6047] ,
    \all_features[6048] , \all_features[6049] , \all_features[6050] ,
    \all_features[6051] , \all_features[6052] , \all_features[6053] ,
    \all_features[6054] , \all_features[6055] , \all_features[6056] ,
    \all_features[6057] , \all_features[6058] , \all_features[6059] ,
    \all_features[6060] , \all_features[6061] , \all_features[6062] ,
    \all_features[6063] , \all_features[6064] , \all_features[6065] ,
    \all_features[6066] , \all_features[6067] , \all_features[6068] ,
    \all_features[6069] , \all_features[6070] , \all_features[6071] ,
    \all_features[6072] , \all_features[6073] , \all_features[6074] ,
    \all_features[6075] , \all_features[6076] , \all_features[6077] ,
    \all_features[6078] , \all_features[6079] , \all_features[6080] ,
    \all_features[6081] , \all_features[6082] , \all_features[6083] ,
    \all_features[6084] , \all_features[6085] , \all_features[6086] ,
    \all_features[6087] , \all_features[6088] , \all_features[6089] ,
    \all_features[6090] , \all_features[6091] , \all_features[6092] ,
    \all_features[6093] , \all_features[6094] , \all_features[6095] ,
    \all_features[6096] , \all_features[6097] , \all_features[6098] ,
    \all_features[6099] , \all_features[6100] , \all_features[6101] ,
    \all_features[6102] , \all_features[6103] , \all_features[6104] ,
    \all_features[6105] , \all_features[6106] , \all_features[6107] ,
    \all_features[6108] , \all_features[6109] , \all_features[6110] ,
    \all_features[6111] , \all_features[6112] , \all_features[6113] ,
    \all_features[6114] , \all_features[6115] , \all_features[6116] ,
    \all_features[6117] , \all_features[6118] , \all_features[6119] ,
    \all_features[6120] , \all_features[6121] , \all_features[6122] ,
    \all_features[6123] , \all_features[6124] , \all_features[6125] ,
    \all_features[6126] , \all_features[6127] , \all_features[6128] ,
    \all_features[6129] , \all_features[6130] , \all_features[6131] ,
    \all_features[6132] , \all_features[6133] , \all_features[6134] ,
    \all_features[6135] , \all_features[6136] , \all_features[6137] ,
    \all_features[6138] , \all_features[6139] , \all_features[6140] ,
    \all_features[6141] , \all_features[6142] , \all_features[6143] ,
    \all_features[6144] , \all_features[6145] , \all_features[6146] ,
    \all_features[6147] , \all_features[6148] , \all_features[6149] ,
    \all_features[6150] , \all_features[6151] , \all_features[6152] ,
    \all_features[6153] , \all_features[6154] , \all_features[6155] ,
    \all_features[6156] , \all_features[6157] , \all_features[6158] ,
    \all_features[6159] , \all_features[6160] , \all_features[6161] ,
    \all_features[6162] , \all_features[6163] , \all_features[6164] ,
    \all_features[6165] , \all_features[6166] , \all_features[6167] ,
    \all_features[6168] , \all_features[6169] , \all_features[6170] ,
    \all_features[6171] , \all_features[6172] , \all_features[6173] ,
    \all_features[6174] , \all_features[6175] , \all_features[6176] ,
    \all_features[6177] , \all_features[6178] , \all_features[6179] ,
    \all_features[6180] , \all_features[6181] , \all_features[6182] ,
    \all_features[6183] , \all_features[6184] , \all_features[6185] ,
    \all_features[6186] , \all_features[6187] , \all_features[6188] ,
    \all_features[6189] , \all_features[6190] , \all_features[6191] ,
    \all_features[6192] , \all_features[6193] , \all_features[6194] ,
    \all_features[6195] , \all_features[6196] , \all_features[6197] ,
    \all_features[6198] , \all_features[6199] , \all_features[6200] ,
    \all_features[6201] , \all_features[6202] , \all_features[6203] ,
    \all_features[6204] , \all_features[6205] , \all_features[6206] ,
    \all_features[6207] , \all_features[6208] , \all_features[6209] ,
    \all_features[6210] , \all_features[6211] , \all_features[6212] ,
    \all_features[6213] , \all_features[6214] , \all_features[6215] ,
    \all_features[6216] , \all_features[6217] , \all_features[6218] ,
    \all_features[6219] , \all_features[6220] , \all_features[6221] ,
    \all_features[6222] , \all_features[6223] , \all_features[6224] ,
    \all_features[6225] , \all_features[6226] , \all_features[6227] ,
    \all_features[6228] , \all_features[6229] , \all_features[6230] ,
    \all_features[6231] , \all_features[6232] , \all_features[6233] ,
    \all_features[6234] , \all_features[6235] , \all_features[6236] ,
    \all_features[6237] , \all_features[6238] , \all_features[6239] ,
    \all_features[6240] , \all_features[6241] , \all_features[6242] ,
    \all_features[6243] , \all_features[6244] , \all_features[6245] ,
    \all_features[6246] , \all_features[6247] , \all_features[6248] ,
    \all_features[6249] , \all_features[6250] , \all_features[6251] ,
    \all_features[6252] , \all_features[6253] , \all_features[6254] ,
    \all_features[6255] , \all_features[6256] , \all_features[6257] ,
    \all_features[6258] , \all_features[6259] , \all_features[6260] ,
    \all_features[6261] , \all_features[6262] , \all_features[6263] ,
    \all_features[6264] , \all_features[6265] , \all_features[6266] ,
    \all_features[6267] , \all_features[6268] , \all_features[6269] ,
    \all_features[6270] , \all_features[6271] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] ,
    \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] ,
    \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] ,
    \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] ,
    \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] ,
    \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] ,
    \o[64] , \o[65] , \o[66] , \o[67] , \o[68] , \o[69] ;
  wire new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_,
    new_n6590_, new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_,
    new_n6596_, new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_,
    new_n6602_, new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_,
    new_n6608_, new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_,
    new_n6614_, new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_,
    new_n6620_, new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_,
    new_n6626_, new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_,
    new_n6632_, new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_,
    new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_,
    new_n6644_, new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_,
    new_n6650_, new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_,
    new_n6656_, new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_,
    new_n6662_, new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_,
    new_n6668_, new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_,
    new_n6674_, new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_,
    new_n6680_, new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_,
    new_n6686_, new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_,
    new_n6692_, new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_,
    new_n6698_, new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_,
    new_n6704_, new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_,
    new_n6710_, new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_,
    new_n6716_, new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_,
    new_n6722_, new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_,
    new_n6728_, new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_,
    new_n6734_, new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_,
    new_n6740_, new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_,
    new_n6746_, new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_,
    new_n6752_, new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_,
    new_n6758_, new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_,
    new_n6764_, new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_,
    new_n6770_, new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_,
    new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_,
    new_n6782_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_,
    new_n7304_, new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_,
    new_n7310_, new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_,
    new_n7316_, new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_,
    new_n7322_, new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_,
    new_n7328_, new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_,
    new_n7334_, new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_,
    new_n7340_, new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_,
    new_n7346_, new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_,
    new_n7352_, new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_,
    new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_,
    new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_,
    new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7375_,
    new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_, new_n7381_,
    new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_, new_n7387_,
    new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_, new_n7393_,
    new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_, new_n7399_,
    new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_, new_n7405_,
    new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_, new_n7411_,
    new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_, new_n7417_,
    new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_, new_n7423_,
    new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_, new_n7429_,
    new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_, new_n7435_,
    new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_, new_n7441_,
    new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_, new_n7447_,
    new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_, new_n7453_,
    new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_, new_n7459_,
    new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_, new_n7465_,
    new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_, new_n7471_,
    new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_, new_n7477_,
    new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_, new_n7483_,
    new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_, new_n7489_,
    new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_, new_n7495_,
    new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_, new_n7501_,
    new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_, new_n7507_,
    new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_, new_n7513_,
    new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_, new_n7519_,
    new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_, new_n7525_,
    new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_, new_n7531_,
    new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_, new_n7537_,
    new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_, new_n7543_,
    new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7762_, new_n7763_, new_n7764_, new_n7765_,
    new_n7766_, new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_,
    new_n7772_, new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_,
    new_n7778_, new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_,
    new_n7784_, new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_,
    new_n7790_, new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_,
    new_n7796_, new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_,
    new_n7802_, new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_,
    new_n7808_, new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_,
    new_n7814_, new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_,
    new_n7820_, new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_,
    new_n7826_, new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_,
    new_n7832_, new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_,
    new_n7838_, new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_,
    new_n7844_, new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_,
    new_n7850_, new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_,
    new_n7856_, new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_,
    new_n7862_, new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_,
    new_n7868_, new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_,
    new_n7874_, new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_,
    new_n7880_, new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_,
    new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_,
    new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_,
    new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_,
    new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_,
    new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_,
    new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_,
    new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_,
    new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_,
    new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_,
    new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_,
    new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_,
    new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_,
    new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_, new_n7963_,
    new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_, new_n7969_,
    new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_, new_n7975_,
    new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_, new_n7981_,
    new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_, new_n7987_,
    new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_, new_n7993_,
    new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_, new_n7999_,
    new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_, new_n8005_,
    new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_, new_n8011_,
    new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_, new_n8017_,
    new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_, new_n8023_,
    new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_, new_n8029_,
    new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_, new_n8035_,
    new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_, new_n8041_,
    new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_, new_n8047_,
    new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_,
    new_n8216_, new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_,
    new_n8222_, new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_,
    new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_,
    new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_,
    new_n8240_, new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_,
    new_n8252_, new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_,
    new_n8258_, new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_,
    new_n8264_, new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_,
    new_n8270_, new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_,
    new_n8276_, new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_,
    new_n8282_, new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_,
    new_n8288_, new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_,
    new_n8294_, new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_,
    new_n8300_, new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_,
    new_n8306_, new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_,
    new_n8312_, new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_,
    new_n8318_, new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_,
    new_n8324_, new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_,
    new_n8330_, new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_,
    new_n8336_, new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_,
    new_n8342_, new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_,
    new_n8348_, new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_,
    new_n8354_, new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_,
    new_n8360_, new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_,
    new_n8366_, new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8371_,
    new_n8372_, new_n8373_, new_n8374_, new_n8375_, new_n8376_, new_n8377_,
    new_n8378_, new_n8379_, new_n8380_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8389_,
    new_n8390_, new_n8391_, new_n8392_, new_n8393_, new_n8394_, new_n8395_,
    new_n8396_, new_n8397_, new_n8398_, new_n8399_, new_n8400_, new_n8401_,
    new_n8402_, new_n8403_, new_n8404_, new_n8405_, new_n8406_, new_n8407_,
    new_n8408_, new_n8409_, new_n8410_, new_n8411_, new_n8412_, new_n8413_,
    new_n8414_, new_n8415_, new_n8416_, new_n8417_, new_n8418_, new_n8419_,
    new_n8420_, new_n8421_, new_n8422_, new_n8423_, new_n8424_, new_n8425_,
    new_n8426_, new_n8427_, new_n8428_, new_n8429_, new_n8430_, new_n8431_,
    new_n8432_, new_n8433_, new_n8434_, new_n8435_, new_n8436_, new_n8437_,
    new_n8438_, new_n8439_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8448_, new_n8449_,
    new_n8450_, new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_,
    new_n8456_, new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8461_,
    new_n8462_, new_n8463_, new_n8464_, new_n8465_, new_n8466_, new_n8467_,
    new_n8468_, new_n8469_, new_n8470_, new_n8471_, new_n8472_, new_n8473_,
    new_n8474_, new_n8475_, new_n8476_, new_n8477_, new_n8478_, new_n8479_,
    new_n8480_, new_n8481_, new_n8482_, new_n8483_, new_n8484_, new_n8485_,
    new_n8486_, new_n8487_, new_n8488_, new_n8489_, new_n8490_, new_n8491_,
    new_n8492_, new_n8493_, new_n8494_, new_n8495_, new_n8496_, new_n8497_,
    new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_, new_n8503_,
    new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_, new_n8515_,
    new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_,
    new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_,
    new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_,
    new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_,
    new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_,
    new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_,
    new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_,
    new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_,
    new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_,
    new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_,
    new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_,
    new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_,
    new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_,
    new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_,
    new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_,
    new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_,
    new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_,
    new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_,
    new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_,
    new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_,
    new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_,
    new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_,
    new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_,
    new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_,
    new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_,
    new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_,
    new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_, new_n8959_,
    new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_,
    new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_,
    new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_,
    new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_,
    new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_,
    new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_,
    new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_,
    new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_,
    new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_,
    new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_,
    new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_,
    new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_,
    new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_,
    new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_,
    new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_,
    new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_, new_n9289_,
    new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_, new_n9295_,
    new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_, new_n9301_,
    new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_, new_n9307_,
    new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_, new_n9313_,
    new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_, new_n9319_,
    new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_, new_n9325_,
    new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_, new_n9331_,
    new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_, new_n9337_,
    new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_, new_n9343_,
    new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_, new_n9349_,
    new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_, new_n9355_,
    new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_, new_n9361_,
    new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_, new_n9367_,
    new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_, new_n9373_,
    new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_, new_n9379_,
    new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_, new_n9385_,
    new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_, new_n9391_,
    new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_, new_n9397_,
    new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_, new_n9403_,
    new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_, new_n9409_,
    new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_, new_n9415_,
    new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_, new_n9421_,
    new_n9422_, new_n9423_, new_n9424_, new_n9425_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9432_, new_n9433_,
    new_n9434_, new_n9435_, new_n9436_, new_n9437_, new_n9438_, new_n9439_,
    new_n9440_, new_n9441_, new_n9442_, new_n9443_, new_n9444_, new_n9445_,
    new_n9446_, new_n9447_, new_n9448_, new_n9449_, new_n9450_, new_n9451_,
    new_n9452_, new_n9453_, new_n9454_, new_n9455_, new_n9456_, new_n9457_,
    new_n9458_, new_n9459_, new_n9460_, new_n9461_, new_n9462_, new_n9463_,
    new_n9464_, new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_,
    new_n9470_, new_n9471_, new_n9472_, new_n9473_, new_n9474_, new_n9475_,
    new_n9476_, new_n9477_, new_n9478_, new_n9479_, new_n9480_, new_n9481_,
    new_n9482_, new_n9483_, new_n9484_, new_n9485_, new_n9486_, new_n9487_,
    new_n9488_, new_n9489_, new_n9490_, new_n9491_, new_n9492_, new_n9493_,
    new_n9494_, new_n9495_, new_n9496_, new_n9497_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9502_, new_n9503_, new_n9504_, new_n9505_,
    new_n9506_, new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9511_,
    new_n9512_, new_n9513_, new_n9514_, new_n9515_, new_n9516_, new_n9517_,
    new_n9518_, new_n9519_, new_n9520_, new_n9521_, new_n9522_, new_n9523_,
    new_n9524_, new_n9525_, new_n9526_, new_n9527_, new_n9528_, new_n9529_,
    new_n9530_, new_n9531_, new_n9532_, new_n9533_, new_n9534_, new_n9535_,
    new_n9536_, new_n9537_, new_n9538_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9589_,
    new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_,
    new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9601_,
    new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_, new_n9607_,
    new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_, new_n9613_,
    new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_, new_n9619_,
    new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_, new_n9625_,
    new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_, new_n9631_,
    new_n9632_, new_n9633_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_,
    new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_,
    new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_,
    new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_,
    new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_,
    new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_,
    new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_,
    new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_,
    new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_,
    new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9956_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11602_,
    new_n11603_, new_n11604_, new_n11605_, new_n11606_, new_n11607_,
    new_n11608_, new_n11609_, new_n11610_, new_n11611_, new_n11612_,
    new_n11613_, new_n11614_, new_n11615_, new_n11616_, new_n11617_,
    new_n11618_, new_n11619_, new_n11620_, new_n11621_, new_n11622_,
    new_n11623_, new_n11624_, new_n11625_, new_n11626_, new_n11627_,
    new_n11628_, new_n11629_, new_n11630_, new_n11631_, new_n11632_,
    new_n11633_, new_n11634_, new_n11635_, new_n11636_, new_n11637_,
    new_n11638_, new_n11639_, new_n11640_, new_n11641_, new_n11642_,
    new_n11643_, new_n11644_, new_n11645_, new_n11646_, new_n11647_,
    new_n11648_, new_n11649_, new_n11650_, new_n11651_, new_n11652_,
    new_n11653_, new_n11654_, new_n11655_, new_n11656_, new_n11657_,
    new_n11658_, new_n11659_, new_n11660_, new_n11661_, new_n11662_,
    new_n11663_, new_n11664_, new_n11665_, new_n11666_, new_n11667_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11732_,
    new_n11733_, new_n11734_, new_n11735_, new_n11736_, new_n11737_,
    new_n11738_, new_n11739_, new_n11740_, new_n11741_, new_n11742_,
    new_n11743_, new_n11744_, new_n11745_, new_n11746_, new_n11747_,
    new_n11748_, new_n11749_, new_n11750_, new_n11751_, new_n11752_,
    new_n11753_, new_n11754_, new_n11755_, new_n11756_, new_n11757_,
    new_n11758_, new_n11759_, new_n11760_, new_n11761_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11804_, new_n11805_, new_n11806_, new_n11807_,
    new_n11808_, new_n11809_, new_n11810_, new_n11811_, new_n11812_,
    new_n11813_, new_n11814_, new_n11815_, new_n11816_, new_n11817_,
    new_n11818_, new_n11819_, new_n11820_, new_n11821_, new_n11822_,
    new_n11823_, new_n11824_, new_n11825_, new_n11826_, new_n11827_,
    new_n11828_, new_n11829_, new_n11830_, new_n11831_, new_n11832_,
    new_n11833_, new_n11834_, new_n11835_, new_n11836_, new_n11837_,
    new_n11838_, new_n11839_, new_n11840_, new_n11841_, new_n11842_,
    new_n11843_, new_n11844_, new_n11845_, new_n11846_, new_n11847_,
    new_n11848_, new_n11849_, new_n11850_, new_n11851_, new_n11852_,
    new_n11853_, new_n11854_, new_n11855_, new_n11856_, new_n11857_,
    new_n11858_, new_n11859_, new_n11860_, new_n11861_, new_n11862_,
    new_n11863_, new_n11864_, new_n11865_, new_n11866_, new_n11867_,
    new_n11868_, new_n11869_, new_n11870_, new_n11871_, new_n11872_,
    new_n11873_, new_n11874_, new_n11875_, new_n11876_, new_n11877_,
    new_n11878_, new_n11879_, new_n11880_, new_n11881_, new_n11882_,
    new_n11883_, new_n11884_, new_n11885_, new_n11886_, new_n11887_,
    new_n11888_, new_n11889_, new_n11890_, new_n11891_, new_n11892_,
    new_n11893_, new_n11894_, new_n11895_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12008_, new_n12009_, new_n12010_, new_n12011_, new_n12012_,
    new_n12013_, new_n12014_, new_n12015_, new_n12016_, new_n12017_,
    new_n12018_, new_n12019_, new_n12020_, new_n12021_, new_n12022_,
    new_n12023_, new_n12024_, new_n12025_, new_n12026_, new_n12027_,
    new_n12028_, new_n12029_, new_n12030_, new_n12031_, new_n12032_,
    new_n12033_, new_n12034_, new_n12035_, new_n12036_, new_n12037_,
    new_n12038_, new_n12039_, new_n12040_, new_n12041_, new_n12042_,
    new_n12043_, new_n12044_, new_n12045_, new_n12046_, new_n12047_,
    new_n12048_, new_n12049_, new_n12050_, new_n12051_, new_n12052_,
    new_n12053_, new_n12054_, new_n12055_, new_n12056_, new_n12057_,
    new_n12058_, new_n12059_, new_n12060_, new_n12061_, new_n12062_,
    new_n12063_, new_n12064_, new_n12065_, new_n12066_, new_n12067_,
    new_n12068_, new_n12069_, new_n12070_, new_n12071_, new_n12072_,
    new_n12073_, new_n12074_, new_n12075_, new_n12076_, new_n12077_,
    new_n12078_, new_n12079_, new_n12080_, new_n12081_, new_n12082_,
    new_n12083_, new_n12084_, new_n12085_, new_n12086_, new_n12087_,
    new_n12088_, new_n12089_, new_n12090_, new_n12091_, new_n12092_,
    new_n12093_, new_n12094_, new_n12095_, new_n12096_, new_n12097_,
    new_n12098_, new_n12099_, new_n12100_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12226_, new_n12227_,
    new_n12228_, new_n12229_, new_n12230_, new_n12231_, new_n12232_,
    new_n12233_, new_n12234_, new_n12235_, new_n12236_, new_n12237_,
    new_n12238_, new_n12239_, new_n12240_, new_n12241_, new_n12242_,
    new_n12243_, new_n12244_, new_n12245_, new_n12246_, new_n12247_,
    new_n12248_, new_n12249_, new_n12250_, new_n12251_, new_n12252_,
    new_n12253_, new_n12254_, new_n12255_, new_n12256_, new_n12257_,
    new_n12258_, new_n12259_, new_n12260_, new_n12261_, new_n12262_,
    new_n12263_, new_n12264_, new_n12265_, new_n12266_, new_n12267_,
    new_n12268_, new_n12269_, new_n12270_, new_n12271_, new_n12272_,
    new_n12273_, new_n12274_, new_n12275_, new_n12276_, new_n12277_,
    new_n12278_, new_n12279_, new_n12280_, new_n12281_, new_n12282_,
    new_n12283_, new_n12284_, new_n12285_, new_n12286_, new_n12287_,
    new_n12288_, new_n12289_, new_n12290_, new_n12291_, new_n12292_,
    new_n12293_, new_n12294_, new_n12295_, new_n12296_, new_n12297_,
    new_n12298_, new_n12299_, new_n12300_, new_n12301_, new_n12302_,
    new_n12303_, new_n12304_, new_n12305_, new_n12306_, new_n12307_,
    new_n12308_, new_n12309_, new_n12310_, new_n12311_, new_n12312_,
    new_n12313_, new_n12314_, new_n12315_, new_n12316_, new_n12317_,
    new_n12318_, new_n12319_, new_n12320_, new_n12321_, new_n12322_,
    new_n12323_, new_n12324_, new_n12325_, new_n12326_, new_n12327_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12417_,
    new_n12418_, new_n12419_, new_n12420_, new_n12421_, new_n12422_,
    new_n12423_, new_n12424_, new_n12425_, new_n12426_, new_n12427_,
    new_n12428_, new_n12429_, new_n12430_, new_n12431_, new_n12432_,
    new_n12433_, new_n12434_, new_n12435_, new_n12436_, new_n12437_,
    new_n12438_, new_n12439_, new_n12440_, new_n12441_, new_n12442_,
    new_n12443_, new_n12444_, new_n12445_, new_n12446_, new_n12447_,
    new_n12448_, new_n12449_, new_n12450_, new_n12451_, new_n12452_,
    new_n12453_, new_n12454_, new_n12455_, new_n12456_, new_n12457_,
    new_n12458_, new_n12459_, new_n12460_, new_n12461_, new_n12462_,
    new_n12463_, new_n12464_, new_n12465_, new_n12466_, new_n12467_,
    new_n12468_, new_n12469_, new_n12470_, new_n12471_, new_n12472_,
    new_n12473_, new_n12474_, new_n12475_, new_n12476_, new_n12477_,
    new_n12478_, new_n12479_, new_n12480_, new_n12481_, new_n12482_,
    new_n12483_, new_n12484_, new_n12485_, new_n12486_, new_n12487_,
    new_n12488_, new_n12489_, new_n12490_, new_n12491_, new_n12492_,
    new_n12493_, new_n12494_, new_n12495_, new_n12496_, new_n12497_,
    new_n12498_, new_n12499_, new_n12500_, new_n12501_, new_n12502_,
    new_n12503_, new_n12504_, new_n12505_, new_n12506_, new_n12507_,
    new_n12508_, new_n12509_, new_n12510_, new_n12511_, new_n12512_,
    new_n12513_, new_n12514_, new_n12515_, new_n12516_, new_n12517_,
    new_n12518_, new_n12519_, new_n12520_, new_n12521_, new_n12522_,
    new_n12523_, new_n12524_, new_n12525_, new_n12526_, new_n12527_,
    new_n12528_, new_n12529_, new_n12530_, new_n12531_, new_n12532_,
    new_n12533_, new_n12534_, new_n12535_, new_n12536_, new_n12537_,
    new_n12538_, new_n12539_, new_n12540_, new_n12541_, new_n12542_,
    new_n12543_, new_n12544_, new_n12545_, new_n12546_, new_n12547_,
    new_n12548_, new_n12549_, new_n12550_, new_n12551_, new_n12552_,
    new_n12553_, new_n12554_, new_n12555_, new_n12556_, new_n12557_,
    new_n12558_, new_n12559_, new_n12560_, new_n12561_, new_n12562_,
    new_n12563_, new_n12564_, new_n12565_, new_n12566_, new_n12567_,
    new_n12568_, new_n12569_, new_n12570_, new_n12571_, new_n12572_,
    new_n12573_, new_n12574_, new_n12575_, new_n12576_, new_n12577_,
    new_n12578_, new_n12579_, new_n12580_, new_n12581_, new_n12582_,
    new_n12583_, new_n12584_, new_n12585_, new_n12586_, new_n12587_,
    new_n12588_, new_n12589_, new_n12590_, new_n12591_, new_n12592_,
    new_n12593_, new_n12594_, new_n12595_, new_n12596_, new_n12597_,
    new_n12598_, new_n12599_, new_n12600_, new_n12601_, new_n12602_,
    new_n12603_, new_n12604_, new_n12605_, new_n12606_, new_n12607_,
    new_n12608_, new_n12609_, new_n12610_, new_n12611_, new_n12612_,
    new_n12613_, new_n12614_, new_n12615_, new_n12616_, new_n12617_,
    new_n12618_, new_n12619_, new_n12620_, new_n12621_, new_n12622_,
    new_n12623_, new_n12624_, new_n12625_, new_n12626_, new_n12627_,
    new_n12628_, new_n12629_, new_n12630_, new_n12631_, new_n12632_,
    new_n12633_, new_n12634_, new_n12635_, new_n12636_, new_n12637_,
    new_n12638_, new_n12639_, new_n12640_, new_n12641_, new_n12642_,
    new_n12643_, new_n12644_, new_n12645_, new_n12646_, new_n12647_,
    new_n12648_, new_n12649_, new_n12650_, new_n12651_, new_n12652_,
    new_n12653_, new_n12654_, new_n12655_, new_n12656_, new_n12657_,
    new_n12658_, new_n12659_, new_n12660_, new_n12661_, new_n12662_,
    new_n12663_, new_n12664_, new_n12665_, new_n12666_, new_n12667_,
    new_n12668_, new_n12669_, new_n12670_, new_n12671_, new_n12672_,
    new_n12673_, new_n12674_, new_n12675_, new_n12676_, new_n12677_,
    new_n12678_, new_n12679_, new_n12680_, new_n12681_, new_n12682_,
    new_n12683_, new_n12684_, new_n12685_, new_n12686_, new_n12687_,
    new_n12688_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12801_, new_n12802_,
    new_n12803_, new_n12804_, new_n12805_, new_n12806_, new_n12807_,
    new_n12808_, new_n12809_, new_n12810_, new_n12811_, new_n12812_,
    new_n12813_, new_n12814_, new_n12815_, new_n12816_, new_n12817_,
    new_n12818_, new_n12819_, new_n12820_, new_n12821_, new_n12822_,
    new_n12823_, new_n12824_, new_n12825_, new_n12826_, new_n12827_,
    new_n12828_, new_n12829_, new_n12830_, new_n12831_, new_n12832_,
    new_n12833_, new_n12834_, new_n12835_, new_n12836_, new_n12837_,
    new_n12838_, new_n12839_, new_n12840_, new_n12841_, new_n12842_,
    new_n12843_, new_n12844_, new_n12845_, new_n12846_, new_n12847_,
    new_n12848_, new_n12849_, new_n12850_, new_n12851_, new_n12852_,
    new_n12853_, new_n12854_, new_n12855_, new_n12856_, new_n12857_,
    new_n12858_, new_n12859_, new_n12860_, new_n12861_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12900_, new_n12901_, new_n12902_, new_n12903_,
    new_n12904_, new_n12905_, new_n12906_, new_n12907_, new_n12908_,
    new_n12909_, new_n12910_, new_n12911_, new_n12912_, new_n12913_,
    new_n12914_, new_n12915_, new_n12916_, new_n12917_, new_n12918_,
    new_n12919_, new_n12920_, new_n12921_, new_n12922_, new_n12923_,
    new_n12924_, new_n12925_, new_n12926_, new_n12927_, new_n12928_,
    new_n12929_, new_n12930_, new_n12931_, new_n12932_, new_n12933_,
    new_n12934_, new_n12935_, new_n12936_, new_n12937_, new_n12938_,
    new_n12939_, new_n12940_, new_n12941_, new_n12942_, new_n12943_,
    new_n12944_, new_n12945_, new_n12946_, new_n12947_, new_n12948_,
    new_n12949_, new_n12950_, new_n12951_, new_n12952_, new_n12953_,
    new_n12954_, new_n12955_, new_n12956_, new_n12957_, new_n12958_,
    new_n12959_, new_n12960_, new_n12961_, new_n12962_, new_n12963_,
    new_n12964_, new_n12965_, new_n12966_, new_n12967_, new_n12968_,
    new_n12969_, new_n12970_, new_n12971_, new_n12972_, new_n12973_,
    new_n12974_, new_n12975_, new_n12976_, new_n12977_, new_n12978_,
    new_n12979_, new_n12980_, new_n12981_, new_n12982_, new_n12983_,
    new_n12984_, new_n12985_, new_n12986_, new_n12987_, new_n12988_,
    new_n12989_, new_n12990_, new_n12991_, new_n12992_, new_n12993_,
    new_n12994_, new_n12995_, new_n12996_, new_n12997_, new_n12998_,
    new_n12999_, new_n13000_, new_n13001_, new_n13002_, new_n13003_,
    new_n13004_, new_n13005_, new_n13006_, new_n13007_, new_n13008_,
    new_n13009_, new_n13010_, new_n13011_, new_n13012_, new_n13013_,
    new_n13014_, new_n13015_, new_n13016_, new_n13017_, new_n13018_,
    new_n13019_, new_n13020_, new_n13021_, new_n13022_, new_n13023_,
    new_n13024_, new_n13025_, new_n13026_, new_n13027_, new_n13028_,
    new_n13029_, new_n13030_, new_n13031_, new_n13032_, new_n13033_,
    new_n13034_, new_n13035_, new_n13036_, new_n13037_, new_n13038_,
    new_n13039_, new_n13040_, new_n13041_, new_n13042_, new_n13043_,
    new_n13044_, new_n13045_, new_n13046_, new_n13047_, new_n13048_,
    new_n13049_, new_n13050_, new_n13051_, new_n13052_, new_n13053_,
    new_n13054_, new_n13055_, new_n13056_, new_n13057_, new_n13058_,
    new_n13059_, new_n13060_, new_n13061_, new_n13062_, new_n13063_,
    new_n13064_, new_n13065_, new_n13066_, new_n13067_, new_n13068_,
    new_n13069_, new_n13070_, new_n13071_, new_n13072_, new_n13073_,
    new_n13074_, new_n13075_, new_n13076_, new_n13077_, new_n13078_,
    new_n13079_, new_n13080_, new_n13081_, new_n13082_, new_n13083_,
    new_n13084_, new_n13085_, new_n13086_, new_n13087_, new_n13088_,
    new_n13089_, new_n13090_, new_n13091_, new_n13092_, new_n13093_,
    new_n13094_, new_n13095_, new_n13096_, new_n13097_, new_n13098_,
    new_n13099_, new_n13100_, new_n13101_, new_n13102_, new_n13103_,
    new_n13104_, new_n13105_, new_n13106_, new_n13107_, new_n13108_,
    new_n13109_, new_n13110_, new_n13111_, new_n13112_, new_n13113_,
    new_n13114_, new_n13115_, new_n13116_, new_n13117_, new_n13118_,
    new_n13119_, new_n13120_, new_n13121_, new_n13122_, new_n13123_,
    new_n13124_, new_n13125_, new_n13126_, new_n13127_, new_n13128_,
    new_n13129_, new_n13130_, new_n13131_, new_n13132_, new_n13133_,
    new_n13134_, new_n13135_, new_n13136_, new_n13137_, new_n13138_,
    new_n13139_, new_n13140_, new_n13141_, new_n13142_, new_n13143_,
    new_n13144_, new_n13145_, new_n13146_, new_n13147_, new_n13148_,
    new_n13149_, new_n13150_, new_n13151_, new_n13152_, new_n13153_,
    new_n13154_, new_n13155_, new_n13156_, new_n13157_, new_n13158_,
    new_n13159_, new_n13160_, new_n13161_, new_n13162_, new_n13163_,
    new_n13164_, new_n13165_, new_n13166_, new_n13167_, new_n13168_,
    new_n13169_, new_n13170_, new_n13171_, new_n13172_, new_n13173_,
    new_n13174_, new_n13175_, new_n13176_, new_n13177_, new_n13178_,
    new_n13179_, new_n13180_, new_n13181_, new_n13182_, new_n13183_,
    new_n13184_, new_n13185_, new_n13186_, new_n13187_, new_n13188_,
    new_n13189_, new_n13190_, new_n13191_, new_n13192_, new_n13193_,
    new_n13194_, new_n13195_, new_n13196_, new_n13197_, new_n13198_,
    new_n13199_, new_n13200_, new_n13201_, new_n13202_, new_n13203_,
    new_n13204_, new_n13205_, new_n13206_, new_n13207_, new_n13208_,
    new_n13209_, new_n13210_, new_n13211_, new_n13212_, new_n13213_,
    new_n13214_, new_n13215_, new_n13216_, new_n13217_, new_n13218_,
    new_n13219_, new_n13220_, new_n13221_, new_n13222_, new_n13223_,
    new_n13224_, new_n13225_, new_n13226_, new_n13227_, new_n13228_,
    new_n13229_, new_n13230_, new_n13231_, new_n13232_, new_n13233_,
    new_n13234_, new_n13235_, new_n13236_, new_n13237_, new_n13238_,
    new_n13239_, new_n13240_, new_n13241_, new_n13242_, new_n13243_,
    new_n13244_, new_n13245_, new_n13246_, new_n13247_, new_n13248_,
    new_n13249_, new_n13250_, new_n13251_, new_n13252_, new_n13253_,
    new_n13254_, new_n13255_, new_n13256_, new_n13257_, new_n13258_,
    new_n13259_, new_n13260_, new_n13261_, new_n13262_, new_n13263_,
    new_n13264_, new_n13265_, new_n13266_, new_n13267_, new_n13268_,
    new_n13269_, new_n13270_, new_n13271_, new_n13272_, new_n13273_,
    new_n13274_, new_n13275_, new_n13276_, new_n13277_, new_n13278_,
    new_n13279_, new_n13280_, new_n13281_, new_n13282_, new_n13283_,
    new_n13284_, new_n13285_, new_n13286_, new_n13287_, new_n13288_,
    new_n13289_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13380_, new_n13381_, new_n13382_, new_n13383_,
    new_n13384_, new_n13385_, new_n13386_, new_n13387_, new_n13388_,
    new_n13389_, new_n13390_, new_n13391_, new_n13392_, new_n13393_,
    new_n13394_, new_n13395_, new_n13396_, new_n13397_, new_n13398_,
    new_n13399_, new_n13400_, new_n13401_, new_n13402_, new_n13403_,
    new_n13404_, new_n13405_, new_n13406_, new_n13407_, new_n13408_,
    new_n13409_, new_n13410_, new_n13411_, new_n13412_, new_n13413_,
    new_n13414_, new_n13415_, new_n13416_, new_n13417_, new_n13418_,
    new_n13419_, new_n13420_, new_n13421_, new_n13422_, new_n13423_,
    new_n13424_, new_n13425_, new_n13426_, new_n13427_, new_n13428_,
    new_n13429_, new_n13430_, new_n13431_, new_n13432_, new_n13433_,
    new_n13434_, new_n13435_, new_n13436_, new_n13437_, new_n13438_,
    new_n13439_, new_n13440_, new_n13441_, new_n13442_, new_n13443_,
    new_n13444_, new_n13445_, new_n13446_, new_n13447_, new_n13448_,
    new_n13449_, new_n13450_, new_n13451_, new_n13452_, new_n13453_,
    new_n13454_, new_n13455_, new_n13456_, new_n13457_, new_n13458_,
    new_n13459_, new_n13460_, new_n13461_, new_n13462_, new_n13463_,
    new_n13464_, new_n13465_, new_n13466_, new_n13467_, new_n13468_,
    new_n13469_, new_n13470_, new_n13471_, new_n13472_, new_n13473_,
    new_n13474_, new_n13475_, new_n13476_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13648_, new_n13649_, new_n13650_, new_n13652_, new_n13653_,
    new_n13654_, new_n13655_, new_n13656_, new_n13657_, new_n13659_,
    new_n13660_, new_n13661_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13831_,
    new_n13832_, new_n13833_, new_n13834_, new_n13835_, new_n13836_,
    new_n13837_, new_n13838_, new_n13839_, new_n13840_, new_n13841_,
    new_n13842_, new_n13843_, new_n13844_, new_n13845_, new_n13846_,
    new_n13847_, new_n13848_, new_n13849_, new_n13850_, new_n13851_,
    new_n13852_, new_n13853_, new_n13854_, new_n13855_, new_n13856_,
    new_n13857_, new_n13858_, new_n13859_, new_n13860_, new_n13861_,
    new_n13862_, new_n13863_, new_n13864_, new_n13865_, new_n13866_,
    new_n13867_, new_n13868_, new_n13869_, new_n13870_, new_n13871_,
    new_n13872_, new_n13873_, new_n13874_, new_n13875_, new_n13876_,
    new_n13877_, new_n13878_, new_n13879_, new_n13880_, new_n13881_,
    new_n13882_, new_n13883_, new_n13884_, new_n13885_, new_n13886_,
    new_n13887_, new_n13888_, new_n13889_, new_n13890_, new_n13891_,
    new_n13892_, new_n13893_, new_n13894_, new_n13895_, new_n13896_,
    new_n13897_, new_n13898_, new_n13899_, new_n13900_, new_n13901_,
    new_n13902_, new_n13903_, new_n13904_, new_n13905_, new_n13906_,
    new_n13907_, new_n13908_, new_n13909_, new_n13910_, new_n13911_,
    new_n13912_, new_n13913_, new_n13914_, new_n13915_, new_n13916_,
    new_n13917_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13979_, new_n13980_, new_n13981_,
    new_n13982_, new_n13983_, new_n13984_, new_n13985_, new_n13986_,
    new_n13987_, new_n13988_, new_n13989_, new_n13990_, new_n13991_,
    new_n13992_, new_n13993_, new_n13994_, new_n13995_, new_n13996_,
    new_n13997_, new_n13998_, new_n13999_, new_n14000_, new_n14001_,
    new_n14002_, new_n14003_, new_n14004_, new_n14005_, new_n14006_,
    new_n14007_, new_n14008_, new_n14009_, new_n14010_, new_n14011_,
    new_n14012_, new_n14013_, new_n14014_, new_n14015_, new_n14016_,
    new_n14017_, new_n14018_, new_n14019_, new_n14020_, new_n14021_,
    new_n14022_, new_n14023_, new_n14024_, new_n14025_, new_n14026_,
    new_n14027_, new_n14028_, new_n14029_, new_n14030_, new_n14031_,
    new_n14032_, new_n14033_, new_n14034_, new_n14035_, new_n14036_,
    new_n14037_, new_n14038_, new_n14039_, new_n14040_, new_n14041_,
    new_n14042_, new_n14043_, new_n14044_, new_n14045_, new_n14046_,
    new_n14047_, new_n14048_, new_n14049_, new_n14050_, new_n14051_,
    new_n14052_, new_n14053_, new_n14054_, new_n14055_, new_n14056_,
    new_n14057_, new_n14058_, new_n14059_, new_n14060_, new_n14061_,
    new_n14062_, new_n14063_, new_n14064_, new_n14065_, new_n14066_,
    new_n14067_, new_n14068_, new_n14069_, new_n14070_, new_n14071_,
    new_n14072_, new_n14073_, new_n14074_, new_n14075_, new_n14076_,
    new_n14077_, new_n14078_, new_n14079_, new_n14080_, new_n14081_,
    new_n14082_, new_n14083_, new_n14084_, new_n14085_, new_n14086_,
    new_n14087_, new_n14088_, new_n14089_, new_n14090_, new_n14091_,
    new_n14092_, new_n14093_, new_n14094_, new_n14095_, new_n14096_,
    new_n14097_, new_n14098_, new_n14099_, new_n14100_, new_n14101_,
    new_n14102_, new_n14103_, new_n14104_, new_n14105_, new_n14106_,
    new_n14107_, new_n14108_, new_n14109_, new_n14110_, new_n14111_,
    new_n14112_, new_n14113_, new_n14114_, new_n14115_, new_n14116_,
    new_n14117_, new_n14118_, new_n14119_, new_n14120_, new_n14121_,
    new_n14122_, new_n14123_, new_n14124_, new_n14125_, new_n14126_,
    new_n14127_, new_n14128_, new_n14129_, new_n14130_, new_n14131_,
    new_n14132_, new_n14133_, new_n14134_, new_n14135_, new_n14136_,
    new_n14137_, new_n14138_, new_n14139_, new_n14140_, new_n14141_,
    new_n14142_, new_n14143_, new_n14144_, new_n14145_, new_n14146_,
    new_n14147_, new_n14148_, new_n14149_, new_n14150_, new_n14151_,
    new_n14152_, new_n14153_, new_n14154_, new_n14155_, new_n14156_,
    new_n14157_, new_n14158_, new_n14159_, new_n14160_, new_n14161_,
    new_n14162_, new_n14163_, new_n14164_, new_n14165_, new_n14166_,
    new_n14167_, new_n14168_, new_n14169_, new_n14170_, new_n14171_,
    new_n14172_, new_n14173_, new_n14174_, new_n14175_, new_n14176_,
    new_n14177_, new_n14178_, new_n14179_, new_n14180_, new_n14181_,
    new_n14182_, new_n14183_, new_n14184_, new_n14185_, new_n14186_,
    new_n14187_, new_n14188_, new_n14189_, new_n14190_, new_n14191_,
    new_n14192_, new_n14193_, new_n14194_, new_n14195_, new_n14196_,
    new_n14197_, new_n14198_, new_n14199_, new_n14200_, new_n14201_,
    new_n14202_, new_n14203_, new_n14204_, new_n14205_, new_n14206_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14257_, new_n14258_, new_n14259_, new_n14260_, new_n14261_,
    new_n14262_, new_n14263_, new_n14264_, new_n14265_, new_n14266_,
    new_n14267_, new_n14268_, new_n14269_, new_n14270_, new_n14271_,
    new_n14272_, new_n14273_, new_n14274_, new_n14275_, new_n14276_,
    new_n14277_, new_n14278_, new_n14279_, new_n14280_, new_n14281_,
    new_n14282_, new_n14283_, new_n14284_, new_n14285_, new_n14286_,
    new_n14287_, new_n14288_, new_n14289_, new_n14290_, new_n14291_,
    new_n14292_, new_n14293_, new_n14294_, new_n14295_, new_n14296_,
    new_n14297_, new_n14298_, new_n14299_, new_n14300_, new_n14301_,
    new_n14302_, new_n14303_, new_n14304_, new_n14305_, new_n14306_,
    new_n14307_, new_n14308_, new_n14309_, new_n14310_, new_n14311_,
    new_n14312_, new_n14313_, new_n14314_, new_n14315_, new_n14316_,
    new_n14317_, new_n14318_, new_n14319_, new_n14320_, new_n14321_,
    new_n14322_, new_n14323_, new_n14324_, new_n14325_, new_n14326_,
    new_n14327_, new_n14328_, new_n14329_, new_n14330_, new_n14331_,
    new_n14332_, new_n14333_, new_n14334_, new_n14335_, new_n14336_,
    new_n14337_, new_n14338_, new_n14339_, new_n14340_, new_n14341_,
    new_n14342_, new_n14343_, new_n14344_, new_n14345_, new_n14346_,
    new_n14347_, new_n14348_, new_n14349_, new_n14350_, new_n14351_,
    new_n14352_, new_n14353_, new_n14354_, new_n14355_, new_n14356_,
    new_n14357_, new_n14358_, new_n14359_, new_n14360_, new_n14361_,
    new_n14362_, new_n14363_, new_n14364_, new_n14365_, new_n14366_,
    new_n14367_, new_n14368_, new_n14369_, new_n14370_, new_n14371_,
    new_n14372_, new_n14373_, new_n14374_, new_n14375_, new_n14376_,
    new_n14377_, new_n14378_, new_n14379_, new_n14380_, new_n14381_,
    new_n14382_, new_n14383_, new_n14384_, new_n14385_, new_n14386_,
    new_n14387_, new_n14388_, new_n14389_, new_n14390_, new_n14391_,
    new_n14392_, new_n14393_, new_n14394_, new_n14395_, new_n14396_,
    new_n14397_, new_n14398_, new_n14399_, new_n14400_, new_n14401_,
    new_n14402_, new_n14403_, new_n14404_, new_n14405_, new_n14406_,
    new_n14407_, new_n14408_, new_n14409_, new_n14410_, new_n14411_,
    new_n14412_, new_n14413_, new_n14414_, new_n14415_, new_n14416_,
    new_n14417_, new_n14418_, new_n14419_, new_n14420_, new_n14421_,
    new_n14422_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14455_, new_n14456_,
    new_n14457_, new_n14458_, new_n14459_, new_n14460_, new_n14461_,
    new_n14462_, new_n14463_, new_n14464_, new_n14465_, new_n14466_,
    new_n14467_, new_n14468_, new_n14469_, new_n14470_, new_n14471_,
    new_n14472_, new_n14473_, new_n14474_, new_n14475_, new_n14476_,
    new_n14477_, new_n14478_, new_n14479_, new_n14480_, new_n14481_,
    new_n14482_, new_n14483_, new_n14484_, new_n14485_, new_n14486_,
    new_n14487_, new_n14488_, new_n14489_, new_n14490_, new_n14491_,
    new_n14492_, new_n14493_, new_n14494_, new_n14495_, new_n14496_,
    new_n14497_, new_n14498_, new_n14499_, new_n14500_, new_n14501_,
    new_n14502_, new_n14503_, new_n14504_, new_n14505_, new_n14506_,
    new_n14507_, new_n14508_, new_n14509_, new_n14510_, new_n14511_,
    new_n14512_, new_n14513_, new_n14514_, new_n14515_, new_n14516_,
    new_n14517_, new_n14518_, new_n14519_, new_n14520_, new_n14521_,
    new_n14522_, new_n14523_, new_n14524_, new_n14525_, new_n14526_,
    new_n14527_, new_n14528_, new_n14529_, new_n14530_, new_n14531_,
    new_n14532_, new_n14533_, new_n14534_, new_n14535_, new_n14536_,
    new_n14537_, new_n14538_, new_n14539_, new_n14540_, new_n14541_,
    new_n14542_, new_n14543_, new_n14544_, new_n14545_, new_n14546_,
    new_n14547_, new_n14548_, new_n14549_, new_n14550_, new_n14551_,
    new_n14552_, new_n14553_, new_n14554_, new_n14555_, new_n14556_,
    new_n14557_, new_n14558_, new_n14559_, new_n14560_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14581_,
    new_n14582_, new_n14583_, new_n14584_, new_n14585_, new_n14586_,
    new_n14587_, new_n14588_, new_n14589_, new_n14590_, new_n14591_,
    new_n14592_, new_n14593_, new_n14594_, new_n14595_, new_n14596_,
    new_n14597_, new_n14598_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14639_, new_n14640_, new_n14641_,
    new_n14642_, new_n14643_, new_n14644_, new_n14645_, new_n14646_,
    new_n14647_, new_n14648_, new_n14649_, new_n14650_, new_n14651_,
    new_n14652_, new_n14653_, new_n14654_, new_n14655_, new_n14656_,
    new_n14657_, new_n14658_, new_n14659_, new_n14660_, new_n14661_,
    new_n14662_, new_n14663_, new_n14664_, new_n14665_, new_n14666_,
    new_n14667_, new_n14668_, new_n14669_, new_n14670_, new_n14671_,
    new_n14672_, new_n14673_, new_n14674_, new_n14675_, new_n14676_,
    new_n14677_, new_n14678_, new_n14679_, new_n14680_, new_n14681_,
    new_n14682_, new_n14683_, new_n14684_, new_n14685_, new_n14686_,
    new_n14687_, new_n14688_, new_n14689_, new_n14690_, new_n14691_,
    new_n14692_, new_n14693_, new_n14694_, new_n14695_, new_n14696_,
    new_n14697_, new_n14698_, new_n14699_, new_n14700_, new_n14701_,
    new_n14702_, new_n14703_, new_n14704_, new_n14705_, new_n14706_,
    new_n14707_, new_n14708_, new_n14709_, new_n14710_, new_n14711_,
    new_n14712_, new_n14713_, new_n14714_, new_n14715_, new_n14716_,
    new_n14717_, new_n14718_, new_n14719_, new_n14720_, new_n14721_,
    new_n14722_, new_n14723_, new_n14724_, new_n14725_, new_n14726_,
    new_n14727_, new_n14728_, new_n14729_, new_n14730_, new_n14731_,
    new_n14732_, new_n14733_, new_n14734_, new_n14735_, new_n14736_,
    new_n14737_, new_n14738_, new_n14739_, new_n14740_, new_n14741_,
    new_n14742_, new_n14743_, new_n14744_, new_n14745_, new_n14746_,
    new_n14747_, new_n14748_, new_n14749_, new_n14750_, new_n14751_,
    new_n14752_, new_n14753_, new_n14754_, new_n14755_, new_n14756_,
    new_n14757_, new_n14758_, new_n14759_, new_n14760_, new_n14761_,
    new_n14762_, new_n14763_, new_n14764_, new_n14765_, new_n14766_,
    new_n14767_, new_n14768_, new_n14769_, new_n14770_, new_n14771_,
    new_n14772_, new_n14773_, new_n14774_, new_n14775_, new_n14776_,
    new_n14777_, new_n14778_, new_n14779_, new_n14780_, new_n14781_,
    new_n14782_, new_n14783_, new_n14784_, new_n14785_, new_n14786_,
    new_n14787_, new_n14788_, new_n14789_, new_n14790_, new_n14791_,
    new_n14792_, new_n14793_, new_n14794_, new_n14795_, new_n14796_,
    new_n14797_, new_n14798_, new_n14799_, new_n14800_, new_n14801_,
    new_n14802_, new_n14803_, new_n14804_, new_n14805_, new_n14806_,
    new_n14807_, new_n14808_, new_n14809_, new_n14810_, new_n14811_,
    new_n14812_, new_n14813_, new_n14814_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14958_, new_n14959_, new_n14960_, new_n14961_,
    new_n14962_, new_n14963_, new_n14964_, new_n14965_, new_n14966_,
    new_n14967_, new_n14968_, new_n14969_, new_n14970_, new_n14971_,
    new_n14972_, new_n14973_, new_n14974_, new_n14975_, new_n14976_,
    new_n14977_, new_n14978_, new_n14979_, new_n14980_, new_n14981_,
    new_n14982_, new_n14983_, new_n14984_, new_n14985_, new_n14986_,
    new_n14987_, new_n14988_, new_n14989_, new_n14990_, new_n14991_,
    new_n14992_, new_n14993_, new_n14994_, new_n14995_, new_n14996_,
    new_n14997_, new_n14998_, new_n14999_, new_n15000_, new_n15001_,
    new_n15002_, new_n15003_, new_n15004_, new_n15005_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15036_,
    new_n15037_, new_n15038_, new_n15039_, new_n15040_, new_n15041_,
    new_n15042_, new_n15043_, new_n15044_, new_n15045_, new_n15046_,
    new_n15047_, new_n15048_, new_n15049_, new_n15050_, new_n15051_,
    new_n15052_, new_n15053_, new_n15054_, new_n15055_, new_n15056_,
    new_n15057_, new_n15058_, new_n15059_, new_n15060_, new_n15061_,
    new_n15062_, new_n15063_, new_n15064_, new_n15065_, new_n15066_,
    new_n15067_, new_n15068_, new_n15069_, new_n15070_, new_n15071_,
    new_n15072_, new_n15073_, new_n15074_, new_n15075_, new_n15076_,
    new_n15077_, new_n15078_, new_n15079_, new_n15080_, new_n15081_,
    new_n15082_, new_n15083_, new_n15084_, new_n15085_, new_n15086_,
    new_n15087_, new_n15088_, new_n15089_, new_n15090_, new_n15091_,
    new_n15092_, new_n15093_, new_n15094_, new_n15095_, new_n15096_,
    new_n15097_, new_n15098_, new_n15099_, new_n15100_, new_n15101_,
    new_n15102_, new_n15103_, new_n15104_, new_n15105_, new_n15106_,
    new_n15107_, new_n15108_, new_n15109_, new_n15110_, new_n15111_,
    new_n15112_, new_n15113_, new_n15114_, new_n15115_, new_n15116_,
    new_n15117_, new_n15118_, new_n15119_, new_n15120_, new_n15121_,
    new_n15122_, new_n15123_, new_n15124_, new_n15125_, new_n15126_,
    new_n15127_, new_n15128_, new_n15129_, new_n15130_, new_n15131_,
    new_n15132_, new_n15133_, new_n15134_, new_n15135_, new_n15136_,
    new_n15137_, new_n15138_, new_n15139_, new_n15140_, new_n15141_,
    new_n15142_, new_n15143_, new_n15144_, new_n15145_, new_n15146_,
    new_n15147_, new_n15148_, new_n15149_, new_n15150_, new_n15151_,
    new_n15152_, new_n15153_, new_n15154_, new_n15155_, new_n15156_,
    new_n15157_, new_n15158_, new_n15159_, new_n15160_, new_n15161_,
    new_n15162_, new_n15163_, new_n15164_, new_n15165_, new_n15166_,
    new_n15167_, new_n15168_, new_n15169_, new_n15170_, new_n15171_,
    new_n15172_, new_n15173_, new_n15174_, new_n15175_, new_n15176_,
    new_n15177_, new_n15178_, new_n15179_, new_n15180_, new_n15181_,
    new_n15182_, new_n15183_, new_n15184_, new_n15185_, new_n15186_,
    new_n15187_, new_n15188_, new_n15189_, new_n15190_, new_n15191_,
    new_n15192_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15215_, new_n15216_,
    new_n15217_, new_n15218_, new_n15219_, new_n15220_, new_n15221_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15228_, new_n15229_, new_n15230_, new_n15231_,
    new_n15232_, new_n15233_, new_n15234_, new_n15235_, new_n15236_,
    new_n15237_, new_n15238_, new_n15239_, new_n15240_, new_n15241_,
    new_n15242_, new_n15243_, new_n15244_, new_n15245_, new_n15246_,
    new_n15247_, new_n15248_, new_n15249_, new_n15250_, new_n15251_,
    new_n15252_, new_n15253_, new_n15254_, new_n15255_, new_n15256_,
    new_n15257_, new_n15258_, new_n15259_, new_n15260_, new_n15261_,
    new_n15262_, new_n15263_, new_n15264_, new_n15265_, new_n15266_,
    new_n15267_, new_n15268_, new_n15269_, new_n15270_, new_n15271_,
    new_n15272_, new_n15273_, new_n15274_, new_n15275_, new_n15276_,
    new_n15277_, new_n15278_, new_n15279_, new_n15280_, new_n15281_,
    new_n15282_, new_n15283_, new_n15284_, new_n15285_, new_n15286_,
    new_n15287_, new_n15288_, new_n15289_, new_n15290_, new_n15291_,
    new_n15292_, new_n15293_, new_n15294_, new_n15295_, new_n15296_,
    new_n15297_, new_n15298_, new_n15299_, new_n15300_, new_n15301_,
    new_n15302_, new_n15303_, new_n15304_, new_n15305_, new_n15306_,
    new_n15307_, new_n15308_, new_n15309_, new_n15310_, new_n15311_,
    new_n15312_, new_n15313_, new_n15314_, new_n15315_, new_n15316_,
    new_n15317_, new_n15318_, new_n15319_, new_n15320_, new_n15321_,
    new_n15322_, new_n15323_, new_n15324_, new_n15325_, new_n15326_,
    new_n15327_, new_n15328_, new_n15329_, new_n15330_, new_n15331_,
    new_n15332_, new_n15333_, new_n15334_, new_n15335_, new_n15336_,
    new_n15337_, new_n15338_, new_n15339_, new_n15340_, new_n15341_,
    new_n15342_, new_n15343_, new_n15344_, new_n15345_, new_n15346_,
    new_n15347_, new_n15348_, new_n15349_, new_n15350_, new_n15351_,
    new_n15352_, new_n15353_, new_n15354_, new_n15355_, new_n15356_,
    new_n15357_, new_n15358_, new_n15359_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15410_, new_n15411_,
    new_n15412_, new_n15413_, new_n15414_, new_n15415_, new_n15416_,
    new_n15417_, new_n15418_, new_n15419_, new_n15420_, new_n15421_,
    new_n15422_, new_n15423_, new_n15424_, new_n15425_, new_n15426_,
    new_n15427_, new_n15428_, new_n15429_, new_n15430_, new_n15431_,
    new_n15432_, new_n15433_, new_n15434_, new_n15435_, new_n15436_,
    new_n15437_, new_n15438_, new_n15439_, new_n15440_, new_n15441_,
    new_n15442_, new_n15443_, new_n15444_, new_n15445_, new_n15446_,
    new_n15447_, new_n15448_, new_n15449_, new_n15450_, new_n15451_,
    new_n15452_, new_n15453_, new_n15454_, new_n15455_, new_n15456_,
    new_n15457_, new_n15458_, new_n15459_, new_n15460_, new_n15461_,
    new_n15462_, new_n15463_, new_n15464_, new_n15465_, new_n15466_,
    new_n15467_, new_n15468_, new_n15469_, new_n15470_, new_n15471_,
    new_n15472_, new_n15473_, new_n15474_, new_n15475_, new_n15476_,
    new_n15477_, new_n15478_, new_n15479_, new_n15480_, new_n15481_,
    new_n15482_, new_n15483_, new_n15484_, new_n15485_, new_n15486_,
    new_n15487_, new_n15488_, new_n15489_, new_n15490_, new_n15491_,
    new_n15492_, new_n15493_, new_n15494_, new_n15495_, new_n15496_,
    new_n15497_, new_n15498_, new_n15499_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15540_, new_n15541_, new_n15542_, new_n15543_,
    new_n15544_, new_n15545_, new_n15546_, new_n15547_, new_n15548_,
    new_n15549_, new_n15550_, new_n15551_, new_n15552_, new_n15553_,
    new_n15554_, new_n15555_, new_n15556_, new_n15557_, new_n15558_,
    new_n15559_, new_n15560_, new_n15561_, new_n15562_, new_n15563_,
    new_n15564_, new_n15565_, new_n15566_, new_n15567_, new_n15568_,
    new_n15569_, new_n15570_, new_n15571_, new_n15572_, new_n15573_,
    new_n15574_, new_n15575_, new_n15576_, new_n15577_, new_n15578_,
    new_n15579_, new_n15580_, new_n15581_, new_n15582_, new_n15583_,
    new_n15584_, new_n15585_, new_n15586_, new_n15587_, new_n15588_,
    new_n15589_, new_n15590_, new_n15591_, new_n15592_, new_n15593_,
    new_n15594_, new_n15595_, new_n15596_, new_n15597_, new_n15598_,
    new_n15599_, new_n15600_, new_n15601_, new_n15602_, new_n15603_,
    new_n15604_, new_n15605_, new_n15606_, new_n15607_, new_n15608_,
    new_n15609_, new_n15610_, new_n15611_, new_n15612_, new_n15613_,
    new_n15614_, new_n15615_, new_n15616_, new_n15617_, new_n15618_,
    new_n15619_, new_n15620_, new_n15621_, new_n15622_, new_n15623_,
    new_n15624_, new_n15625_, new_n15626_, new_n15627_, new_n15628_,
    new_n15629_, new_n15630_, new_n15631_, new_n15632_, new_n15633_,
    new_n15634_, new_n15635_, new_n15636_, new_n15637_, new_n15638_,
    new_n15639_, new_n15640_, new_n15641_, new_n15642_, new_n15643_,
    new_n15644_, new_n15645_, new_n15646_, new_n15647_, new_n15648_,
    new_n15649_, new_n15650_, new_n15651_, new_n15652_, new_n15653_,
    new_n15654_, new_n15655_, new_n15656_, new_n15657_, new_n15658_,
    new_n15659_, new_n15660_, new_n15661_, new_n15662_, new_n15663_,
    new_n15664_, new_n15665_, new_n15666_, new_n15667_, new_n15668_,
    new_n15669_, new_n15670_, new_n15671_, new_n15672_, new_n15673_,
    new_n15674_, new_n15675_, new_n15676_, new_n15677_, new_n15678_,
    new_n15679_, new_n15680_, new_n15681_, new_n15682_, new_n15683_,
    new_n15684_, new_n15685_, new_n15686_, new_n15687_, new_n15688_,
    new_n15689_, new_n15690_, new_n15691_, new_n15692_, new_n15693_,
    new_n15694_, new_n15695_, new_n15696_, new_n15697_, new_n15698_,
    new_n15699_, new_n15700_, new_n15701_, new_n15702_, new_n15703_,
    new_n15704_, new_n15705_, new_n15706_, new_n15707_, new_n15708_,
    new_n15709_, new_n15710_, new_n15711_, new_n15712_, new_n15713_,
    new_n15714_, new_n15715_, new_n15716_, new_n15717_, new_n15718_,
    new_n15719_, new_n15720_, new_n15721_, new_n15722_, new_n15723_,
    new_n15724_, new_n15725_, new_n15726_, new_n15727_, new_n15728_,
    new_n15729_, new_n15730_, new_n15731_, new_n15732_, new_n15733_,
    new_n15734_, new_n15735_, new_n15736_, new_n15737_, new_n15738_,
    new_n15739_, new_n15740_, new_n15741_, new_n15742_, new_n15743_,
    new_n15744_, new_n15745_, new_n15746_, new_n15747_, new_n15748_,
    new_n15749_, new_n15750_, new_n15751_, new_n15752_, new_n15753_,
    new_n15754_, new_n15755_, new_n15756_, new_n15757_, new_n15758_,
    new_n15759_, new_n15760_, new_n15761_, new_n15762_, new_n15763_,
    new_n15764_, new_n15765_, new_n15766_, new_n15767_, new_n15768_,
    new_n15769_, new_n15770_, new_n15771_, new_n15772_, new_n15773_,
    new_n15774_, new_n15775_, new_n15776_, new_n15777_, new_n15778_,
    new_n15779_, new_n15780_, new_n15781_, new_n15782_, new_n15783_,
    new_n15784_, new_n15785_, new_n15786_, new_n15787_, new_n15788_,
    new_n15789_, new_n15790_, new_n15791_, new_n15792_, new_n15793_,
    new_n15794_, new_n15795_, new_n15796_, new_n15797_, new_n15798_,
    new_n15799_, new_n15800_, new_n15801_, new_n15802_, new_n15803_,
    new_n15804_, new_n15805_, new_n15806_, new_n15807_, new_n15808_,
    new_n15809_, new_n15810_, new_n15811_, new_n15812_, new_n15813_,
    new_n15814_, new_n15815_, new_n15816_, new_n15817_, new_n15818_,
    new_n15819_, new_n15820_, new_n15821_, new_n15822_, new_n15823_,
    new_n15824_, new_n15825_, new_n15826_, new_n15827_, new_n15828_,
    new_n15829_, new_n15830_, new_n15831_, new_n15832_, new_n15833_,
    new_n15834_, new_n15835_, new_n15836_, new_n15837_, new_n15838_,
    new_n15839_, new_n15840_, new_n15841_, new_n15842_, new_n15843_,
    new_n15844_, new_n15845_, new_n15846_, new_n15847_, new_n15848_,
    new_n15849_, new_n15850_, new_n15851_, new_n15852_, new_n15853_,
    new_n15854_, new_n15855_, new_n15856_, new_n15857_, new_n15858_,
    new_n15859_, new_n15860_, new_n15861_, new_n15862_, new_n15863_,
    new_n15864_, new_n15865_, new_n15866_, new_n15867_, new_n15868_,
    new_n15869_, new_n15870_, new_n15871_, new_n15872_, new_n15873_,
    new_n15874_, new_n15875_, new_n15876_, new_n15877_, new_n15878_,
    new_n15879_, new_n15880_, new_n15881_, new_n15882_, new_n15883_,
    new_n15884_, new_n15885_, new_n15886_, new_n15887_, new_n15888_,
    new_n15889_, new_n15890_, new_n15891_, new_n15892_, new_n15893_,
    new_n15894_, new_n15895_, new_n15896_, new_n15897_, new_n15898_,
    new_n15899_, new_n15900_, new_n15901_, new_n15902_, new_n15903_,
    new_n15904_, new_n15905_, new_n15906_, new_n15907_, new_n15908_,
    new_n15909_, new_n15910_, new_n15911_, new_n15912_, new_n15913_,
    new_n15914_, new_n15915_, new_n15916_, new_n15917_, new_n15918_,
    new_n15919_, new_n15920_, new_n15921_, new_n15922_, new_n15923_,
    new_n15924_, new_n15925_, new_n15926_, new_n15927_, new_n15928_,
    new_n15929_, new_n15930_, new_n15931_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15939_, new_n15940_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15947_, new_n15948_,
    new_n15949_, new_n15950_, new_n15951_, new_n15952_, new_n15953_,
    new_n15954_, new_n15955_, new_n15956_, new_n15957_, new_n15958_,
    new_n15959_, new_n15960_, new_n15961_, new_n15962_, new_n15963_,
    new_n15964_, new_n15965_, new_n15966_, new_n15967_, new_n15968_,
    new_n15969_, new_n15970_, new_n15971_, new_n15972_, new_n15973_,
    new_n15974_, new_n15975_, new_n15976_, new_n15977_, new_n15978_,
    new_n15979_, new_n15980_, new_n15981_, new_n15982_, new_n15983_,
    new_n15984_, new_n15985_, new_n15986_, new_n15987_, new_n15988_,
    new_n15989_, new_n15990_, new_n15991_, new_n15992_, new_n15993_,
    new_n15994_, new_n15995_, new_n15996_, new_n15997_, new_n15998_,
    new_n15999_, new_n16000_, new_n16001_, new_n16002_, new_n16003_,
    new_n16004_, new_n16005_, new_n16006_, new_n16007_, new_n16008_,
    new_n16009_, new_n16010_, new_n16011_, new_n16012_, new_n16013_,
    new_n16014_, new_n16015_, new_n16016_, new_n16017_, new_n16018_,
    new_n16019_, new_n16020_, new_n16021_, new_n16022_, new_n16023_,
    new_n16024_, new_n16025_, new_n16026_, new_n16027_, new_n16028_,
    new_n16029_, new_n16030_, new_n16031_, new_n16032_, new_n16033_,
    new_n16034_, new_n16035_, new_n16036_, new_n16037_, new_n16038_,
    new_n16039_, new_n16040_, new_n16041_, new_n16042_, new_n16043_,
    new_n16044_, new_n16045_, new_n16046_, new_n16047_, new_n16048_,
    new_n16049_, new_n16050_, new_n16051_, new_n16052_, new_n16053_,
    new_n16054_, new_n16055_, new_n16056_, new_n16057_, new_n16058_,
    new_n16059_, new_n16060_, new_n16061_, new_n16062_, new_n16063_,
    new_n16064_, new_n16065_, new_n16066_, new_n16067_, new_n16068_,
    new_n16069_, new_n16070_, new_n16071_, new_n16072_, new_n16073_,
    new_n16074_, new_n16075_, new_n16076_, new_n16077_, new_n16078_,
    new_n16079_, new_n16080_, new_n16081_, new_n16082_, new_n16083_,
    new_n16084_, new_n16085_, new_n16086_, new_n16087_, new_n16088_,
    new_n16089_, new_n16090_, new_n16091_, new_n16092_, new_n16093_,
    new_n16094_, new_n16095_, new_n16096_, new_n16097_, new_n16098_,
    new_n16099_, new_n16100_, new_n16101_, new_n16102_, new_n16103_,
    new_n16104_, new_n16105_, new_n16106_, new_n16107_, new_n16108_,
    new_n16109_, new_n16110_, new_n16111_, new_n16112_, new_n16113_,
    new_n16114_, new_n16115_, new_n16116_, new_n16117_, new_n16118_,
    new_n16119_, new_n16120_, new_n16121_, new_n16122_, new_n16123_,
    new_n16124_, new_n16125_, new_n16126_, new_n16127_, new_n16128_,
    new_n16129_, new_n16130_, new_n16131_, new_n16132_, new_n16133_,
    new_n16134_, new_n16135_, new_n16136_, new_n16137_, new_n16138_,
    new_n16139_, new_n16140_, new_n16141_, new_n16142_, new_n16143_,
    new_n16144_, new_n16145_, new_n16146_, new_n16147_, new_n16148_,
    new_n16149_, new_n16150_, new_n16151_, new_n16152_, new_n16153_,
    new_n16154_, new_n16155_, new_n16156_, new_n16157_, new_n16158_,
    new_n16159_, new_n16160_, new_n16161_, new_n16162_, new_n16163_,
    new_n16164_, new_n16165_, new_n16166_, new_n16167_, new_n16168_,
    new_n16169_, new_n16170_, new_n16171_, new_n16172_, new_n16173_,
    new_n16174_, new_n16175_, new_n16176_, new_n16177_, new_n16178_,
    new_n16179_, new_n16180_, new_n16181_, new_n16182_, new_n16183_,
    new_n16184_, new_n16185_, new_n16186_, new_n16187_, new_n16188_,
    new_n16189_, new_n16190_, new_n16191_, new_n16192_, new_n16193_,
    new_n16194_, new_n16195_, new_n16196_, new_n16197_, new_n16198_,
    new_n16199_, new_n16200_, new_n16201_, new_n16202_, new_n16203_,
    new_n16204_, new_n16205_, new_n16206_, new_n16207_, new_n16208_,
    new_n16209_, new_n16210_, new_n16211_, new_n16212_, new_n16213_,
    new_n16214_, new_n16215_, new_n16216_, new_n16217_, new_n16218_,
    new_n16219_, new_n16220_, new_n16221_, new_n16222_, new_n16223_,
    new_n16224_, new_n16225_, new_n16226_, new_n16227_, new_n16228_,
    new_n16229_, new_n16230_, new_n16231_, new_n16232_, new_n16233_,
    new_n16234_, new_n16235_, new_n16236_, new_n16237_, new_n16238_,
    new_n16239_, new_n16240_, new_n16241_, new_n16242_, new_n16243_,
    new_n16244_, new_n16245_, new_n16246_, new_n16247_, new_n16248_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16255_, new_n16256_, new_n16257_, new_n16258_,
    new_n16259_, new_n16260_, new_n16261_, new_n16262_, new_n16263_,
    new_n16264_, new_n16265_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16270_, new_n16271_, new_n16272_, new_n16273_,
    new_n16274_, new_n16275_, new_n16276_, new_n16277_, new_n16278_,
    new_n16279_, new_n16280_, new_n16281_, new_n16282_, new_n16283_,
    new_n16284_, new_n16285_, new_n16286_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16291_, new_n16292_, new_n16293_,
    new_n16294_, new_n16295_, new_n16296_, new_n16297_, new_n16298_,
    new_n16299_, new_n16300_, new_n16301_, new_n16302_, new_n16303_,
    new_n16304_, new_n16305_, new_n16306_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16313_,
    new_n16314_, new_n16315_, new_n16316_, new_n16317_, new_n16318_,
    new_n16319_, new_n16320_, new_n16321_, new_n16322_, new_n16323_,
    new_n16324_, new_n16325_, new_n16326_, new_n16327_, new_n16328_,
    new_n16329_, new_n16330_, new_n16331_, new_n16332_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16346_, new_n16347_, new_n16348_,
    new_n16349_, new_n16350_, new_n16351_, new_n16352_, new_n16353_,
    new_n16354_, new_n16355_, new_n16356_, new_n16357_, new_n16358_,
    new_n16359_, new_n16360_, new_n16361_, new_n16362_, new_n16363_,
    new_n16364_, new_n16365_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16463_,
    new_n16464_, new_n16465_, new_n16466_, new_n16467_, new_n16468_,
    new_n16469_, new_n16470_, new_n16471_, new_n16472_, new_n16473_,
    new_n16474_, new_n16475_, new_n16476_, new_n16477_, new_n16478_,
    new_n16479_, new_n16480_, new_n16481_, new_n16482_, new_n16483_,
    new_n16484_, new_n16485_, new_n16486_, new_n16487_, new_n16488_,
    new_n16489_, new_n16490_, new_n16491_, new_n16492_, new_n16493_,
    new_n16494_, new_n16495_, new_n16496_, new_n16497_, new_n16498_,
    new_n16499_, new_n16500_, new_n16501_, new_n16502_, new_n16503_,
    new_n16504_, new_n16505_, new_n16506_, new_n16507_, new_n16508_,
    new_n16509_, new_n16510_, new_n16511_, new_n16512_, new_n16513_,
    new_n16514_, new_n16515_, new_n16516_, new_n16517_, new_n16518_,
    new_n16519_, new_n16520_, new_n16521_, new_n16522_, new_n16523_,
    new_n16524_, new_n16525_, new_n16526_, new_n16527_, new_n16528_,
    new_n16529_, new_n16530_, new_n16531_, new_n16532_, new_n16533_,
    new_n16534_, new_n16535_, new_n16536_, new_n16537_, new_n16538_,
    new_n16539_, new_n16540_, new_n16541_, new_n16542_, new_n16543_,
    new_n16544_, new_n16545_, new_n16546_, new_n16547_, new_n16548_,
    new_n16549_, new_n16550_, new_n16551_, new_n16552_, new_n16553_,
    new_n16554_, new_n16555_, new_n16556_, new_n16557_, new_n16558_,
    new_n16559_, new_n16560_, new_n16561_, new_n16562_, new_n16563_,
    new_n16564_, new_n16565_, new_n16566_, new_n16567_, new_n16568_,
    new_n16569_, new_n16570_, new_n16571_, new_n16572_, new_n16573_,
    new_n16574_, new_n16575_, new_n16576_, new_n16577_, new_n16578_,
    new_n16579_, new_n16580_, new_n16581_, new_n16582_, new_n16583_,
    new_n16584_, new_n16585_, new_n16586_, new_n16587_, new_n16588_,
    new_n16589_, new_n16590_, new_n16591_, new_n16592_, new_n16593_,
    new_n16594_, new_n16595_, new_n16596_, new_n16597_, new_n16598_,
    new_n16599_, new_n16600_, new_n16601_, new_n16602_, new_n16603_,
    new_n16604_, new_n16605_, new_n16606_, new_n16607_, new_n16608_,
    new_n16609_, new_n16610_, new_n16611_, new_n16612_, new_n16613_,
    new_n16614_, new_n16615_, new_n16616_, new_n16617_, new_n16618_,
    new_n16619_, new_n16620_, new_n16621_, new_n16622_, new_n16623_,
    new_n16624_, new_n16625_, new_n16626_, new_n16627_, new_n16628_,
    new_n16629_, new_n16630_, new_n16631_, new_n16632_, new_n16633_,
    new_n16634_, new_n16635_, new_n16636_, new_n16637_, new_n16638_,
    new_n16639_, new_n16640_, new_n16641_, new_n16642_, new_n16643_,
    new_n16644_, new_n16645_, new_n16646_, new_n16647_, new_n16648_,
    new_n16649_, new_n16650_, new_n16651_, new_n16652_, new_n16653_,
    new_n16654_, new_n16655_, new_n16656_, new_n16657_, new_n16658_,
    new_n16659_, new_n16660_, new_n16661_, new_n16662_, new_n16663_,
    new_n16664_, new_n16665_, new_n16666_, new_n16667_, new_n16668_,
    new_n16669_, new_n16670_, new_n16671_, new_n16672_, new_n16673_,
    new_n16674_, new_n16675_, new_n16676_, new_n16677_, new_n16678_,
    new_n16679_, new_n16680_, new_n16681_, new_n16682_, new_n16683_,
    new_n16684_, new_n16685_, new_n16686_, new_n16687_, new_n16688_,
    new_n16689_, new_n16690_, new_n16691_, new_n16692_, new_n16693_,
    new_n16694_, new_n16695_, new_n16696_, new_n16697_, new_n16698_,
    new_n16699_, new_n16700_, new_n16701_, new_n16702_, new_n16703_,
    new_n16704_, new_n16705_, new_n16706_, new_n16707_, new_n16708_,
    new_n16709_, new_n16710_, new_n16711_, new_n16712_, new_n16713_,
    new_n16714_, new_n16715_, new_n16716_, new_n16717_, new_n16718_,
    new_n16719_, new_n16720_, new_n16721_, new_n16722_, new_n16723_,
    new_n16724_, new_n16725_, new_n16726_, new_n16727_, new_n16728_,
    new_n16729_, new_n16730_, new_n16731_, new_n16732_, new_n16733_,
    new_n16734_, new_n16735_, new_n16736_, new_n16737_, new_n16738_,
    new_n16739_, new_n16740_, new_n16741_, new_n16742_, new_n16743_,
    new_n16744_, new_n16745_, new_n16746_, new_n16747_, new_n16748_,
    new_n16749_, new_n16750_, new_n16751_, new_n16752_, new_n16753_,
    new_n16754_, new_n16755_, new_n16756_, new_n16757_, new_n16758_,
    new_n16759_, new_n16760_, new_n16761_, new_n16762_, new_n16763_,
    new_n16764_, new_n16765_, new_n16766_, new_n16767_, new_n16768_,
    new_n16769_, new_n16770_, new_n16771_, new_n16772_, new_n16773_,
    new_n16774_, new_n16775_, new_n16776_, new_n16777_, new_n16778_,
    new_n16779_, new_n16780_, new_n16781_, new_n16782_, new_n16783_,
    new_n16784_, new_n16785_, new_n16786_, new_n16787_, new_n16788_,
    new_n16789_, new_n16790_, new_n16791_, new_n16792_, new_n16793_,
    new_n16794_, new_n16795_, new_n16796_, new_n16797_, new_n16798_,
    new_n16799_, new_n16800_, new_n16801_, new_n16802_, new_n16803_,
    new_n16804_, new_n16805_, new_n16806_, new_n16807_, new_n16808_,
    new_n16809_, new_n16810_, new_n16811_, new_n16812_, new_n16813_,
    new_n16814_, new_n16815_, new_n16816_, new_n16817_, new_n16818_,
    new_n16819_, new_n16820_, new_n16821_, new_n16822_, new_n16823_,
    new_n16824_, new_n16825_, new_n16826_, new_n16827_, new_n16828_,
    new_n16829_, new_n16830_, new_n16831_, new_n16832_, new_n16833_,
    new_n16834_, new_n16835_, new_n16836_, new_n16837_, new_n16838_,
    new_n16839_, new_n16840_, new_n16841_, new_n16842_, new_n16843_,
    new_n16844_, new_n16845_, new_n16846_, new_n16847_, new_n16848_,
    new_n16849_, new_n16850_, new_n16851_, new_n16852_, new_n16853_,
    new_n16854_, new_n16855_, new_n16856_, new_n16857_, new_n16858_,
    new_n16859_, new_n16860_, new_n16861_, new_n16862_, new_n16863_,
    new_n16864_, new_n16865_, new_n16866_, new_n16867_, new_n16868_,
    new_n16869_, new_n16870_, new_n16871_, new_n16872_, new_n16873_,
    new_n16874_, new_n16875_, new_n16876_, new_n16877_, new_n16878_,
    new_n16879_, new_n16880_, new_n16881_, new_n16882_, new_n16883_,
    new_n16884_, new_n16885_, new_n16886_, new_n16887_, new_n16888_,
    new_n16889_, new_n16890_, new_n16891_, new_n16892_, new_n16893_,
    new_n16894_, new_n16895_, new_n16896_, new_n16897_, new_n16898_,
    new_n16899_, new_n16900_, new_n16901_, new_n16902_, new_n16903_,
    new_n16904_, new_n16905_, new_n16906_, new_n16907_, new_n16908_,
    new_n16909_, new_n16910_, new_n16911_, new_n16912_, new_n16913_,
    new_n16914_, new_n16915_, new_n16916_, new_n16917_, new_n16918_,
    new_n16919_, new_n16920_, new_n16921_, new_n16922_, new_n16923_,
    new_n16924_, new_n16925_, new_n16926_, new_n16927_, new_n16928_,
    new_n16929_, new_n16930_, new_n16931_, new_n16932_, new_n16933_,
    new_n16934_, new_n16935_, new_n16936_, new_n16937_, new_n16938_,
    new_n16939_, new_n16940_, new_n16941_, new_n16942_, new_n16943_,
    new_n16944_, new_n16945_, new_n16946_, new_n16947_, new_n16948_,
    new_n16949_, new_n16950_, new_n16951_, new_n16952_, new_n16953_,
    new_n16954_, new_n16955_, new_n16956_, new_n16957_, new_n16958_,
    new_n16959_, new_n16960_, new_n16961_, new_n16962_, new_n16963_,
    new_n16964_, new_n16965_, new_n16966_, new_n16967_, new_n16968_,
    new_n16969_, new_n16970_, new_n16971_, new_n16972_, new_n16973_,
    new_n16974_, new_n16975_, new_n16976_, new_n16977_, new_n16978_,
    new_n16979_, new_n16980_, new_n16981_, new_n16982_, new_n16983_,
    new_n16984_, new_n16985_, new_n16986_, new_n16987_, new_n16988_,
    new_n16989_, new_n16990_, new_n16991_, new_n16992_, new_n16993_,
    new_n16994_, new_n16995_, new_n16996_, new_n16997_, new_n16998_,
    new_n16999_, new_n17000_, new_n17001_, new_n17002_, new_n17003_,
    new_n17004_, new_n17005_, new_n17006_, new_n17007_, new_n17008_,
    new_n17009_, new_n17010_, new_n17011_, new_n17012_, new_n17013_,
    new_n17015_, new_n17016_, new_n17017_, new_n17018_, new_n17019_,
    new_n17020_, new_n17021_, new_n17022_, new_n17023_, new_n17024_,
    new_n17025_, new_n17026_, new_n17027_, new_n17028_, new_n17029_,
    new_n17030_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17041_, new_n17042_, new_n17043_, new_n17044_, new_n17045_,
    new_n17046_, new_n17047_, new_n17048_, new_n17049_, new_n17050_,
    new_n17051_, new_n17052_, new_n17053_, new_n17054_, new_n17055_,
    new_n17056_, new_n17057_, new_n17058_, new_n17059_, new_n17060_,
    new_n17061_, new_n17062_, new_n17063_, new_n17064_, new_n17065_,
    new_n17066_, new_n17067_, new_n17068_, new_n17069_, new_n17070_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17106_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17125_, new_n17126_, new_n17127_, new_n17128_,
    new_n17129_, new_n17130_, new_n17131_, new_n17132_, new_n17133_,
    new_n17135_, new_n17136_, new_n17137_, new_n17138_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17283_, new_n17284_, new_n17285_, new_n17286_,
    new_n17287_, new_n17288_, new_n17289_, new_n17290_, new_n17291_,
    new_n17292_, new_n17293_, new_n17294_, new_n17295_, new_n17296_,
    new_n17297_, new_n17298_, new_n17299_, new_n17300_, new_n17301_,
    new_n17302_, new_n17303_, new_n17304_, new_n17305_, new_n17306_,
    new_n17307_, new_n17308_, new_n17309_, new_n17310_, new_n17311_,
    new_n17312_, new_n17313_, new_n17314_, new_n17315_, new_n17316_,
    new_n17317_, new_n17318_, new_n17319_, new_n17320_, new_n17321_,
    new_n17322_, new_n17323_, new_n17324_, new_n17325_, new_n17326_,
    new_n17327_, new_n17328_, new_n17329_, new_n17330_, new_n17331_,
    new_n17332_, new_n17333_, new_n17334_, new_n17335_, new_n17336_,
    new_n17337_, new_n17338_, new_n17339_, new_n17340_, new_n17341_,
    new_n17342_, new_n17343_, new_n17344_, new_n17345_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17398_, new_n17399_, new_n17400_, new_n17401_,
    new_n17402_, new_n17403_, new_n17404_, new_n17405_, new_n17406_,
    new_n17407_, new_n17408_, new_n17409_, new_n17410_, new_n17411_,
    new_n17412_, new_n17413_, new_n17414_, new_n17415_, new_n17416_,
    new_n17417_, new_n17418_, new_n17419_, new_n17420_, new_n17421_,
    new_n17422_, new_n17423_, new_n17424_, new_n17425_, new_n17426_,
    new_n17427_, new_n17428_, new_n17429_, new_n17430_, new_n17431_,
    new_n17432_, new_n17433_, new_n17434_, new_n17435_, new_n17436_,
    new_n17437_, new_n17438_, new_n17439_, new_n17440_, new_n17441_,
    new_n17442_, new_n17443_, new_n17444_, new_n17445_, new_n17446_,
    new_n17447_, new_n17448_, new_n17449_, new_n17450_, new_n17451_,
    new_n17452_, new_n17453_, new_n17454_, new_n17455_, new_n17456_,
    new_n17457_, new_n17458_, new_n17459_, new_n17460_, new_n17461_,
    new_n17462_, new_n17463_, new_n17464_, new_n17465_, new_n17466_,
    new_n17467_, new_n17468_, new_n17469_, new_n17470_, new_n17471_,
    new_n17472_, new_n17473_, new_n17474_, new_n17475_, new_n17476_,
    new_n17477_, new_n17478_, new_n17479_, new_n17480_, new_n17481_,
    new_n17482_, new_n17483_, new_n17484_, new_n17485_, new_n17486_,
    new_n17487_, new_n17488_, new_n17489_, new_n17490_, new_n17491_,
    new_n17492_, new_n17493_, new_n17494_, new_n17495_, new_n17496_,
    new_n17497_, new_n17498_, new_n17499_, new_n17500_, new_n17501_,
    new_n17502_, new_n17503_, new_n17504_, new_n17505_, new_n17506_,
    new_n17507_, new_n17508_, new_n17509_, new_n17510_, new_n17511_,
    new_n17512_, new_n17513_, new_n17514_, new_n17515_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17560_, new_n17561_, new_n17562_,
    new_n17563_, new_n17564_, new_n17565_, new_n17566_, new_n17567_,
    new_n17568_, new_n17569_, new_n17570_, new_n17571_, new_n17572_,
    new_n17573_, new_n17574_, new_n17575_, new_n17576_, new_n17577_,
    new_n17578_, new_n17579_, new_n17580_, new_n17581_, new_n17582_,
    new_n17583_, new_n17584_, new_n17585_, new_n17586_, new_n17587_,
    new_n17588_, new_n17589_, new_n17590_, new_n17591_, new_n17592_,
    new_n17593_, new_n17594_, new_n17595_, new_n17596_, new_n17597_,
    new_n17598_, new_n17599_, new_n17600_, new_n17601_, new_n17602_,
    new_n17603_, new_n17604_, new_n17605_, new_n17606_, new_n17607_,
    new_n17608_, new_n17609_, new_n17610_, new_n17611_, new_n17612_,
    new_n17613_, new_n17614_, new_n17615_, new_n17616_, new_n17617_,
    new_n17618_, new_n17619_, new_n17620_, new_n17621_, new_n17622_,
    new_n17623_, new_n17624_, new_n17625_, new_n17626_, new_n17627_,
    new_n17628_, new_n17629_, new_n17630_, new_n17631_, new_n17632_,
    new_n17633_, new_n17634_, new_n17635_, new_n17636_, new_n17637_,
    new_n17638_, new_n17639_, new_n17640_, new_n17641_, new_n17642_,
    new_n17643_, new_n17644_, new_n17645_, new_n17646_, new_n17647_,
    new_n17648_, new_n17649_, new_n17650_, new_n17651_, new_n17652_,
    new_n17653_, new_n17654_, new_n17655_, new_n17656_, new_n17657_,
    new_n17658_, new_n17659_, new_n17660_, new_n17661_, new_n17662_,
    new_n17663_, new_n17664_, new_n17665_, new_n17666_, new_n17667_,
    new_n17668_, new_n17669_, new_n17670_, new_n17671_, new_n17672_,
    new_n17673_, new_n17674_, new_n17675_, new_n17676_, new_n17677_,
    new_n17678_, new_n17679_, new_n17680_, new_n17681_, new_n17682_,
    new_n17683_, new_n17684_, new_n17685_, new_n17686_, new_n17687_,
    new_n17688_, new_n17689_, new_n17690_, new_n17691_, new_n17692_,
    new_n17693_, new_n17694_, new_n17695_, new_n17696_, new_n17697_,
    new_n17698_, new_n17699_, new_n17700_, new_n17701_, new_n17702_,
    new_n17703_, new_n17704_, new_n17705_, new_n17706_, new_n17707_,
    new_n17708_, new_n17709_, new_n17710_, new_n17711_, new_n17712_,
    new_n17713_, new_n17714_, new_n17715_, new_n17716_, new_n17717_,
    new_n17718_, new_n17719_, new_n17720_, new_n17721_, new_n17722_,
    new_n17723_, new_n17724_, new_n17725_, new_n17726_, new_n17727_,
    new_n17728_, new_n17729_, new_n17730_, new_n17731_, new_n17732_,
    new_n17733_, new_n17734_, new_n17735_, new_n17736_, new_n17737_,
    new_n17738_, new_n17739_, new_n17740_, new_n17741_, new_n17742_,
    new_n17743_, new_n17744_, new_n17745_, new_n17746_, new_n17747_,
    new_n17748_, new_n17749_, new_n17750_, new_n17751_, new_n17752_,
    new_n17753_, new_n17754_, new_n17755_, new_n17756_, new_n17757_,
    new_n17758_, new_n17759_, new_n17760_, new_n17761_, new_n17762_,
    new_n17763_, new_n17764_, new_n17765_, new_n17766_, new_n17767_,
    new_n17768_, new_n17769_, new_n17770_, new_n17771_, new_n17772_,
    new_n17773_, new_n17774_, new_n17775_, new_n17776_, new_n17777_,
    new_n17778_, new_n17779_, new_n17780_, new_n17781_, new_n17782_,
    new_n17783_, new_n17784_, new_n17785_, new_n17786_, new_n17787_,
    new_n17788_, new_n17789_, new_n17790_, new_n17791_, new_n17792_,
    new_n17793_, new_n17794_, new_n17795_, new_n17796_, new_n17797_,
    new_n17798_, new_n17799_, new_n17800_, new_n17801_, new_n17802_,
    new_n17803_, new_n17804_, new_n17805_, new_n17806_, new_n17807_,
    new_n17808_, new_n17809_, new_n17810_, new_n17811_, new_n17812_,
    new_n17813_, new_n17814_, new_n17815_, new_n17816_, new_n17817_,
    new_n17818_, new_n17819_, new_n17820_, new_n17821_, new_n17822_,
    new_n17823_, new_n17824_, new_n17825_, new_n17826_, new_n17827_,
    new_n17828_, new_n17829_, new_n17830_, new_n17831_, new_n17832_,
    new_n17833_, new_n17834_, new_n17835_, new_n17836_, new_n17837_,
    new_n17838_, new_n17839_, new_n17840_, new_n17841_, new_n17842_,
    new_n17843_, new_n17844_, new_n17845_, new_n17846_, new_n17847_,
    new_n17848_, new_n17849_, new_n17850_, new_n17851_, new_n17852_,
    new_n17853_, new_n17854_, new_n17855_, new_n17856_, new_n17857_,
    new_n17858_, new_n17859_, new_n17860_, new_n17861_, new_n17862_,
    new_n17863_, new_n17864_, new_n17865_, new_n17866_, new_n17867_,
    new_n17868_, new_n17869_, new_n17870_, new_n17871_, new_n17872_,
    new_n17873_, new_n17874_, new_n17875_, new_n17876_, new_n17877_,
    new_n17878_, new_n17879_, new_n17880_, new_n17881_, new_n17882_,
    new_n17883_, new_n17884_, new_n17885_, new_n17886_, new_n17887_,
    new_n17888_, new_n17889_, new_n17890_, new_n17891_, new_n17892_,
    new_n17893_, new_n17894_, new_n17895_, new_n17896_, new_n17897_,
    new_n17898_, new_n17899_, new_n17900_, new_n17901_, new_n17902_,
    new_n17903_, new_n17904_, new_n17905_, new_n17906_, new_n17907_,
    new_n17908_, new_n17909_, new_n17910_, new_n17911_, new_n17912_,
    new_n17913_, new_n17914_, new_n17915_, new_n17916_, new_n17917_,
    new_n17918_, new_n17919_, new_n17920_, new_n17921_, new_n17922_,
    new_n17923_, new_n17924_, new_n17925_, new_n17926_, new_n17927_,
    new_n17928_, new_n17929_, new_n17930_, new_n17931_, new_n17932_,
    new_n17933_, new_n17934_, new_n17935_, new_n17936_, new_n17937_,
    new_n17938_, new_n17939_, new_n17940_, new_n17941_, new_n17942_,
    new_n17943_, new_n17944_, new_n17945_, new_n17946_, new_n17947_,
    new_n17948_, new_n17949_, new_n17950_, new_n17951_, new_n17952_,
    new_n17953_, new_n17954_, new_n17955_, new_n17956_, new_n17957_,
    new_n17958_, new_n17959_, new_n17960_, new_n17961_, new_n17962_,
    new_n17963_, new_n17964_, new_n17965_, new_n17966_, new_n17967_,
    new_n17968_, new_n17969_, new_n17970_, new_n17971_, new_n17972_,
    new_n17973_, new_n17974_, new_n17975_, new_n17976_, new_n17977_,
    new_n17978_, new_n17979_, new_n17980_, new_n17981_, new_n17982_,
    new_n17983_, new_n17984_, new_n17985_, new_n17986_, new_n17987_,
    new_n17988_, new_n17989_, new_n17990_, new_n17991_, new_n17992_,
    new_n17993_, new_n17994_, new_n17995_, new_n17996_, new_n17997_,
    new_n17998_, new_n17999_, new_n18000_, new_n18001_, new_n18002_,
    new_n18003_, new_n18004_, new_n18005_, new_n18006_, new_n18007_,
    new_n18008_, new_n18009_, new_n18010_, new_n18011_, new_n18012_,
    new_n18013_, new_n18014_, new_n18015_, new_n18016_, new_n18017_,
    new_n18018_, new_n18019_, new_n18020_, new_n18021_, new_n18022_,
    new_n18023_, new_n18024_, new_n18025_, new_n18026_, new_n18027_,
    new_n18028_, new_n18029_, new_n18030_, new_n18031_, new_n18032_,
    new_n18033_, new_n18034_, new_n18035_, new_n18036_, new_n18037_,
    new_n18038_, new_n18039_, new_n18040_, new_n18041_, new_n18042_,
    new_n18043_, new_n18044_, new_n18045_, new_n18046_, new_n18047_,
    new_n18048_, new_n18049_, new_n18050_, new_n18051_, new_n18052_,
    new_n18053_, new_n18054_, new_n18055_, new_n18056_, new_n18057_,
    new_n18058_, new_n18059_, new_n18060_, new_n18061_, new_n18062_,
    new_n18063_, new_n18064_, new_n18065_, new_n18066_, new_n18067_,
    new_n18068_, new_n18069_, new_n18070_, new_n18071_, new_n18072_,
    new_n18073_, new_n18074_, new_n18075_, new_n18076_, new_n18077_,
    new_n18078_, new_n18079_, new_n18080_, new_n18081_, new_n18082_,
    new_n18083_, new_n18084_, new_n18085_, new_n18086_, new_n18087_,
    new_n18088_, new_n18089_, new_n18090_, new_n18091_, new_n18092_,
    new_n18093_, new_n18094_, new_n18095_, new_n18096_, new_n18097_,
    new_n18098_, new_n18099_, new_n18100_, new_n18101_, new_n18102_,
    new_n18103_, new_n18104_, new_n18105_, new_n18106_, new_n18107_,
    new_n18108_, new_n18109_, new_n18110_, new_n18111_, new_n18112_,
    new_n18113_, new_n18114_, new_n18115_, new_n18116_, new_n18117_,
    new_n18118_, new_n18119_, new_n18120_, new_n18121_, new_n18123_,
    new_n18124_, new_n18125_, new_n18126_, new_n18127_, new_n18128_,
    new_n18129_, new_n18130_, new_n18131_, new_n18132_, new_n18133_,
    new_n18134_, new_n18135_, new_n18136_, new_n18137_, new_n18138_,
    new_n18139_, new_n18140_, new_n18141_, new_n18142_, new_n18143_,
    new_n18144_, new_n18145_, new_n18146_, new_n18147_, new_n18148_,
    new_n18149_, new_n18150_, new_n18151_, new_n18152_, new_n18153_,
    new_n18154_, new_n18155_, new_n18156_, new_n18157_, new_n18158_,
    new_n18159_, new_n18160_, new_n18161_, new_n18162_, new_n18163_,
    new_n18164_, new_n18165_, new_n18166_, new_n18167_, new_n18168_,
    new_n18169_, new_n18170_, new_n18171_, new_n18172_, new_n18173_,
    new_n18174_, new_n18175_, new_n18176_, new_n18177_, new_n18178_,
    new_n18179_, new_n18180_, new_n18181_, new_n18182_, new_n18183_,
    new_n18184_, new_n18185_, new_n18186_, new_n18187_, new_n18188_,
    new_n18189_, new_n18190_, new_n18191_, new_n18192_, new_n18193_,
    new_n18194_, new_n18195_, new_n18196_, new_n18197_, new_n18198_,
    new_n18199_, new_n18200_, new_n18201_, new_n18202_, new_n18203_,
    new_n18204_, new_n18205_, new_n18206_, new_n18207_, new_n18208_,
    new_n18209_, new_n18210_, new_n18211_, new_n18212_, new_n18213_,
    new_n18214_, new_n18215_, new_n18216_, new_n18217_, new_n18218_,
    new_n18219_, new_n18220_, new_n18221_, new_n18222_, new_n18223_,
    new_n18224_, new_n18225_, new_n18226_, new_n18227_, new_n18228_,
    new_n18229_, new_n18230_, new_n18231_, new_n18232_, new_n18233_,
    new_n18234_, new_n18235_, new_n18236_, new_n18237_, new_n18238_,
    new_n18239_, new_n18240_, new_n18241_, new_n18242_, new_n18243_,
    new_n18244_, new_n18245_, new_n18246_, new_n18247_, new_n18248_,
    new_n18249_, new_n18250_, new_n18251_, new_n18252_, new_n18253_,
    new_n18254_, new_n18255_, new_n18256_, new_n18257_, new_n18258_,
    new_n18259_, new_n18260_, new_n18261_, new_n18262_, new_n18263_,
    new_n18264_, new_n18265_, new_n18266_, new_n18267_, new_n18268_,
    new_n18269_, new_n18270_, new_n18271_, new_n18272_, new_n18273_,
    new_n18274_, new_n18275_, new_n18276_, new_n18277_, new_n18278_,
    new_n18279_, new_n18280_, new_n18281_, new_n18282_, new_n18283_,
    new_n18284_, new_n18285_, new_n18286_, new_n18287_, new_n18288_,
    new_n18289_, new_n18290_, new_n18291_, new_n18292_, new_n18293_,
    new_n18294_, new_n18295_, new_n18296_, new_n18297_, new_n18298_,
    new_n18299_, new_n18300_, new_n18301_, new_n18302_, new_n18303_,
    new_n18304_, new_n18305_, new_n18306_, new_n18307_, new_n18308_,
    new_n18309_, new_n18310_, new_n18311_, new_n18312_, new_n18313_,
    new_n18314_, new_n18315_, new_n18316_, new_n18317_, new_n18318_,
    new_n18319_, new_n18320_, new_n18321_, new_n18322_, new_n18323_,
    new_n18324_, new_n18325_, new_n18326_, new_n18327_, new_n18328_,
    new_n18329_, new_n18330_, new_n18331_, new_n18332_, new_n18333_,
    new_n18334_, new_n18335_, new_n18336_, new_n18337_, new_n18338_,
    new_n18339_, new_n18340_, new_n18341_, new_n18342_, new_n18343_,
    new_n18344_, new_n18345_, new_n18346_, new_n18347_, new_n18348_,
    new_n18349_, new_n18350_, new_n18351_, new_n18352_, new_n18353_,
    new_n18354_, new_n18355_, new_n18356_, new_n18357_, new_n18358_,
    new_n18359_, new_n18360_, new_n18361_, new_n18362_, new_n18363_,
    new_n18364_, new_n18365_, new_n18366_, new_n18367_, new_n18368_,
    new_n18369_, new_n18370_, new_n18371_, new_n18372_, new_n18373_,
    new_n18374_, new_n18375_, new_n18376_, new_n18377_, new_n18378_,
    new_n18379_, new_n18380_, new_n18381_, new_n18382_, new_n18383_,
    new_n18384_, new_n18385_, new_n18386_, new_n18387_, new_n18388_,
    new_n18389_, new_n18390_, new_n18391_, new_n18392_, new_n18393_,
    new_n18394_, new_n18395_, new_n18396_, new_n18397_, new_n18398_,
    new_n18399_, new_n18400_, new_n18401_, new_n18402_, new_n18403_,
    new_n18404_, new_n18405_, new_n18406_, new_n18407_, new_n18408_,
    new_n18409_, new_n18410_, new_n18411_, new_n18412_, new_n18413_,
    new_n18414_, new_n18415_, new_n18416_, new_n18417_, new_n18418_,
    new_n18419_, new_n18420_, new_n18421_, new_n18422_, new_n18423_,
    new_n18424_, new_n18425_, new_n18426_, new_n18427_, new_n18428_,
    new_n18429_, new_n18430_, new_n18431_, new_n18432_, new_n18433_,
    new_n18434_, new_n18435_, new_n18436_, new_n18437_, new_n18438_,
    new_n18439_, new_n18440_, new_n18441_, new_n18442_, new_n18443_,
    new_n18444_, new_n18445_, new_n18446_, new_n18447_, new_n18448_,
    new_n18449_, new_n18450_, new_n18451_, new_n18452_, new_n18453_,
    new_n18454_, new_n18455_, new_n18456_, new_n18457_, new_n18458_,
    new_n18459_, new_n18460_, new_n18461_, new_n18462_, new_n18463_,
    new_n18464_, new_n18465_, new_n18466_, new_n18467_, new_n18468_,
    new_n18469_, new_n18470_, new_n18471_, new_n18472_, new_n18473_,
    new_n18474_, new_n18475_, new_n18476_, new_n18477_, new_n18478_,
    new_n18479_, new_n18480_, new_n18481_, new_n18482_, new_n18483_,
    new_n18484_, new_n18485_, new_n18486_, new_n18487_, new_n18488_,
    new_n18489_, new_n18490_, new_n18491_, new_n18492_, new_n18493_,
    new_n18494_, new_n18495_, new_n18496_, new_n18497_, new_n18498_,
    new_n18499_, new_n18500_, new_n18501_, new_n18502_, new_n18503_,
    new_n18504_, new_n18505_, new_n18506_, new_n18507_, new_n18508_,
    new_n18509_, new_n18510_, new_n18511_, new_n18512_, new_n18513_,
    new_n18514_, new_n18515_, new_n18516_, new_n18517_, new_n18518_,
    new_n18519_, new_n18520_, new_n18521_, new_n18522_, new_n18523_,
    new_n18524_, new_n18525_, new_n18526_, new_n18527_, new_n18528_,
    new_n18529_, new_n18530_, new_n18531_, new_n18532_, new_n18533_,
    new_n18534_, new_n18535_, new_n18536_, new_n18537_, new_n18538_,
    new_n18539_, new_n18540_, new_n18541_, new_n18542_, new_n18543_,
    new_n18544_, new_n18545_, new_n18546_, new_n18547_, new_n18548_,
    new_n18549_, new_n18550_, new_n18551_, new_n18552_, new_n18553_,
    new_n18554_, new_n18555_, new_n18556_, new_n18557_, new_n18558_,
    new_n18559_, new_n18560_, new_n18561_, new_n18562_, new_n18563_,
    new_n18564_, new_n18565_, new_n18566_, new_n18567_, new_n18568_,
    new_n18569_, new_n18570_, new_n18571_, new_n18572_, new_n18573_,
    new_n18574_, new_n18575_, new_n18576_, new_n18577_, new_n18578_,
    new_n18579_, new_n18580_, new_n18581_, new_n18582_, new_n18583_,
    new_n18584_, new_n18585_, new_n18586_, new_n18587_, new_n18588_,
    new_n18589_, new_n18590_, new_n18591_, new_n18592_, new_n18593_,
    new_n18594_, new_n18595_, new_n18596_, new_n18597_, new_n18598_,
    new_n18599_, new_n18600_, new_n18601_, new_n18602_, new_n18603_,
    new_n18604_, new_n18605_, new_n18606_, new_n18607_, new_n18608_,
    new_n18609_, new_n18610_, new_n18611_, new_n18612_, new_n18613_,
    new_n18614_, new_n18615_, new_n18616_, new_n18617_, new_n18618_,
    new_n18619_, new_n18620_, new_n18621_, new_n18622_, new_n18623_,
    new_n18624_, new_n18625_, new_n18626_, new_n18627_, new_n18628_,
    new_n18629_, new_n18630_, new_n18631_, new_n18632_, new_n18633_,
    new_n18634_, new_n18635_, new_n18636_, new_n18637_, new_n18638_,
    new_n18639_, new_n18640_, new_n18641_, new_n18642_, new_n18643_,
    new_n18644_, new_n18645_, new_n18646_, new_n18647_, new_n18648_,
    new_n18649_, new_n18650_, new_n18651_, new_n18652_, new_n18653_,
    new_n18654_, new_n18655_, new_n18656_, new_n18657_, new_n18658_,
    new_n18659_, new_n18660_, new_n18661_, new_n18662_, new_n18663_,
    new_n18664_, new_n18665_, new_n18666_, new_n18667_, new_n18668_,
    new_n18669_, new_n18670_, new_n18671_, new_n18672_, new_n18673_,
    new_n18674_, new_n18675_, new_n18676_, new_n18677_, new_n18678_,
    new_n18679_, new_n18680_, new_n18681_, new_n18682_, new_n18683_,
    new_n18684_, new_n18685_, new_n18686_, new_n18687_, new_n18688_,
    new_n18689_, new_n18690_, new_n18691_, new_n18692_, new_n18693_,
    new_n18694_, new_n18695_, new_n18696_, new_n18697_, new_n18698_,
    new_n18699_, new_n18700_, new_n18701_, new_n18702_, new_n18703_,
    new_n18704_, new_n18705_, new_n18706_, new_n18707_, new_n18708_,
    new_n18709_, new_n18710_, new_n18711_, new_n18712_, new_n18713_,
    new_n18714_, new_n18715_, new_n18716_, new_n18717_, new_n18718_,
    new_n18719_, new_n18720_, new_n18721_, new_n18722_, new_n18723_,
    new_n18724_, new_n18725_, new_n18726_, new_n18727_, new_n18728_,
    new_n18729_, new_n18730_, new_n18731_, new_n18732_, new_n18733_,
    new_n18734_, new_n18735_, new_n18736_, new_n18737_, new_n18738_,
    new_n18739_, new_n18740_, new_n18741_, new_n18742_, new_n18743_,
    new_n18744_, new_n18745_, new_n18746_, new_n18747_, new_n18748_,
    new_n18749_, new_n18750_, new_n18751_, new_n18752_, new_n18753_,
    new_n18754_, new_n18755_, new_n18756_, new_n18757_, new_n18758_,
    new_n18759_, new_n18760_, new_n18761_, new_n18762_, new_n18763_,
    new_n18764_, new_n18765_, new_n18766_, new_n18767_, new_n18768_,
    new_n18769_, new_n18770_, new_n18771_, new_n18772_, new_n18773_,
    new_n18774_, new_n18775_, new_n18776_, new_n18777_, new_n18778_,
    new_n18779_, new_n18780_, new_n18782_, new_n18783_, new_n18784_,
    new_n18785_, new_n18786_, new_n18787_, new_n18788_, new_n18789_,
    new_n18790_, new_n18791_, new_n18792_, new_n18793_, new_n18794_,
    new_n18795_, new_n18796_, new_n18797_, new_n18798_, new_n18799_,
    new_n18800_, new_n18801_, new_n18802_, new_n18803_, new_n18804_,
    new_n18805_, new_n18806_, new_n18807_, new_n18808_, new_n18809_,
    new_n18810_, new_n18811_, new_n18812_, new_n18813_, new_n18814_,
    new_n18815_, new_n18816_, new_n18817_, new_n18818_, new_n18819_,
    new_n18820_, new_n18821_, new_n18822_, new_n18823_, new_n18824_,
    new_n18825_, new_n18826_, new_n18827_, new_n18828_, new_n18829_,
    new_n18830_, new_n18831_, new_n18832_, new_n18833_, new_n18834_,
    new_n18835_, new_n18836_, new_n18837_, new_n18838_, new_n18839_,
    new_n18840_, new_n18841_, new_n18842_, new_n18843_, new_n18844_,
    new_n18845_, new_n18846_, new_n18847_, new_n18848_, new_n18849_,
    new_n18850_, new_n18851_, new_n18852_, new_n18853_, new_n18854_,
    new_n18855_, new_n18856_, new_n18857_, new_n18858_, new_n18859_,
    new_n18860_, new_n18861_, new_n18862_, new_n18863_, new_n18864_,
    new_n18865_, new_n18866_, new_n18867_, new_n18868_, new_n18869_,
    new_n18870_, new_n18871_, new_n18872_, new_n18873_, new_n18874_,
    new_n18875_, new_n18876_, new_n18877_, new_n18878_, new_n18879_,
    new_n18880_, new_n18881_, new_n18882_, new_n18883_, new_n18884_,
    new_n18885_, new_n18886_, new_n18887_, new_n18888_, new_n18889_,
    new_n18890_, new_n18891_, new_n18892_, new_n18893_, new_n18894_,
    new_n18895_, new_n18896_, new_n18897_, new_n18898_, new_n18899_,
    new_n18900_, new_n18901_, new_n18902_, new_n18903_, new_n18904_,
    new_n18905_, new_n18906_, new_n18907_, new_n18908_, new_n18909_,
    new_n18910_, new_n18911_, new_n18912_, new_n18913_, new_n18914_,
    new_n18915_, new_n18916_, new_n18917_, new_n18918_, new_n18919_,
    new_n18920_, new_n18921_, new_n18922_, new_n18923_, new_n18924_,
    new_n18925_, new_n18926_, new_n18927_, new_n18928_, new_n18929_,
    new_n18930_, new_n18931_, new_n18932_, new_n18933_, new_n18934_,
    new_n18935_, new_n18936_, new_n18937_, new_n18938_, new_n18939_,
    new_n18940_, new_n18941_, new_n18942_, new_n18943_, new_n18944_,
    new_n18945_, new_n18946_, new_n18947_, new_n18948_, new_n18949_,
    new_n18950_, new_n18951_, new_n18952_, new_n18953_, new_n18954_,
    new_n18955_, new_n18956_, new_n18957_, new_n18958_, new_n18959_,
    new_n18960_, new_n18961_, new_n18962_, new_n18963_, new_n18964_,
    new_n18965_, new_n18966_, new_n18967_, new_n18968_, new_n18969_,
    new_n18970_, new_n18971_, new_n18972_, new_n18973_, new_n18974_,
    new_n18975_, new_n18976_, new_n18977_, new_n18978_, new_n18979_,
    new_n18980_, new_n18981_, new_n18982_, new_n18983_, new_n18984_,
    new_n18985_, new_n18986_, new_n18987_, new_n18988_, new_n18989_,
    new_n18990_, new_n18991_, new_n18992_, new_n18993_, new_n18994_,
    new_n18995_, new_n18996_, new_n18997_, new_n18998_, new_n18999_,
    new_n19000_, new_n19001_, new_n19002_, new_n19003_, new_n19004_,
    new_n19005_, new_n19006_, new_n19007_, new_n19008_, new_n19009_,
    new_n19010_, new_n19011_, new_n19012_, new_n19013_, new_n19014_,
    new_n19015_, new_n19016_, new_n19017_, new_n19018_, new_n19019_,
    new_n19020_, new_n19021_, new_n19022_, new_n19023_, new_n19024_,
    new_n19025_, new_n19026_, new_n19027_, new_n19028_, new_n19029_,
    new_n19030_, new_n19031_, new_n19032_, new_n19033_, new_n19034_,
    new_n19035_, new_n19036_, new_n19037_, new_n19038_, new_n19039_,
    new_n19040_, new_n19041_, new_n19042_, new_n19043_, new_n19044_,
    new_n19045_, new_n19046_, new_n19047_, new_n19048_, new_n19049_,
    new_n19050_, new_n19051_, new_n19052_, new_n19053_, new_n19054_,
    new_n19055_, new_n19056_, new_n19057_, new_n19058_, new_n19059_,
    new_n19060_, new_n19061_, new_n19062_, new_n19063_, new_n19064_,
    new_n19065_, new_n19066_, new_n19067_, new_n19068_, new_n19069_,
    new_n19070_, new_n19071_, new_n19072_, new_n19073_, new_n19074_,
    new_n19075_, new_n19076_, new_n19077_, new_n19078_, new_n19079_,
    new_n19080_, new_n19081_, new_n19082_, new_n19083_, new_n19084_,
    new_n19085_, new_n19086_, new_n19087_, new_n19088_, new_n19089_,
    new_n19090_, new_n19091_, new_n19092_, new_n19093_, new_n19094_,
    new_n19095_, new_n19096_, new_n19097_, new_n19098_, new_n19099_,
    new_n19100_, new_n19101_, new_n19102_, new_n19103_, new_n19104_,
    new_n19105_, new_n19106_, new_n19107_, new_n19108_, new_n19109_,
    new_n19110_, new_n19111_, new_n19112_, new_n19113_, new_n19114_,
    new_n19115_, new_n19116_, new_n19117_, new_n19118_, new_n19119_,
    new_n19120_, new_n19121_, new_n19122_, new_n19123_, new_n19124_,
    new_n19125_, new_n19126_, new_n19127_, new_n19128_, new_n19129_,
    new_n19130_, new_n19131_, new_n19132_, new_n19133_, new_n19134_,
    new_n19135_, new_n19136_, new_n19137_, new_n19138_, new_n19139_,
    new_n19140_, new_n19141_, new_n19142_, new_n19143_, new_n19144_,
    new_n19145_, new_n19146_, new_n19147_, new_n19148_, new_n19149_,
    new_n19150_, new_n19151_, new_n19152_, new_n19153_, new_n19154_,
    new_n19155_, new_n19156_, new_n19157_, new_n19158_, new_n19159_,
    new_n19160_, new_n19161_, new_n19162_, new_n19163_, new_n19164_,
    new_n19165_, new_n19166_, new_n19167_, new_n19168_, new_n19169_,
    new_n19170_, new_n19171_, new_n19172_, new_n19173_, new_n19174_,
    new_n19175_, new_n19176_, new_n19177_, new_n19178_, new_n19179_,
    new_n19180_, new_n19181_, new_n19182_, new_n19183_, new_n19184_,
    new_n19185_, new_n19186_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19456_, new_n19457_, new_n19458_, new_n19459_,
    new_n19460_, new_n19461_, new_n19462_, new_n19463_, new_n19464_,
    new_n19465_, new_n19466_, new_n19467_, new_n19468_, new_n19469_,
    new_n19470_, new_n19471_, new_n19472_, new_n19473_, new_n19474_,
    new_n19475_, new_n19476_, new_n19477_, new_n19478_, new_n19479_,
    new_n19480_, new_n19481_, new_n19482_, new_n19483_, new_n19484_,
    new_n19485_, new_n19486_, new_n19487_, new_n19488_, new_n19489_,
    new_n19490_, new_n19491_, new_n19492_, new_n19493_, new_n19494_,
    new_n19495_, new_n19496_, new_n19497_, new_n19498_, new_n19499_,
    new_n19500_, new_n19501_, new_n19502_, new_n19503_, new_n19504_,
    new_n19505_, new_n19506_, new_n19507_, new_n19508_, new_n19509_,
    new_n19510_, new_n19511_, new_n19512_, new_n19513_, new_n19514_,
    new_n19515_, new_n19516_, new_n19517_, new_n19518_, new_n19519_,
    new_n19520_, new_n19521_, new_n19522_, new_n19523_, new_n19524_,
    new_n19525_, new_n19526_, new_n19527_, new_n19528_, new_n19529_,
    new_n19530_, new_n19531_, new_n19532_, new_n19533_, new_n19534_,
    new_n19535_, new_n19536_, new_n19537_, new_n19538_, new_n19539_,
    new_n19540_, new_n19541_, new_n19542_, new_n19543_, new_n19544_,
    new_n19545_, new_n19546_, new_n19547_, new_n19548_, new_n19549_,
    new_n19550_, new_n19551_, new_n19552_, new_n19553_, new_n19554_,
    new_n19555_, new_n19556_, new_n19557_, new_n19558_, new_n19559_,
    new_n19560_, new_n19561_, new_n19562_, new_n19563_, new_n19564_,
    new_n19565_, new_n19566_, new_n19567_, new_n19568_, new_n19569_,
    new_n19570_, new_n19571_, new_n19572_, new_n19573_, new_n19574_,
    new_n19575_, new_n19576_, new_n19577_, new_n19578_, new_n19579_,
    new_n19580_, new_n19581_, new_n19582_, new_n19583_, new_n19584_,
    new_n19585_, new_n19586_, new_n19587_, new_n19588_, new_n19589_,
    new_n19590_, new_n19591_, new_n19592_, new_n19593_, new_n19594_,
    new_n19595_, new_n19596_, new_n19597_, new_n19598_, new_n19599_,
    new_n19600_, new_n19601_, new_n19602_, new_n19603_, new_n19604_,
    new_n19605_, new_n19606_, new_n19607_, new_n19608_, new_n19609_,
    new_n19610_, new_n19611_, new_n19612_, new_n19613_, new_n19614_,
    new_n19615_, new_n19616_, new_n19617_, new_n19618_, new_n19619_,
    new_n19620_, new_n19621_, new_n19622_, new_n19623_, new_n19624_,
    new_n19625_, new_n19626_, new_n19627_, new_n19628_, new_n19629_,
    new_n19630_, new_n19631_, new_n19632_, new_n19633_, new_n19634_,
    new_n19635_, new_n19636_, new_n19637_, new_n19638_, new_n19639_,
    new_n19640_, new_n19641_, new_n19642_, new_n19643_, new_n19644_,
    new_n19645_, new_n19646_, new_n19647_, new_n19648_, new_n19649_,
    new_n19650_, new_n19651_, new_n19652_, new_n19653_, new_n19654_,
    new_n19655_, new_n19656_, new_n19657_, new_n19658_, new_n19659_,
    new_n19660_, new_n19661_, new_n19662_, new_n19663_, new_n19664_,
    new_n19665_, new_n19666_, new_n19667_, new_n19668_, new_n19669_,
    new_n19670_, new_n19671_, new_n19672_, new_n19673_, new_n19674_,
    new_n19675_, new_n19676_, new_n19677_, new_n19678_, new_n19679_,
    new_n19680_, new_n19681_, new_n19682_, new_n19683_, new_n19684_,
    new_n19685_, new_n19686_, new_n19687_, new_n19688_, new_n19689_,
    new_n19690_, new_n19691_, new_n19692_, new_n19693_, new_n19694_,
    new_n19695_, new_n19696_, new_n19697_, new_n19698_, new_n19699_,
    new_n19700_, new_n19701_, new_n19702_, new_n19703_, new_n19704_,
    new_n19705_, new_n19706_, new_n19707_, new_n19708_, new_n19709_,
    new_n19710_, new_n19711_, new_n19712_, new_n19713_, new_n19714_,
    new_n19715_, new_n19716_, new_n19717_, new_n19718_, new_n19719_,
    new_n19720_, new_n19721_, new_n19722_, new_n19723_, new_n19724_,
    new_n19725_, new_n19726_, new_n19727_, new_n19728_, new_n19729_,
    new_n19730_, new_n19731_, new_n19732_, new_n19733_, new_n19734_,
    new_n19735_, new_n19736_, new_n19737_, new_n19738_, new_n19739_,
    new_n19740_, new_n19741_, new_n19742_, new_n19743_, new_n19744_,
    new_n19745_, new_n19746_, new_n19747_, new_n19748_, new_n19749_,
    new_n19750_, new_n19751_, new_n19752_, new_n19753_, new_n19754_,
    new_n19755_, new_n19756_, new_n19757_, new_n19758_, new_n19759_,
    new_n19760_, new_n19761_, new_n19762_, new_n19763_, new_n19764_,
    new_n19765_, new_n19766_, new_n19767_, new_n19768_, new_n19769_,
    new_n19770_, new_n19771_, new_n19772_, new_n19773_, new_n19774_,
    new_n19775_, new_n19776_, new_n19777_, new_n19778_, new_n19779_,
    new_n19780_, new_n19781_, new_n19782_, new_n19783_, new_n19784_,
    new_n19785_, new_n19786_, new_n19787_, new_n19788_, new_n19789_,
    new_n19790_, new_n19791_, new_n19792_, new_n19793_, new_n19794_,
    new_n19795_, new_n19796_, new_n19797_, new_n19798_, new_n19799_,
    new_n19800_, new_n19801_, new_n19802_, new_n19803_, new_n19804_,
    new_n19805_, new_n19806_, new_n19807_, new_n19808_, new_n19809_,
    new_n19810_, new_n19811_, new_n19812_, new_n19813_, new_n19814_,
    new_n19815_, new_n19816_, new_n19817_, new_n19818_, new_n19819_,
    new_n19820_, new_n19821_, new_n19822_, new_n19823_, new_n19824_,
    new_n19825_, new_n19826_, new_n19827_, new_n19828_, new_n19829_,
    new_n19830_, new_n19831_, new_n19832_, new_n19833_, new_n19834_,
    new_n19835_, new_n19836_, new_n19837_, new_n19838_, new_n19839_,
    new_n19840_, new_n19841_, new_n19842_, new_n19843_, new_n19844_,
    new_n19845_, new_n19846_, new_n19847_, new_n19848_, new_n19849_,
    new_n19850_, new_n19851_, new_n19852_, new_n19853_, new_n19854_,
    new_n19855_, new_n19856_, new_n19857_, new_n19858_, new_n19859_,
    new_n19860_, new_n19861_, new_n19862_, new_n19863_, new_n19864_,
    new_n19865_, new_n19866_, new_n19867_, new_n19868_, new_n19869_,
    new_n19870_, new_n19871_, new_n19872_, new_n19873_, new_n19874_,
    new_n19875_, new_n19876_, new_n19877_, new_n19878_, new_n19879_,
    new_n19880_, new_n19881_, new_n19882_, new_n19883_, new_n19884_,
    new_n19885_, new_n19886_, new_n19887_, new_n19888_, new_n19889_,
    new_n19890_, new_n19891_, new_n19892_, new_n19893_, new_n19894_,
    new_n19895_, new_n19896_, new_n19897_, new_n19898_, new_n19899_,
    new_n19901_, new_n19902_, new_n19903_, new_n19904_, new_n19905_,
    new_n19906_, new_n19907_, new_n19908_, new_n19909_, new_n19910_,
    new_n19911_, new_n19912_, new_n19913_, new_n19914_, new_n19915_,
    new_n19916_, new_n19917_, new_n19918_, new_n19919_, new_n19920_,
    new_n19921_, new_n19922_, new_n19923_, new_n19924_, new_n19925_,
    new_n19926_, new_n19927_, new_n19928_, new_n19929_, new_n19930_,
    new_n19931_, new_n19932_, new_n19933_, new_n19934_, new_n19935_,
    new_n19936_, new_n19937_, new_n19938_, new_n19939_, new_n19940_,
    new_n19941_, new_n19942_, new_n19943_, new_n19944_, new_n19945_,
    new_n19946_, new_n19947_, new_n19948_, new_n19949_, new_n19950_,
    new_n19951_, new_n19952_, new_n19953_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19991_, new_n19992_,
    new_n19993_, new_n19994_, new_n19995_, new_n19996_, new_n19997_,
    new_n19998_, new_n19999_, new_n20000_, new_n20001_, new_n20002_,
    new_n20003_, new_n20004_, new_n20005_, new_n20006_, new_n20007_,
    new_n20008_, new_n20009_, new_n20011_, new_n20012_, new_n20013_,
    new_n20014_, new_n20015_, new_n20016_, new_n20017_, new_n20018_,
    new_n20019_, new_n20021_, new_n20022_, new_n20023_, new_n20024_,
    new_n20027_, new_n20028_, new_n20029_, new_n20030_, new_n20031_,
    new_n20032_, new_n20033_, new_n20034_, new_n20035_, new_n20036_,
    new_n20037_, new_n20038_, new_n20039_, new_n20040_, new_n20041_,
    new_n20042_, new_n20043_, new_n20044_, new_n20045_, new_n20046_,
    new_n20047_, new_n20048_, new_n20049_, new_n20050_, new_n20051_,
    new_n20052_, new_n20053_, new_n20054_, new_n20055_, new_n20056_,
    new_n20057_, new_n20058_, new_n20059_, new_n20060_, new_n20061_,
    new_n20062_, new_n20063_, new_n20064_, new_n20065_, new_n20066_,
    new_n20067_, new_n20068_, new_n20069_, new_n20070_, new_n20071_,
    new_n20072_, new_n20073_, new_n20074_, new_n20075_, new_n20076_,
    new_n20077_, new_n20078_, new_n20079_, new_n20080_, new_n20081_,
    new_n20082_, new_n20083_, new_n20084_, new_n20085_, new_n20086_,
    new_n20087_, new_n20088_, new_n20089_, new_n20090_, new_n20091_,
    new_n20092_, new_n20093_, new_n20094_, new_n20095_, new_n20096_,
    new_n20097_, new_n20098_, new_n20099_, new_n20100_, new_n20101_,
    new_n20102_, new_n20103_, new_n20104_, new_n20105_, new_n20106_,
    new_n20107_, new_n20108_, new_n20109_, new_n20110_, new_n20111_,
    new_n20112_, new_n20113_, new_n20114_, new_n20115_, new_n20116_,
    new_n20117_, new_n20118_, new_n20119_, new_n20120_, new_n20121_,
    new_n20122_, new_n20123_, new_n20124_, new_n20125_, new_n20126_,
    new_n20127_, new_n20128_, new_n20129_, new_n20130_, new_n20131_,
    new_n20132_, new_n20133_, new_n20134_, new_n20135_, new_n20136_,
    new_n20137_, new_n20138_, new_n20139_, new_n20140_, new_n20141_,
    new_n20142_, new_n20143_, new_n20144_, new_n20145_, new_n20146_,
    new_n20147_, new_n20148_, new_n20149_, new_n20150_, new_n20151_,
    new_n20152_, new_n20153_, new_n20154_, new_n20155_, new_n20156_,
    new_n20157_, new_n20158_, new_n20159_, new_n20160_, new_n20161_,
    new_n20162_, new_n20163_, new_n20164_, new_n20165_, new_n20166_,
    new_n20167_, new_n20168_, new_n20169_, new_n20170_, new_n20171_,
    new_n20172_, new_n20173_, new_n20174_, new_n20175_, new_n20176_,
    new_n20177_, new_n20178_, new_n20179_, new_n20180_, new_n20181_,
    new_n20182_, new_n20183_, new_n20184_, new_n20185_, new_n20186_,
    new_n20187_, new_n20188_, new_n20189_, new_n20190_, new_n20191_,
    new_n20192_, new_n20193_, new_n20194_, new_n20195_, new_n20196_,
    new_n20197_, new_n20198_, new_n20199_, new_n20200_, new_n20201_,
    new_n20202_, new_n20203_, new_n20204_, new_n20205_, new_n20206_,
    new_n20207_, new_n20208_, new_n20209_, new_n20210_, new_n20211_,
    new_n20212_, new_n20213_, new_n20214_, new_n20215_, new_n20216_,
    new_n20217_, new_n20218_, new_n20219_, new_n20220_, new_n20221_,
    new_n20222_, new_n20223_, new_n20224_, new_n20225_, new_n20226_,
    new_n20227_, new_n20228_, new_n20229_, new_n20230_, new_n20231_,
    new_n20232_, new_n20233_, new_n20234_, new_n20235_, new_n20236_,
    new_n20237_, new_n20238_, new_n20239_, new_n20240_, new_n20241_,
    new_n20242_, new_n20243_, new_n20244_, new_n20245_, new_n20246_,
    new_n20247_, new_n20248_, new_n20249_, new_n20250_, new_n20251_,
    new_n20252_, new_n20253_, new_n20254_, new_n20255_, new_n20256_,
    new_n20257_, new_n20258_, new_n20259_, new_n20260_, new_n20261_,
    new_n20262_, new_n20263_, new_n20264_, new_n20265_, new_n20266_,
    new_n20267_, new_n20268_, new_n20269_, new_n20270_, new_n20271_,
    new_n20272_, new_n20273_, new_n20274_, new_n20275_, new_n20276_,
    new_n20277_, new_n20278_, new_n20279_, new_n20280_, new_n20281_,
    new_n20282_, new_n20283_, new_n20284_, new_n20285_, new_n20286_,
    new_n20287_, new_n20288_, new_n20289_, new_n20290_, new_n20291_,
    new_n20292_, new_n20293_, new_n20294_, new_n20295_, new_n20296_,
    new_n20297_, new_n20298_, new_n20299_, new_n20300_, new_n20301_,
    new_n20302_, new_n20303_, new_n20304_, new_n20305_, new_n20306_,
    new_n20307_, new_n20308_, new_n20309_, new_n20310_, new_n20311_,
    new_n20312_, new_n20313_, new_n20314_, new_n20315_, new_n20316_,
    new_n20317_, new_n20318_, new_n20319_, new_n20320_, new_n20321_,
    new_n20322_, new_n20323_, new_n20324_, new_n20325_, new_n20326_,
    new_n20327_, new_n20328_, new_n20329_, new_n20330_, new_n20331_,
    new_n20332_, new_n20333_, new_n20334_, new_n20335_, new_n20336_,
    new_n20337_, new_n20338_, new_n20339_, new_n20340_, new_n20341_,
    new_n20342_, new_n20343_, new_n20344_, new_n20345_, new_n20346_,
    new_n20347_, new_n20348_, new_n20349_, new_n20350_, new_n20351_,
    new_n20352_, new_n20353_, new_n20354_, new_n20355_, new_n20356_,
    new_n20357_, new_n20358_, new_n20359_, new_n20360_, new_n20361_,
    new_n20362_, new_n20363_, new_n20364_, new_n20365_, new_n20366_,
    new_n20367_, new_n20368_, new_n20369_, new_n20370_, new_n20371_,
    new_n20372_, new_n20373_, new_n20374_, new_n20375_, new_n20376_,
    new_n20377_, new_n20378_, new_n20379_, new_n20380_, new_n20381_,
    new_n20382_, new_n20383_, new_n20384_, new_n20385_, new_n20386_,
    new_n20387_, new_n20388_, new_n20389_, new_n20390_, new_n20391_,
    new_n20392_, new_n20393_, new_n20394_, new_n20395_, new_n20396_,
    new_n20397_, new_n20398_, new_n20399_, new_n20400_, new_n20401_,
    new_n20402_, new_n20403_, new_n20404_, new_n20405_, new_n20406_,
    new_n20407_, new_n20408_, new_n20409_, new_n20410_, new_n20411_,
    new_n20412_, new_n20413_, new_n20414_, new_n20415_, new_n20416_,
    new_n20417_, new_n20418_, new_n20419_, new_n20420_, new_n20421_,
    new_n20422_, new_n20423_, new_n20424_, new_n20425_, new_n20426_,
    new_n20427_, new_n20428_, new_n20429_, new_n20430_, new_n20431_,
    new_n20432_, new_n20433_, new_n20434_, new_n20435_, new_n20436_,
    new_n20437_, new_n20438_, new_n20439_, new_n20440_, new_n20441_,
    new_n20442_, new_n20443_, new_n20444_, new_n20445_, new_n20446_,
    new_n20447_, new_n20448_, new_n20449_, new_n20450_, new_n20451_,
    new_n20452_, new_n20453_, new_n20454_, new_n20455_, new_n20456_,
    new_n20457_, new_n20458_, new_n20459_, new_n20460_, new_n20461_,
    new_n20462_, new_n20463_, new_n20464_, new_n20465_, new_n20466_,
    new_n20467_, new_n20468_, new_n20469_, new_n20470_, new_n20471_,
    new_n20472_, new_n20473_, new_n20474_, new_n20475_, new_n20476_,
    new_n20477_, new_n20478_, new_n20479_, new_n20480_, new_n20481_,
    new_n20482_, new_n20483_, new_n20484_, new_n20485_, new_n20486_,
    new_n20487_, new_n20488_, new_n20489_, new_n20490_, new_n20491_,
    new_n20492_, new_n20493_, new_n20494_, new_n20495_, new_n20496_,
    new_n20497_, new_n20498_, new_n20499_, new_n20500_, new_n20501_,
    new_n20502_, new_n20503_, new_n20504_, new_n20505_, new_n20506_,
    new_n20507_, new_n20508_, new_n20509_, new_n20510_, new_n20511_,
    new_n20512_, new_n20513_, new_n20514_, new_n20515_, new_n20516_,
    new_n20517_, new_n20518_, new_n20519_, new_n20520_, new_n20521_,
    new_n20522_, new_n20523_, new_n20524_, new_n20525_, new_n20526_,
    new_n20527_, new_n20528_, new_n20529_, new_n20530_, new_n20531_,
    new_n20532_, new_n20533_, new_n20534_, new_n20535_, new_n20536_,
    new_n20537_, new_n20538_, new_n20539_, new_n20540_, new_n20541_,
    new_n20542_, new_n20543_, new_n20544_, new_n20545_, new_n20546_,
    new_n20547_, new_n20548_, new_n20549_, new_n20550_, new_n20551_,
    new_n20552_, new_n20553_, new_n20554_, new_n20555_, new_n20556_,
    new_n20557_, new_n20558_, new_n20559_, new_n20560_, new_n20561_,
    new_n20562_, new_n20563_, new_n20564_, new_n20565_, new_n20566_,
    new_n20567_, new_n20568_, new_n20569_, new_n20570_, new_n20571_,
    new_n20572_, new_n20573_, new_n20574_, new_n20575_, new_n20576_,
    new_n20577_, new_n20578_, new_n20579_, new_n20580_, new_n20581_,
    new_n20582_, new_n20583_, new_n20584_, new_n20585_, new_n20586_,
    new_n20587_, new_n20588_, new_n20589_, new_n20590_, new_n20591_,
    new_n20592_, new_n20593_, new_n20594_, new_n20595_, new_n20596_,
    new_n20597_, new_n20598_, new_n20599_, new_n20600_, new_n20601_,
    new_n20602_, new_n20603_, new_n20604_, new_n20605_, new_n20606_,
    new_n20607_, new_n20608_, new_n20609_, new_n20610_, new_n20611_,
    new_n20612_, new_n20613_, new_n20614_, new_n20615_, new_n20616_,
    new_n20617_, new_n20618_, new_n20619_, new_n20620_, new_n20621_,
    new_n20622_, new_n20623_, new_n20624_, new_n20625_, new_n20626_,
    new_n20627_, new_n20628_, new_n20629_, new_n20630_, new_n20631_,
    new_n20632_, new_n20633_, new_n20634_, new_n20635_, new_n20636_,
    new_n20637_, new_n20638_, new_n20639_, new_n20640_, new_n20641_,
    new_n20642_, new_n20643_, new_n20644_, new_n20645_, new_n20646_,
    new_n20647_, new_n20648_, new_n20649_, new_n20650_, new_n20651_,
    new_n20652_, new_n20653_, new_n20654_, new_n20655_, new_n20656_,
    new_n20657_, new_n20658_, new_n20659_, new_n20660_, new_n20661_,
    new_n20662_, new_n20663_, new_n20664_, new_n20665_, new_n20666_,
    new_n20667_, new_n20668_, new_n20669_, new_n20670_, new_n20671_,
    new_n20672_, new_n20673_, new_n20674_, new_n20675_, new_n20676_,
    new_n20677_, new_n20678_, new_n20679_, new_n20680_, new_n20681_,
    new_n20682_, new_n20683_, new_n20684_, new_n20685_, new_n20686_,
    new_n20687_, new_n20688_, new_n20689_, new_n20690_, new_n20691_,
    new_n20692_, new_n20693_, new_n20694_, new_n20695_, new_n20696_,
    new_n20697_, new_n20698_, new_n20699_, new_n20700_, new_n20701_,
    new_n20702_, new_n20703_, new_n20704_, new_n20705_, new_n20706_,
    new_n20707_, new_n20708_, new_n20709_, new_n20710_, new_n20711_,
    new_n20712_, new_n20713_, new_n20714_, new_n20715_, new_n20716_,
    new_n20717_, new_n20718_, new_n20719_, new_n20720_, new_n20721_,
    new_n20722_, new_n20723_, new_n20724_, new_n20725_, new_n20726_,
    new_n20727_, new_n20728_, new_n20729_, new_n20730_, new_n20731_,
    new_n20732_, new_n20733_, new_n20734_, new_n20735_, new_n20736_,
    new_n20737_, new_n20738_, new_n20739_, new_n20740_, new_n20741_,
    new_n20742_, new_n20743_, new_n20744_, new_n20745_, new_n20746_,
    new_n20747_, new_n20748_, new_n20749_, new_n20750_, new_n20751_,
    new_n20752_, new_n20753_, new_n20754_, new_n20755_, new_n20756_,
    new_n20757_, new_n20758_, new_n20759_, new_n20760_, new_n20761_,
    new_n20762_, new_n20763_, new_n20764_, new_n20765_, new_n20766_,
    new_n20767_, new_n20768_, new_n20769_, new_n20770_, new_n20771_,
    new_n20772_, new_n20773_, new_n20774_, new_n20775_, new_n20776_,
    new_n20777_, new_n20778_, new_n20779_, new_n20780_, new_n20781_,
    new_n20782_, new_n20783_, new_n20784_, new_n20785_, new_n20786_,
    new_n20787_, new_n20788_, new_n20789_, new_n20790_, new_n20791_,
    new_n20792_, new_n20793_, new_n20794_, new_n20795_, new_n20796_,
    new_n20797_, new_n20798_, new_n20799_, new_n20800_, new_n20801_,
    new_n20802_, new_n20803_, new_n20804_, new_n20805_, new_n20806_,
    new_n20807_, new_n20808_, new_n20809_, new_n20810_, new_n20811_,
    new_n20812_, new_n20813_, new_n20814_, new_n20815_, new_n20816_,
    new_n20817_, new_n20818_, new_n20819_, new_n20820_, new_n20821_,
    new_n20822_, new_n20823_, new_n20824_, new_n20825_, new_n20826_,
    new_n20827_, new_n20828_, new_n20829_, new_n20830_, new_n20831_,
    new_n20832_, new_n20833_, new_n20834_, new_n20835_, new_n20836_,
    new_n20837_, new_n20838_, new_n20839_, new_n20840_, new_n20841_,
    new_n20842_, new_n20843_, new_n20844_, new_n20845_, new_n20846_,
    new_n20847_, new_n20848_, new_n20849_, new_n20850_, new_n20851_,
    new_n20852_, new_n20853_, new_n20854_, new_n20855_, new_n20856_,
    new_n20857_, new_n20858_, new_n20859_, new_n20860_, new_n20861_,
    new_n20862_, new_n20863_, new_n20864_, new_n20865_, new_n20866_,
    new_n20867_, new_n20868_, new_n20869_, new_n20870_, new_n20871_,
    new_n20872_, new_n20873_, new_n20874_, new_n20875_, new_n20876_,
    new_n20877_, new_n20878_, new_n20879_, new_n20880_, new_n20881_,
    new_n20882_, new_n20883_, new_n20884_, new_n20885_, new_n20886_,
    new_n20887_, new_n20888_, new_n20889_, new_n20890_, new_n20891_,
    new_n20892_, new_n20893_, new_n20894_, new_n20895_, new_n20896_,
    new_n20897_, new_n20898_, new_n20899_, new_n20900_, new_n20901_,
    new_n20902_, new_n20903_, new_n20904_, new_n20905_, new_n20906_,
    new_n20907_, new_n20908_, new_n20909_, new_n20910_, new_n20911_,
    new_n20912_, new_n20913_, new_n20914_, new_n20915_, new_n20916_,
    new_n20917_, new_n20918_, new_n20919_, new_n20920_, new_n20921_,
    new_n20922_, new_n20923_, new_n20924_, new_n20925_, new_n20926_,
    new_n20927_, new_n20928_, new_n20929_, new_n20930_, new_n20931_,
    new_n20932_, new_n20933_, new_n20934_, new_n20935_, new_n20936_,
    new_n20937_, new_n20938_, new_n20939_, new_n20940_, new_n20941_,
    new_n20942_, new_n20943_, new_n20944_, new_n20945_, new_n20946_,
    new_n20947_, new_n20948_, new_n20949_, new_n20950_, new_n20951_,
    new_n20952_, new_n20953_, new_n20954_, new_n20955_, new_n20956_,
    new_n20957_, new_n20958_, new_n20959_, new_n20960_, new_n20961_,
    new_n20962_, new_n20963_, new_n20964_, new_n20965_, new_n20966_,
    new_n20967_, new_n20968_, new_n20969_, new_n20970_, new_n20971_,
    new_n20972_, new_n20973_, new_n20974_, new_n20975_, new_n20976_,
    new_n20977_, new_n20978_, new_n20979_, new_n20980_, new_n20981_,
    new_n20982_, new_n20983_, new_n20984_, new_n20985_, new_n20986_,
    new_n20987_, new_n20988_, new_n20989_, new_n20990_, new_n20991_,
    new_n20992_, new_n20993_, new_n20994_, new_n20995_, new_n20996_,
    new_n20997_, new_n20998_, new_n20999_, new_n21000_, new_n21001_,
    new_n21002_, new_n21003_, new_n21004_, new_n21005_, new_n21006_,
    new_n21007_, new_n21008_, new_n21009_, new_n21010_, new_n21011_,
    new_n21012_, new_n21013_, new_n21014_, new_n21015_, new_n21016_,
    new_n21017_, new_n21018_, new_n21019_, new_n21020_, new_n21021_,
    new_n21022_, new_n21023_, new_n21024_, new_n21025_, new_n21026_,
    new_n21027_, new_n21028_, new_n21029_, new_n21030_, new_n21031_,
    new_n21032_, new_n21033_, new_n21034_, new_n21035_, new_n21036_,
    new_n21037_, new_n21038_, new_n21039_, new_n21040_, new_n21041_,
    new_n21042_, new_n21043_, new_n21044_, new_n21045_, new_n21046_,
    new_n21047_, new_n21048_, new_n21049_, new_n21050_, new_n21051_,
    new_n21052_, new_n21053_, new_n21054_, new_n21055_, new_n21056_,
    new_n21057_, new_n21058_, new_n21059_, new_n21071_, new_n21072_,
    new_n21073_, new_n21075_, new_n21076_, new_n21077_, new_n21078_,
    new_n21079_, new_n21080_, new_n21081_, new_n21082_, new_n21083_,
    new_n21084_, new_n21085_, new_n21086_, new_n21087_, new_n21088_,
    new_n21089_, new_n21090_, new_n21091_, new_n21092_, new_n21093_,
    new_n21094_, new_n21095_, new_n21096_, new_n21097_, new_n21098_,
    new_n21099_, new_n21100_, new_n21101_, new_n21102_, new_n21103_,
    new_n21104_, new_n21105_, new_n21106_, new_n21107_, new_n21108_,
    new_n21109_, new_n21111_, new_n21112_, new_n21113_, new_n21114_,
    new_n21115_, new_n21116_, new_n21117_, new_n21118_, new_n21119_,
    new_n21120_, new_n21121_, new_n21122_, new_n21123_, new_n21124_,
    new_n21125_, new_n21126_, new_n21127_, new_n21128_, new_n21129_,
    new_n21130_, new_n21131_, new_n21132_, new_n21133_, new_n21134_,
    new_n21135_, new_n21136_, new_n21137_, new_n21138_, new_n21139_,
    new_n21140_, new_n21141_, new_n21142_, new_n21143_, new_n21144_,
    new_n21145_, new_n21146_, new_n21147_, new_n21148_, new_n21149_,
    new_n21150_, new_n21151_, new_n21152_, new_n21153_, new_n21154_,
    new_n21155_, new_n21156_, new_n21157_, new_n21158_, new_n21159_,
    new_n21160_, new_n21161_, new_n21162_, new_n21163_, new_n21164_,
    new_n21165_, new_n21166_, new_n21167_, new_n21168_, new_n21169_,
    new_n21170_, new_n21171_, new_n21172_, new_n21173_, new_n21174_,
    new_n21175_, new_n21176_, new_n21177_, new_n21178_, new_n21179_,
    new_n21180_, new_n21181_, new_n21182_, new_n21183_, new_n21184_,
    new_n21185_, new_n21186_, new_n21187_, new_n21188_, new_n21189_,
    new_n21190_, new_n21191_, new_n21192_, new_n21193_, new_n21194_,
    new_n21195_, new_n21196_, new_n21197_, new_n21198_, new_n21199_,
    new_n21200_, new_n21201_, new_n21202_, new_n21203_, new_n21204_,
    new_n21205_, new_n21206_, new_n21207_, new_n21208_, new_n21209_,
    new_n21210_, new_n21211_, new_n21212_, new_n21213_, new_n21214_,
    new_n21215_, new_n21216_, new_n21217_, new_n21218_, new_n21219_,
    new_n21220_, new_n21221_, new_n21222_, new_n21223_, new_n21224_,
    new_n21225_, new_n21226_, new_n21227_, new_n21228_, new_n21229_,
    new_n21230_, new_n21231_, new_n21232_, new_n21233_, new_n21234_,
    new_n21235_, new_n21236_, new_n21237_, new_n21238_, new_n21239_,
    new_n21240_, new_n21241_, new_n21242_, new_n21243_, new_n21244_,
    new_n21245_, new_n21246_, new_n21247_, new_n21248_, new_n21249_,
    new_n21250_, new_n21251_, new_n21252_, new_n21253_, new_n21254_,
    new_n21255_, new_n21256_, new_n21257_, new_n21258_, new_n21259_,
    new_n21260_, new_n21261_, new_n21262_, new_n21263_, new_n21264_,
    new_n21265_, new_n21266_, new_n21267_, new_n21268_, new_n21269_,
    new_n21270_, new_n21271_, new_n21272_, new_n21273_, new_n21274_,
    new_n21275_, new_n21276_, new_n21277_, new_n21278_, new_n21279_,
    new_n21280_, new_n21281_, new_n21282_, new_n21283_, new_n21284_,
    new_n21285_, new_n21286_, new_n21287_, new_n21288_, new_n21289_,
    new_n21290_, new_n21291_, new_n21292_, new_n21293_, new_n21294_,
    new_n21295_, new_n21296_, new_n21297_, new_n21298_, new_n21299_,
    new_n21300_, new_n21301_, new_n21302_, new_n21303_, new_n21304_,
    new_n21305_, new_n21306_, new_n21307_, new_n21308_, new_n21309_,
    new_n21310_, new_n21311_, new_n21312_, new_n21313_, new_n21314_,
    new_n21315_, new_n21316_, new_n21317_, new_n21318_, new_n21319_,
    new_n21320_, new_n21321_, new_n21322_, new_n21323_, new_n21324_,
    new_n21325_, new_n21326_, new_n21327_, new_n21328_, new_n21329_,
    new_n21330_, new_n21331_, new_n21332_, new_n21333_, new_n21334_,
    new_n21335_, new_n21336_, new_n21337_, new_n21338_, new_n21339_,
    new_n21340_, new_n21341_, new_n21342_, new_n21343_, new_n21344_,
    new_n21345_, new_n21346_, new_n21347_, new_n21348_, new_n21349_,
    new_n21350_, new_n21351_, new_n21352_, new_n21353_, new_n21354_,
    new_n21355_, new_n21356_, new_n21357_, new_n21358_, new_n21359_,
    new_n21360_, new_n21361_, new_n21362_, new_n21363_, new_n21364_,
    new_n21365_, new_n21366_, new_n21367_, new_n21368_, new_n21369_,
    new_n21370_, new_n21371_, new_n21372_, new_n21373_, new_n21374_,
    new_n21375_, new_n21376_, new_n21377_, new_n21378_, new_n21379_,
    new_n21380_, new_n21381_, new_n21382_, new_n21383_, new_n21384_,
    new_n21385_, new_n21387_, new_n21388_, new_n21389_, new_n21390_,
    new_n21391_, new_n21392_, new_n21393_, new_n21394_, new_n21395_,
    new_n21396_, new_n21397_, new_n21398_, new_n21399_, new_n21400_,
    new_n21401_, new_n21402_, new_n21403_, new_n21404_, new_n21405_,
    new_n21406_, new_n21407_, new_n21408_, new_n21409_, new_n21410_,
    new_n21411_, new_n21412_, new_n21413_, new_n21414_, new_n21415_,
    new_n21416_, new_n21417_, new_n21418_, new_n21419_, new_n21420_,
    new_n21421_, new_n21422_, new_n21423_, new_n21424_, new_n21425_,
    new_n21426_, new_n21427_, new_n21428_, new_n21429_, new_n21430_,
    new_n21431_, new_n21432_, new_n21433_, new_n21434_, new_n21435_,
    new_n21436_, new_n21437_, new_n21438_, new_n21439_, new_n21440_,
    new_n21441_, new_n21442_, new_n21443_, new_n21444_, new_n21445_,
    new_n21446_, new_n21447_, new_n21448_, new_n21449_, new_n21450_,
    new_n21451_, new_n21452_, new_n21453_, new_n21454_, new_n21455_,
    new_n21456_, new_n21457_, new_n21458_, new_n21459_, new_n21460_,
    new_n21461_, new_n21462_, new_n21463_, new_n21464_, new_n21465_,
    new_n21466_, new_n21467_, new_n21468_, new_n21469_, new_n21470_,
    new_n21471_, new_n21472_, new_n21473_, new_n21474_, new_n21475_,
    new_n21476_, new_n21477_, new_n21478_, new_n21479_, new_n21480_,
    new_n21481_, new_n21482_, new_n21483_, new_n21484_, new_n21485_,
    new_n21486_, new_n21487_, new_n21488_, new_n21489_, new_n21490_,
    new_n21491_, new_n21492_, new_n21493_, new_n21494_, new_n21495_,
    new_n21496_, new_n21497_, new_n21498_, new_n21499_, new_n21500_,
    new_n21501_, new_n21502_, new_n21503_, new_n21504_, new_n21505_,
    new_n21506_, new_n21507_, new_n21508_, new_n21509_, new_n21510_,
    new_n21511_, new_n21512_, new_n21513_, new_n21514_, new_n21515_,
    new_n21516_, new_n21517_, new_n21518_, new_n21519_, new_n21520_,
    new_n21521_, new_n21522_, new_n21523_, new_n21524_, new_n21525_,
    new_n21526_, new_n21527_, new_n21528_, new_n21529_, new_n21530_,
    new_n21531_, new_n21532_, new_n21533_, new_n21534_, new_n21535_,
    new_n21536_, new_n21537_, new_n21538_, new_n21539_, new_n21540_,
    new_n21541_, new_n21542_, new_n21543_, new_n21544_, new_n21545_,
    new_n21546_, new_n21547_, new_n21548_, new_n21549_, new_n21550_,
    new_n21551_, new_n21552_, new_n21553_, new_n21554_, new_n21555_,
    new_n21556_, new_n21557_, new_n21558_, new_n21559_, new_n21560_,
    new_n21561_, new_n21562_, new_n21563_, new_n21564_, new_n21565_,
    new_n21566_, new_n21567_, new_n21568_, new_n21569_, new_n21570_,
    new_n21571_, new_n21572_, new_n21573_, new_n21574_, new_n21575_,
    new_n21576_, new_n21577_, new_n21578_, new_n21579_, new_n21580_,
    new_n21581_, new_n21582_, new_n21583_, new_n21584_, new_n21585_,
    new_n21586_, new_n21587_, new_n21588_, new_n21589_, new_n21590_,
    new_n21591_, new_n21592_, new_n21593_, new_n21594_, new_n21595_,
    new_n21596_, new_n21597_, new_n21598_, new_n21599_, new_n21600_,
    new_n21601_, new_n21602_, new_n21603_, new_n21604_, new_n21605_,
    new_n21606_, new_n21607_, new_n21608_, new_n21609_, new_n21610_,
    new_n21611_, new_n21612_, new_n21613_, new_n21614_, new_n21615_,
    new_n21616_, new_n21617_, new_n21618_, new_n21619_, new_n21620_,
    new_n21621_, new_n21622_, new_n21623_, new_n21624_, new_n21625_,
    new_n21626_, new_n21627_, new_n21628_, new_n21629_, new_n21630_,
    new_n21631_, new_n21632_, new_n21633_, new_n21634_, new_n21635_,
    new_n21636_, new_n21637_, new_n21638_, new_n21639_, new_n21640_,
    new_n21641_, new_n21642_, new_n21643_, new_n21644_, new_n21645_,
    new_n21646_, new_n21647_, new_n21648_, new_n21649_, new_n21650_,
    new_n21651_, new_n21652_, new_n21653_, new_n21654_, new_n21655_,
    new_n21656_, new_n21657_, new_n21658_, new_n21659_, new_n21660_,
    new_n21661_, new_n21662_, new_n21663_, new_n21664_, new_n21665_,
    new_n21666_, new_n21667_, new_n21668_, new_n21669_, new_n21670_,
    new_n21671_, new_n21672_, new_n21673_, new_n21674_, new_n21675_,
    new_n21676_, new_n21677_, new_n21678_, new_n21679_, new_n21680_,
    new_n21681_, new_n21682_, new_n21683_, new_n21684_, new_n21685_,
    new_n21686_, new_n21687_, new_n21688_, new_n21689_, new_n21690_,
    new_n21691_, new_n21692_, new_n21693_, new_n21694_, new_n21695_,
    new_n21696_, new_n21697_, new_n21698_, new_n21699_, new_n21700_,
    new_n21701_, new_n21702_, new_n21703_, new_n21704_, new_n21705_,
    new_n21706_, new_n21707_, new_n21708_, new_n21709_, new_n21710_,
    new_n21711_, new_n21712_, new_n21713_, new_n21714_, new_n21715_,
    new_n21716_, new_n21717_, new_n21718_, new_n21719_, new_n21720_,
    new_n21721_, new_n21722_, new_n21723_, new_n21724_, new_n21725_,
    new_n21726_, new_n21727_, new_n21728_, new_n21729_, new_n21730_,
    new_n21731_, new_n21732_, new_n21733_, new_n21734_, new_n21735_,
    new_n21736_, new_n21737_, new_n21738_, new_n21739_, new_n21740_,
    new_n21741_, new_n21742_, new_n21743_, new_n21744_, new_n21745_,
    new_n21746_, new_n21747_, new_n21748_, new_n21749_, new_n21750_,
    new_n21751_, new_n21752_, new_n21753_, new_n21754_, new_n21755_,
    new_n21756_, new_n21757_, new_n21758_, new_n21759_, new_n21760_,
    new_n21761_, new_n21762_, new_n21763_, new_n21764_, new_n21765_,
    new_n21766_, new_n21767_, new_n21768_, new_n21769_, new_n21770_,
    new_n21771_, new_n21772_, new_n21773_, new_n21774_, new_n21775_,
    new_n21776_, new_n21777_, new_n21778_, new_n21779_, new_n21780_,
    new_n21781_, new_n21782_, new_n21783_, new_n21784_, new_n21785_,
    new_n21786_, new_n21787_, new_n21788_, new_n21789_, new_n21790_,
    new_n21791_, new_n21792_, new_n21793_, new_n21794_, new_n21795_,
    new_n21796_, new_n21797_, new_n21798_, new_n21799_, new_n21800_,
    new_n21801_, new_n21802_, new_n21803_, new_n21804_, new_n21805_,
    new_n21806_, new_n21807_, new_n21808_, new_n21809_, new_n21810_,
    new_n21811_, new_n21812_, new_n21813_, new_n21814_, new_n21815_,
    new_n21816_, new_n21817_, new_n21818_, new_n21819_, new_n21820_,
    new_n21821_, new_n21822_, new_n21823_, new_n21824_, new_n21825_,
    new_n21826_, new_n21827_, new_n21828_, new_n21829_, new_n21830_,
    new_n21831_, new_n21832_, new_n21833_, new_n21834_, new_n21835_,
    new_n21836_, new_n21837_, new_n21838_, new_n21839_, new_n21840_,
    new_n21841_, new_n21842_, new_n21843_, new_n21844_, new_n21845_,
    new_n21846_, new_n21847_, new_n21848_, new_n21849_, new_n21850_,
    new_n21851_, new_n21852_, new_n21853_, new_n21854_, new_n21855_,
    new_n21856_, new_n21857_, new_n21858_, new_n21859_, new_n21860_,
    new_n21861_, new_n21862_, new_n21863_, new_n21864_, new_n21865_,
    new_n21866_, new_n21867_, new_n21868_, new_n21869_, new_n21870_,
    new_n21871_, new_n21872_, new_n21873_, new_n21874_, new_n21875_,
    new_n21876_, new_n21877_, new_n21878_, new_n21879_, new_n21880_,
    new_n21881_, new_n21882_, new_n21883_, new_n21884_, new_n21885_,
    new_n21886_, new_n21887_, new_n21888_, new_n21889_, new_n21890_,
    new_n21891_, new_n21892_, new_n21893_, new_n21894_, new_n21895_,
    new_n21896_, new_n21897_, new_n21898_, new_n21899_, new_n21900_,
    new_n21901_, new_n21902_, new_n21903_, new_n21904_, new_n21905_,
    new_n21906_, new_n21907_, new_n21908_, new_n21909_, new_n21910_,
    new_n21911_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21939_, new_n21940_, new_n21941_, new_n21944_,
    new_n21945_, new_n21946_, new_n21947_, new_n21948_, new_n21949_,
    new_n21950_, new_n21951_, new_n21952_, new_n21953_, new_n21954_,
    new_n21955_, new_n21956_, new_n21957_, new_n21958_, new_n21959_,
    new_n21960_, new_n21961_, new_n21962_, new_n21963_, new_n21964_,
    new_n21965_, new_n21966_, new_n21967_, new_n21968_, new_n21969_,
    new_n21970_, new_n21971_, new_n21972_, new_n21973_, new_n21974_,
    new_n21975_, new_n21976_, new_n21977_, new_n21978_, new_n21979_,
    new_n21980_, new_n21981_, new_n21982_, new_n21983_, new_n21984_,
    new_n21985_, new_n21986_, new_n21987_, new_n21988_, new_n21989_,
    new_n21990_, new_n21991_, new_n21992_, new_n21993_, new_n21994_,
    new_n21995_, new_n21996_, new_n21997_, new_n21998_, new_n21999_,
    new_n22000_, new_n22001_, new_n22002_, new_n22003_, new_n22004_,
    new_n22005_, new_n22006_, new_n22007_, new_n22008_, new_n22009_,
    new_n22010_, new_n22011_, new_n22012_, new_n22013_, new_n22014_,
    new_n22015_, new_n22016_, new_n22017_, new_n22018_, new_n22019_,
    new_n22020_, new_n22021_, new_n22022_, new_n22023_, new_n22024_,
    new_n22025_, new_n22026_, new_n22027_, new_n22028_, new_n22029_,
    new_n22030_, new_n22031_, new_n22032_, new_n22033_, new_n22034_,
    new_n22035_, new_n22036_, new_n22037_, new_n22038_, new_n22039_,
    new_n22040_, new_n22041_, new_n22042_, new_n22043_, new_n22044_,
    new_n22045_, new_n22046_, new_n22047_, new_n22048_, new_n22049_,
    new_n22050_, new_n22051_, new_n22052_, new_n22053_, new_n22054_,
    new_n22055_, new_n22056_, new_n22057_, new_n22058_, new_n22059_,
    new_n22060_, new_n22061_, new_n22062_, new_n22063_, new_n22064_,
    new_n22065_, new_n22066_, new_n22067_, new_n22068_, new_n22069_,
    new_n22070_, new_n22071_, new_n22072_, new_n22073_, new_n22074_,
    new_n22075_, new_n22076_, new_n22077_, new_n22078_, new_n22079_,
    new_n22080_, new_n22081_, new_n22082_, new_n22083_, new_n22085_,
    new_n22086_, new_n22087_, new_n22088_, new_n22089_, new_n22090_,
    new_n22091_, new_n22092_, new_n22093_, new_n22094_, new_n22095_,
    new_n22096_, new_n22097_, new_n22098_, new_n22099_, new_n22100_,
    new_n22101_, new_n22102_, new_n22103_, new_n22104_, new_n22105_,
    new_n22106_, new_n22107_, new_n22108_, new_n22109_, new_n22110_,
    new_n22111_, new_n22112_, new_n22113_, new_n22114_, new_n22115_,
    new_n22116_, new_n22117_, new_n22118_, new_n22119_, new_n22120_,
    new_n22121_, new_n22122_, new_n22123_, new_n22124_, new_n22125_,
    new_n22126_, new_n22127_, new_n22128_, new_n22129_, new_n22130_,
    new_n22131_, new_n22132_, new_n22133_, new_n22134_, new_n22135_,
    new_n22136_, new_n22137_, new_n22138_, new_n22139_, new_n22140_,
    new_n22141_, new_n22142_, new_n22143_, new_n22144_, new_n22145_,
    new_n22146_, new_n22147_, new_n22148_, new_n22149_, new_n22150_,
    new_n22151_, new_n22152_, new_n22153_, new_n22154_, new_n22155_,
    new_n22156_, new_n22157_, new_n22158_, new_n22159_, new_n22160_,
    new_n22161_, new_n22162_, new_n22163_, new_n22164_, new_n22165_,
    new_n22166_, new_n22167_, new_n22168_, new_n22169_, new_n22170_,
    new_n22171_, new_n22172_, new_n22173_, new_n22174_, new_n22175_,
    new_n22176_, new_n22177_, new_n22178_, new_n22179_, new_n22180_,
    new_n22181_, new_n22182_, new_n22183_, new_n22184_, new_n22185_,
    new_n22186_, new_n22187_, new_n22188_, new_n22190_, new_n22191_,
    new_n22192_, new_n22193_, new_n22194_, new_n22195_, new_n22196_,
    new_n22197_, new_n22198_, new_n22199_, new_n22200_, new_n22201_,
    new_n22202_, new_n22203_, new_n22204_, new_n22205_, new_n22206_,
    new_n22207_, new_n22208_, new_n22209_, new_n22210_, new_n22211_,
    new_n22212_, new_n22213_, new_n22214_, new_n22215_, new_n22216_,
    new_n22217_, new_n22218_, new_n22219_, new_n22220_, new_n22221_,
    new_n22222_, new_n22223_, new_n22225_, new_n22226_, new_n22227_,
    new_n22228_, new_n22229_, new_n22230_, new_n22231_, new_n22232_,
    new_n22233_, new_n22234_, new_n22235_, new_n22236_, new_n22237_,
    new_n22238_, new_n22239_, new_n22240_, new_n22241_, new_n22242_,
    new_n22243_, new_n22244_, new_n22246_, new_n22247_, new_n22248_,
    new_n22249_, new_n22250_, new_n22251_, new_n22252_, new_n22253_,
    new_n22254_, new_n22255_, new_n22256_, new_n22258_, new_n22259_,
    new_n22260_, new_n22261_, new_n22262_, new_n22265_, new_n22266_,
    new_n22267_, new_n22268_, new_n22269_, new_n22270_, new_n22271_,
    new_n22272_, new_n22273_, new_n22274_, new_n22275_, new_n22276_,
    new_n22277_, new_n22278_, new_n22279_, new_n22280_, new_n22281_,
    new_n22282_, new_n22283_, new_n22284_, new_n22285_, new_n22286_,
    new_n22287_, new_n22288_, new_n22289_, new_n22290_, new_n22291_,
    new_n22292_, new_n22293_, new_n22294_, new_n22295_, new_n22296_,
    new_n22297_, new_n22298_, new_n22299_, new_n22300_, new_n22301_,
    new_n22302_, new_n22303_, new_n22304_, new_n22305_, new_n22306_,
    new_n22307_, new_n22308_, new_n22309_, new_n22310_, new_n22311_,
    new_n22312_, new_n22313_, new_n22314_, new_n22315_, new_n22316_,
    new_n22317_, new_n22318_, new_n22319_, new_n22320_, new_n22321_,
    new_n22322_, new_n22323_, new_n22324_, new_n22326_, new_n22327_,
    new_n22328_, new_n22329_, new_n22330_, new_n22331_, new_n22332_,
    new_n22333_, new_n22335_, new_n22336_, new_n22337_, new_n22338_,
    new_n22339_, new_n22340_, new_n22341_, new_n22342_, new_n22343_,
    new_n22344_, new_n22345_, new_n22346_, new_n22347_, new_n22348_,
    new_n22349_, new_n22350_, new_n22351_, new_n22352_, new_n22353_,
    new_n22354_, new_n22355_, new_n22356_, new_n22357_, new_n22358_,
    new_n22359_, new_n22360_, new_n22361_, new_n22362_, new_n22363_,
    new_n22364_, new_n22365_, new_n22366_, new_n22367_, new_n22368_,
    new_n22369_, new_n22370_, new_n22371_, new_n22372_, new_n22373_,
    new_n22374_, new_n22375_, new_n22376_, new_n22377_, new_n22378_,
    new_n22379_, new_n22380_, new_n22381_, new_n22382_, new_n22383_,
    new_n22384_, new_n22385_, new_n22386_, new_n22387_, new_n22388_,
    new_n22389_, new_n22390_, new_n22391_, new_n22392_, new_n22393_,
    new_n22394_, new_n22395_, new_n22396_, new_n22397_, new_n22398_,
    new_n22399_, new_n22400_, new_n22401_, new_n22402_, new_n22403_,
    new_n22404_, new_n22405_, new_n22406_, new_n22407_, new_n22408_,
    new_n22409_, new_n22410_, new_n22411_, new_n22412_, new_n22413_,
    new_n22414_, new_n22415_, new_n22416_, new_n22417_, new_n22418_,
    new_n22419_, new_n22420_, new_n22421_, new_n22422_, new_n22423_,
    new_n22424_, new_n22425_, new_n22426_, new_n22427_, new_n22428_,
    new_n22429_, new_n22430_, new_n22431_, new_n22432_, new_n22433_,
    new_n22434_, new_n22435_, new_n22436_, new_n22437_, new_n22438_,
    new_n22439_, new_n22440_, new_n22441_, new_n22442_, new_n22443_,
    new_n22444_, new_n22445_, new_n22446_, new_n22447_, new_n22448_,
    new_n22449_, new_n22450_, new_n22451_, new_n22452_, new_n22453_,
    new_n22454_, new_n22455_, new_n22456_, new_n22457_, new_n22458_,
    new_n22459_, new_n22460_, new_n22461_, new_n22462_, new_n22463_,
    new_n22464_, new_n22465_, new_n22466_, new_n22467_, new_n22468_,
    new_n22469_, new_n22470_, new_n22471_, new_n22472_, new_n22473_,
    new_n22474_, new_n22475_, new_n22476_, new_n22477_, new_n22478_,
    new_n22479_, new_n22480_, new_n22481_, new_n22482_, new_n22483_,
    new_n22484_, new_n22485_, new_n22486_, new_n22487_, new_n22488_,
    new_n22489_, new_n22490_, new_n22491_, new_n22492_, new_n22493_,
    new_n22494_, new_n22495_, new_n22496_, new_n22497_, new_n22498_,
    new_n22499_, new_n22500_, new_n22501_, new_n22502_, new_n22503_,
    new_n22504_, new_n22505_, new_n22506_, new_n22507_, new_n22508_,
    new_n22509_, new_n22510_, new_n22511_, new_n22512_, new_n22513_,
    new_n22514_, new_n22515_, new_n22516_, new_n22517_, new_n22518_,
    new_n22519_, new_n22520_, new_n22521_, new_n22522_, new_n22523_,
    new_n22524_, new_n22525_, new_n22526_, new_n22527_, new_n22528_,
    new_n22529_, new_n22530_, new_n22531_, new_n22532_, new_n22533_,
    new_n22534_, new_n22535_, new_n22536_, new_n22537_, new_n22538_,
    new_n22539_, new_n22540_, new_n22541_, new_n22542_, new_n22543_,
    new_n22544_, new_n22545_, new_n22546_, new_n22547_, new_n22548_,
    new_n22549_, new_n22550_, new_n22551_, new_n22552_, new_n22553_,
    new_n22554_, new_n22555_, new_n22556_, new_n22557_, new_n22558_,
    new_n22559_, new_n22560_, new_n22561_, new_n22562_, new_n22563_,
    new_n22564_, new_n22565_, new_n22566_, new_n22567_, new_n22568_,
    new_n22569_, new_n22570_, new_n22571_, new_n22572_, new_n22573_,
    new_n22574_, new_n22575_, new_n22576_, new_n22577_, new_n22578_,
    new_n22579_, new_n22580_, new_n22581_, new_n22582_, new_n22583_,
    new_n22584_, new_n22585_, new_n22586_, new_n22587_, new_n22588_,
    new_n22589_, new_n22590_, new_n22591_, new_n22592_, new_n22593_,
    new_n22594_, new_n22595_, new_n22596_, new_n22597_, new_n22598_,
    new_n22599_, new_n22600_, new_n22601_, new_n22602_, new_n22603_,
    new_n22604_, new_n22605_, new_n22606_, new_n22607_, new_n22608_,
    new_n22609_, new_n22610_, new_n22611_, new_n22612_, new_n22613_,
    new_n22614_, new_n22615_, new_n22616_, new_n22617_, new_n22618_,
    new_n22619_, new_n22620_, new_n22621_, new_n22622_, new_n22623_,
    new_n22624_, new_n22625_, new_n22626_, new_n22627_, new_n22628_,
    new_n22629_, new_n22630_, new_n22631_, new_n22632_, new_n22633_,
    new_n22634_, new_n22635_, new_n22636_, new_n22637_, new_n22638_,
    new_n22639_, new_n22640_, new_n22641_, new_n22642_, new_n22643_,
    new_n22644_, new_n22645_, new_n22646_, new_n22647_, new_n22648_,
    new_n22649_, new_n22650_, new_n22651_, new_n22652_, new_n22653_,
    new_n22654_, new_n22655_, new_n22656_, new_n22657_, new_n22658_,
    new_n22659_, new_n22660_, new_n22661_, new_n22662_, new_n22663_,
    new_n22664_, new_n22665_, new_n22666_, new_n22667_, new_n22668_,
    new_n22669_, new_n22670_, new_n22671_, new_n22672_, new_n22673_,
    new_n22674_, new_n22675_, new_n22676_, new_n22677_, new_n22678_,
    new_n22679_, new_n22680_, new_n22681_, new_n22682_, new_n22683_,
    new_n22684_, new_n22685_, new_n22686_, new_n22687_, new_n22688_,
    new_n22689_, new_n22690_, new_n22691_, new_n22692_, new_n22693_,
    new_n22694_, new_n22695_, new_n22696_, new_n22697_, new_n22698_,
    new_n22699_, new_n22700_, new_n22701_, new_n22702_, new_n22703_,
    new_n22704_, new_n22705_, new_n22706_, new_n22707_, new_n22708_,
    new_n22709_, new_n22710_, new_n22711_, new_n22712_, new_n22713_,
    new_n22714_, new_n22715_, new_n22716_, new_n22717_, new_n22718_,
    new_n22719_, new_n22720_, new_n22721_, new_n22722_, new_n22723_,
    new_n22724_, new_n22725_, new_n22726_, new_n22727_, new_n22728_,
    new_n22729_, new_n22730_, new_n22731_, new_n22732_, new_n22733_,
    new_n22734_, new_n22735_, new_n22736_, new_n22737_, new_n22738_,
    new_n22739_, new_n22740_, new_n22741_, new_n22742_, new_n22743_,
    new_n22744_, new_n22745_, new_n22746_, new_n22747_, new_n22748_,
    new_n22749_, new_n22750_, new_n22751_, new_n22752_, new_n22753_,
    new_n22754_, new_n22755_, new_n22756_, new_n22757_, new_n22758_,
    new_n22759_, new_n22761_, new_n22762_, new_n22763_, new_n22764_,
    new_n22767_, new_n22768_, new_n22769_, new_n22770_, new_n22771_,
    new_n22772_, new_n22773_, new_n22774_, new_n22775_, new_n22776_,
    new_n22777_, new_n22778_, new_n22779_, new_n22780_, new_n22781_,
    new_n22782_, new_n22783_, new_n22784_, new_n22785_, new_n22786_,
    new_n22787_, new_n22788_, new_n22789_, new_n22790_, new_n22791_,
    new_n22792_, new_n22793_, new_n22794_, new_n22795_, new_n22796_,
    new_n22797_, new_n22798_, new_n22799_, new_n22800_, new_n22801_,
    new_n22802_, new_n22803_, new_n22804_, new_n22805_, new_n22806_,
    new_n22807_, new_n22808_, new_n22809_, new_n22810_, new_n22811_,
    new_n22812_, new_n22813_, new_n22814_, new_n22815_, new_n22816_,
    new_n22817_, new_n22818_, new_n22819_, new_n22820_, new_n22821_,
    new_n22822_, new_n22823_, new_n22824_, new_n22825_, new_n22826_,
    new_n22827_, new_n22828_, new_n22829_, new_n22830_, new_n22831_,
    new_n22832_, new_n22833_, new_n22834_, new_n22835_, new_n22836_,
    new_n22837_, new_n22838_, new_n22839_, new_n22840_, new_n22841_,
    new_n22842_, new_n22843_, new_n22844_, new_n22845_, new_n22846_,
    new_n22847_, new_n22848_, new_n22849_, new_n22850_, new_n22851_,
    new_n22852_, new_n22853_, new_n22854_, new_n22855_, new_n22856_,
    new_n22857_, new_n22858_, new_n22859_, new_n22860_, new_n22861_,
    new_n22862_, new_n22863_, new_n22864_, new_n22865_, new_n22866_,
    new_n22867_, new_n22868_, new_n22869_, new_n22870_, new_n22871_,
    new_n22872_, new_n22873_, new_n22874_, new_n22875_, new_n22876_,
    new_n22877_, new_n22878_, new_n22879_, new_n22880_, new_n22881_,
    new_n22882_, new_n22883_, new_n22884_, new_n22885_, new_n22886_,
    new_n22887_, new_n22888_, new_n22889_, new_n22890_, new_n22891_,
    new_n22892_, new_n22893_, new_n22894_, new_n22895_, new_n22896_,
    new_n22897_, new_n22898_, new_n22899_, new_n22900_, new_n22901_,
    new_n22902_, new_n22903_, new_n22904_, new_n22905_, new_n22906_,
    new_n22907_, new_n22908_, new_n22909_, new_n22910_, new_n22911_,
    new_n22912_, new_n22913_, new_n22914_, new_n22915_, new_n22916_,
    new_n22917_, new_n22918_, new_n22919_, new_n22920_, new_n22921_,
    new_n22922_, new_n22923_, new_n22924_, new_n22925_, new_n22926_,
    new_n22927_, new_n22928_, new_n22929_, new_n22930_, new_n22931_,
    new_n22932_, new_n22933_, new_n22934_, new_n22935_, new_n22936_,
    new_n22937_, new_n22938_, new_n22939_, new_n22940_, new_n22941_,
    new_n22942_, new_n22943_, new_n22944_, new_n22945_, new_n22946_,
    new_n22947_, new_n22948_, new_n22949_, new_n22950_, new_n22951_,
    new_n22952_, new_n22953_, new_n22954_, new_n22955_, new_n22956_,
    new_n22957_, new_n22958_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23001_,
    new_n23002_, new_n23003_, new_n23004_, new_n23005_, new_n23006_,
    new_n23007_, new_n23008_, new_n23009_, new_n23010_, new_n23011_,
    new_n23012_, new_n23013_, new_n23014_, new_n23015_, new_n23016_,
    new_n23017_, new_n23018_, new_n23019_, new_n23020_, new_n23021_,
    new_n23022_, new_n23023_, new_n23024_, new_n23025_, new_n23026_,
    new_n23027_, new_n23028_, new_n23029_, new_n23030_, new_n23031_,
    new_n23032_, new_n23033_, new_n23034_, new_n23035_, new_n23036_,
    new_n23037_, new_n23038_, new_n23039_, new_n23040_, new_n23041_,
    new_n23042_, new_n23043_, new_n23044_, new_n23045_, new_n23046_,
    new_n23047_, new_n23048_, new_n23049_, new_n23050_, new_n23051_,
    new_n23052_, new_n23053_, new_n23054_, new_n23055_, new_n23056_,
    new_n23057_, new_n23058_, new_n23059_, new_n23060_, new_n23061_,
    new_n23062_, new_n23063_, new_n23064_, new_n23065_, new_n23066_,
    new_n23067_, new_n23068_, new_n23069_, new_n23070_, new_n23071_,
    new_n23072_, new_n23073_, new_n23074_, new_n23075_, new_n23076_,
    new_n23077_, new_n23078_, new_n23079_, new_n23080_, new_n23081_,
    new_n23082_, new_n23083_, new_n23084_, new_n23085_, new_n23086_,
    new_n23087_, new_n23088_, new_n23089_, new_n23090_, new_n23091_,
    new_n23092_, new_n23093_, new_n23094_, new_n23095_, new_n23096_,
    new_n23097_, new_n23098_, new_n23099_, new_n23100_, new_n23101_,
    new_n23102_, new_n23103_, new_n23104_, new_n23105_, new_n23106_,
    new_n23107_, new_n23108_, new_n23109_, new_n23110_, new_n23111_,
    new_n23112_, new_n23113_, new_n23114_, new_n23115_, new_n23116_,
    new_n23117_, new_n23118_, new_n23119_, new_n23120_, new_n23121_,
    new_n23122_, new_n23123_, new_n23124_, new_n23125_, new_n23126_,
    new_n23127_, new_n23128_, new_n23129_, new_n23130_, new_n23131_,
    new_n23132_, new_n23133_, new_n23134_, new_n23135_, new_n23136_,
    new_n23137_, new_n23138_, new_n23139_, new_n23140_, new_n23141_,
    new_n23142_, new_n23143_, new_n23144_, new_n23145_, new_n23146_,
    new_n23147_, new_n23148_, new_n23149_, new_n23150_, new_n23151_,
    new_n23152_, new_n23153_, new_n23154_, new_n23155_, new_n23156_,
    new_n23157_, new_n23158_, new_n23159_, new_n23160_, new_n23161_,
    new_n23162_, new_n23163_, new_n23164_, new_n23165_, new_n23166_,
    new_n23167_, new_n23168_, new_n23169_, new_n23170_, new_n23171_,
    new_n23172_, new_n23173_, new_n23174_, new_n23175_, new_n23176_,
    new_n23177_, new_n23178_, new_n23179_, new_n23180_, new_n23181_,
    new_n23182_, new_n23183_, new_n23184_, new_n23185_, new_n23186_,
    new_n23187_, new_n23188_, new_n23189_, new_n23190_, new_n23191_,
    new_n23192_, new_n23193_, new_n23194_, new_n23195_, new_n23196_,
    new_n23197_, new_n23198_, new_n23199_, new_n23200_, new_n23201_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23213_, new_n23214_, new_n23215_, new_n23216_,
    new_n23217_, new_n23218_, new_n23219_, new_n23220_, new_n23221_,
    new_n23222_, new_n23223_, new_n23224_, new_n23225_, new_n23226_,
    new_n23227_, new_n23228_, new_n23229_, new_n23230_, new_n23231_,
    new_n23232_, new_n23233_, new_n23234_, new_n23235_, new_n23236_,
    new_n23237_, new_n23238_, new_n23239_, new_n23240_, new_n23241_,
    new_n23242_, new_n23243_, new_n23244_, new_n23245_, new_n23246_,
    new_n23247_, new_n23248_, new_n23249_, new_n23250_, new_n23251_,
    new_n23252_, new_n23253_, new_n23254_, new_n23255_, new_n23256_,
    new_n23257_, new_n23258_, new_n23259_, new_n23260_, new_n23261_,
    new_n23262_, new_n23263_, new_n23264_, new_n23265_, new_n23266_,
    new_n23267_, new_n23268_, new_n23269_, new_n23270_, new_n23271_,
    new_n23272_, new_n23273_, new_n23274_, new_n23275_, new_n23276_,
    new_n23277_, new_n23278_, new_n23279_, new_n23280_, new_n23281_,
    new_n23282_, new_n23283_, new_n23284_, new_n23285_, new_n23286_,
    new_n23287_, new_n23288_, new_n23289_, new_n23290_, new_n23291_,
    new_n23292_, new_n23293_, new_n23294_, new_n23295_, new_n23296_,
    new_n23297_, new_n23298_, new_n23299_, new_n23300_, new_n23301_,
    new_n23302_, new_n23303_, new_n23304_, new_n23305_, new_n23306_,
    new_n23307_, new_n23308_, new_n23309_, new_n23310_, new_n23311_,
    new_n23312_, new_n23313_, new_n23314_, new_n23315_, new_n23316_,
    new_n23317_, new_n23318_, new_n23319_, new_n23320_, new_n23321_,
    new_n23322_, new_n23323_, new_n23324_, new_n23325_, new_n23326_,
    new_n23327_, new_n23328_, new_n23329_, new_n23330_, new_n23331_,
    new_n23332_, new_n23333_, new_n23334_, new_n23335_, new_n23336_,
    new_n23337_, new_n23338_, new_n23339_, new_n23340_, new_n23341_,
    new_n23342_, new_n23343_, new_n23344_, new_n23346_, new_n23347_,
    new_n23348_, new_n23349_, new_n23350_, new_n23351_, new_n23352_,
    new_n23353_, new_n23354_, new_n23355_, new_n23356_, new_n23357_,
    new_n23358_, new_n23359_, new_n23360_, new_n23361_, new_n23362_,
    new_n23363_, new_n23364_, new_n23365_, new_n23366_, new_n23367_,
    new_n23368_, new_n23369_, new_n23370_, new_n23371_, new_n23372_,
    new_n23373_, new_n23374_, new_n23375_, new_n23376_, new_n23377_,
    new_n23378_, new_n23379_, new_n23380_, new_n23381_, new_n23382_,
    new_n23383_, new_n23384_, new_n23385_, new_n23386_, new_n23387_,
    new_n23389_, new_n23390_, new_n23391_, new_n23392_, new_n23393_,
    new_n23394_, new_n23395_, new_n23396_, new_n23397_, new_n23398_,
    new_n23399_, new_n23400_, new_n23401_, new_n23402_, new_n23403_,
    new_n23404_, new_n23405_, new_n23406_, new_n23407_, new_n23408_,
    new_n23409_, new_n23410_, new_n23411_, new_n23413_, new_n23414_,
    new_n23415_, new_n23416_, new_n23417_, new_n23418_, new_n23419_,
    new_n23420_, new_n23421_, new_n23422_, new_n23423_, new_n23424_,
    new_n23426_, new_n23427_, new_n23428_, new_n23429_, new_n23430_,
    new_n23431_, new_n23433_, new_n23434_, new_n23435_, new_n23438_,
    new_n23439_, new_n23440_, new_n23441_, new_n23442_, new_n23443_,
    new_n23444_, new_n23445_, new_n23446_, new_n23447_, new_n23448_,
    new_n23449_, new_n23450_, new_n23451_, new_n23452_, new_n23453_,
    new_n23454_, new_n23455_, new_n23456_, new_n23457_, new_n23458_,
    new_n23459_, new_n23460_, new_n23461_, new_n23462_, new_n23463_,
    new_n23464_, new_n23465_, new_n23466_, new_n23467_, new_n23468_,
    new_n23469_, new_n23470_, new_n23471_, new_n23472_, new_n23473_,
    new_n23474_, new_n23475_, new_n23476_, new_n23477_, new_n23478_,
    new_n23479_, new_n23480_, new_n23481_, new_n23482_, new_n23483_,
    new_n23484_, new_n23485_, new_n23486_, new_n23487_, new_n23488_,
    new_n23489_, new_n23490_, new_n23491_, new_n23492_, new_n23493_,
    new_n23494_, new_n23495_, new_n23496_, new_n23497_, new_n23498_,
    new_n23499_, new_n23500_, new_n23501_, new_n23502_, new_n23503_,
    new_n23504_, new_n23505_, new_n23506_, new_n23507_, new_n23508_,
    new_n23509_, new_n23510_, new_n23511_, new_n23512_, new_n23513_,
    new_n23514_, new_n23515_, new_n23516_, new_n23517_, new_n23518_,
    new_n23519_, new_n23520_, new_n23521_, new_n23522_, new_n23523_,
    new_n23524_, new_n23525_, new_n23526_, new_n23527_, new_n23528_,
    new_n23529_, new_n23530_, new_n23531_, new_n23532_, new_n23533_,
    new_n23534_, new_n23535_, new_n23536_, new_n23537_, new_n23538_,
    new_n23539_, new_n23540_, new_n23541_, new_n23542_, new_n23543_,
    new_n23544_, new_n23545_, new_n23546_, new_n23547_, new_n23548_,
    new_n23549_, new_n23550_, new_n23551_, new_n23552_, new_n23553_,
    new_n23554_, new_n23555_, new_n23556_, new_n23557_, new_n23558_,
    new_n23559_, new_n23560_, new_n23561_, new_n23562_, new_n23563_,
    new_n23564_, new_n23565_, new_n23566_, new_n23567_, new_n23568_,
    new_n23569_, new_n23570_, new_n23571_, new_n23572_, new_n23573_,
    new_n23574_, new_n23575_, new_n23576_, new_n23577_, new_n23578_,
    new_n23579_, new_n23580_, new_n23581_, new_n23582_, new_n23583_,
    new_n23584_, new_n23585_, new_n23586_, new_n23587_, new_n23588_,
    new_n23589_, new_n23590_, new_n23591_, new_n23592_, new_n23593_,
    new_n23594_, new_n23595_, new_n23596_, new_n23597_, new_n23598_,
    new_n23599_, new_n23600_, new_n23601_, new_n23602_, new_n23603_,
    new_n23604_, new_n23605_, new_n23606_, new_n23607_, new_n23608_,
    new_n23609_, new_n23610_, new_n23611_, new_n23612_, new_n23613_,
    new_n23614_, new_n23615_, new_n23616_, new_n23617_, new_n23618_,
    new_n23619_, new_n23620_, new_n23621_, new_n23622_, new_n23623_,
    new_n23624_, new_n23625_, new_n23626_, new_n23627_, new_n23628_,
    new_n23629_, new_n23630_, new_n23631_, new_n23632_, new_n23633_,
    new_n23634_, new_n23635_, new_n23636_, new_n23637_, new_n23638_,
    new_n23639_, new_n23640_, new_n23641_, new_n23642_, new_n23643_,
    new_n23644_, new_n23645_, new_n23646_, new_n23647_, new_n23648_,
    new_n23649_, new_n23650_, new_n23651_, new_n23652_, new_n23653_,
    new_n23654_, new_n23655_, new_n23656_, new_n23657_, new_n23658_,
    new_n23659_, new_n23660_, new_n23661_, new_n23662_, new_n23663_,
    new_n23664_, new_n23665_, new_n23666_, new_n23667_, new_n23668_,
    new_n23669_, new_n23670_, new_n23671_, new_n23672_, new_n23673_,
    new_n23674_, new_n23675_, new_n23676_, new_n23677_, new_n23678_,
    new_n23679_, new_n23680_, new_n23681_, new_n23682_, new_n23683_,
    new_n23684_, new_n23685_, new_n23686_, new_n23687_, new_n23688_,
    new_n23689_, new_n23690_, new_n23691_, new_n23692_, new_n23693_,
    new_n23694_, new_n23695_, new_n23696_, new_n23697_, new_n23698_,
    new_n23699_, new_n23700_, new_n23701_, new_n23702_, new_n23703_,
    new_n23704_, new_n23705_, new_n23706_, new_n23707_, new_n23708_,
    new_n23709_, new_n23710_, new_n23711_, new_n23712_, new_n23713_,
    new_n23714_, new_n23715_, new_n23716_, new_n23717_, new_n23718_,
    new_n23719_, new_n23720_, new_n23721_, new_n23722_, new_n23723_,
    new_n23724_, new_n23725_, new_n23726_, new_n23727_, new_n23728_,
    new_n23729_, new_n23730_, new_n23731_, new_n23732_, new_n23733_,
    new_n23734_, new_n23735_, new_n23736_, new_n23737_, new_n23738_,
    new_n23739_, new_n23740_, new_n23741_, new_n23742_, new_n23743_,
    new_n23744_, new_n23745_, new_n23746_, new_n23747_, new_n23748_,
    new_n23749_, new_n23750_, new_n23751_, new_n23752_, new_n23753_,
    new_n23754_, new_n23755_, new_n23756_, new_n23757_, new_n23758_,
    new_n23759_, new_n23760_, new_n23761_, new_n23762_, new_n23763_,
    new_n23764_, new_n23765_, new_n23766_, new_n23767_, new_n23768_,
    new_n23769_, new_n23770_, new_n23771_, new_n23772_, new_n23773_,
    new_n23774_, new_n23775_, new_n23776_, new_n23777_, new_n23778_,
    new_n23779_, new_n23780_, new_n23781_, new_n23782_, new_n23783_,
    new_n23784_, new_n23785_, new_n23786_, new_n23787_, new_n23788_,
    new_n23789_, new_n23790_, new_n23791_, new_n23792_, new_n23793_,
    new_n23794_, new_n23795_, new_n23796_, new_n23797_, new_n23798_,
    new_n23799_, new_n23800_, new_n23801_, new_n23802_, new_n23803_,
    new_n23804_, new_n23805_, new_n23806_, new_n23807_, new_n23808_,
    new_n23809_, new_n23810_, new_n23811_, new_n23812_, new_n23813_,
    new_n23814_, new_n23815_, new_n23816_, new_n23817_, new_n23818_,
    new_n23819_, new_n23820_, new_n23821_, new_n23822_, new_n23823_,
    new_n23824_, new_n23825_, new_n23826_, new_n23827_, new_n23828_,
    new_n23829_, new_n23830_, new_n23831_, new_n23832_, new_n23833_,
    new_n23834_, new_n23835_, new_n23836_, new_n23837_, new_n23838_,
    new_n23839_, new_n23840_, new_n23841_, new_n23842_, new_n23843_,
    new_n23844_, new_n23845_, new_n23846_, new_n23847_, new_n23848_,
    new_n23849_, new_n23850_, new_n23851_, new_n23852_, new_n23853_,
    new_n23854_, new_n23855_, new_n23856_, new_n23857_, new_n23858_,
    new_n23859_, new_n23860_, new_n23861_, new_n23862_, new_n23863_,
    new_n23864_, new_n23865_, new_n23866_, new_n23867_, new_n23868_,
    new_n23869_, new_n23870_, new_n23871_, new_n23872_, new_n23873_,
    new_n23874_, new_n23875_, new_n23876_, new_n23877_, new_n23878_,
    new_n23879_, new_n23880_, new_n23881_, new_n23882_, new_n23883_,
    new_n23884_, new_n23885_, new_n23886_, new_n23887_, new_n23888_,
    new_n23889_, new_n23890_, new_n23891_, new_n23892_, new_n23893_,
    new_n23894_, new_n23895_, new_n23896_, new_n23897_, new_n23898_,
    new_n23899_, new_n23900_, new_n23901_, new_n23902_, new_n23903_,
    new_n23904_, new_n23905_, new_n23906_, new_n23907_, new_n23908_,
    new_n23909_, new_n23910_, new_n23911_, new_n23912_, new_n23913_,
    new_n23914_, new_n23915_, new_n23916_, new_n23917_, new_n23918_,
    new_n23919_, new_n23920_, new_n23921_, new_n23922_, new_n23923_,
    new_n23924_, new_n23925_, new_n23926_, new_n23927_, new_n23928_,
    new_n23929_, new_n23930_, new_n23931_, new_n23932_, new_n23933_,
    new_n23934_, new_n23935_, new_n23936_, new_n23937_, new_n23938_,
    new_n23939_, new_n23940_, new_n23941_, new_n23942_, new_n23943_,
    new_n23944_, new_n23945_, new_n23946_, new_n23947_, new_n23948_,
    new_n23949_, new_n23950_, new_n23951_, new_n23952_, new_n23953_,
    new_n23954_, new_n23955_, new_n23956_, new_n23957_, new_n23958_,
    new_n23959_, new_n23960_, new_n23961_, new_n23962_, new_n23963_,
    new_n23964_, new_n23965_, new_n23966_, new_n23967_, new_n23968_,
    new_n23969_, new_n23970_, new_n23971_, new_n23972_, new_n23973_,
    new_n23974_, new_n23975_, new_n23976_, new_n23977_, new_n23978_,
    new_n23979_, new_n23980_, new_n23981_, new_n23982_, new_n23983_,
    new_n23984_, new_n23985_, new_n23986_, new_n23987_, new_n23988_,
    new_n23989_, new_n23990_, new_n23991_, new_n23993_, new_n23994_,
    new_n23995_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24004_, new_n24005_, new_n24006_,
    new_n24007_, new_n24008_, new_n24009_, new_n24010_, new_n24011_,
    new_n24012_, new_n24013_, new_n24014_, new_n24015_, new_n24016_,
    new_n24017_, new_n24018_, new_n24019_, new_n24020_, new_n24021_,
    new_n24022_, new_n24023_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24240_, new_n24241_,
    new_n24242_, new_n24243_, new_n24244_, new_n24245_, new_n24246_,
    new_n24247_, new_n24248_, new_n24249_, new_n24250_, new_n24251_,
    new_n24252_, new_n24253_, new_n24254_, new_n24255_, new_n24256_,
    new_n24257_, new_n24258_, new_n24259_, new_n24260_, new_n24261_,
    new_n24262_, new_n24263_, new_n24264_, new_n24265_, new_n24266_,
    new_n24267_, new_n24268_, new_n24269_, new_n24270_, new_n24271_,
    new_n24272_, new_n24273_, new_n24274_, new_n24275_, new_n24276_,
    new_n24277_, new_n24278_, new_n24279_, new_n24280_, new_n24281_,
    new_n24282_, new_n24283_, new_n24284_, new_n24285_, new_n24286_,
    new_n24287_, new_n24288_, new_n24289_, new_n24290_, new_n24291_,
    new_n24292_, new_n24293_, new_n24294_, new_n24295_, new_n24296_,
    new_n24297_, new_n24298_, new_n24299_, new_n24300_, new_n24301_,
    new_n24302_, new_n24303_, new_n24304_, new_n24305_, new_n24306_,
    new_n24307_, new_n24308_, new_n24309_, new_n24310_, new_n24311_,
    new_n24312_, new_n24313_, new_n24314_, new_n24315_, new_n24316_,
    new_n24317_, new_n24318_, new_n24319_, new_n24320_, new_n24321_,
    new_n24322_, new_n24323_, new_n24324_, new_n24325_, new_n24326_,
    new_n24327_, new_n24328_, new_n24329_, new_n24330_, new_n24331_,
    new_n24332_, new_n24333_, new_n24334_, new_n24335_, new_n24336_,
    new_n24337_, new_n24338_, new_n24339_, new_n24340_, new_n24341_,
    new_n24342_, new_n24343_, new_n24344_, new_n24345_, new_n24346_,
    new_n24347_, new_n24348_, new_n24349_, new_n24350_, new_n24351_,
    new_n24352_, new_n24353_, new_n24354_, new_n24355_, new_n24356_,
    new_n24357_, new_n24358_, new_n24359_, new_n24360_, new_n24361_,
    new_n24362_, new_n24363_, new_n24364_, new_n24365_, new_n24366_,
    new_n24367_, new_n24368_, new_n24369_, new_n24370_, new_n24371_,
    new_n24372_, new_n24373_, new_n24374_, new_n24375_, new_n24376_,
    new_n24377_, new_n24378_, new_n24379_, new_n24380_, new_n24381_,
    new_n24382_, new_n24383_, new_n24384_, new_n24385_, new_n24386_,
    new_n24387_, new_n24388_, new_n24389_, new_n24390_, new_n24391_,
    new_n24392_, new_n24393_, new_n24394_, new_n24395_, new_n24396_,
    new_n24397_, new_n24398_, new_n24399_, new_n24400_, new_n24401_,
    new_n24402_, new_n24403_, new_n24404_, new_n24405_, new_n24406_,
    new_n24407_, new_n24408_, new_n24409_, new_n24410_, new_n24411_,
    new_n24412_, new_n24413_, new_n24414_, new_n24415_, new_n24416_,
    new_n24417_, new_n24418_, new_n24419_, new_n24420_, new_n24421_,
    new_n24422_, new_n24423_, new_n24424_, new_n24425_, new_n24426_,
    new_n24427_, new_n24428_, new_n24429_, new_n24430_, new_n24431_,
    new_n24432_, new_n24433_, new_n24434_, new_n24435_, new_n24436_,
    new_n24437_, new_n24438_, new_n24439_, new_n24440_, new_n24441_,
    new_n24442_, new_n24443_, new_n24444_, new_n24445_, new_n24446_,
    new_n24447_, new_n24448_, new_n24449_, new_n24450_, new_n24451_,
    new_n24452_, new_n24453_, new_n24454_, new_n24455_, new_n24456_,
    new_n24457_, new_n24458_, new_n24459_, new_n24460_, new_n24461_,
    new_n24462_, new_n24463_, new_n24464_, new_n24465_, new_n24466_,
    new_n24467_, new_n24468_, new_n24469_, new_n24470_, new_n24471_,
    new_n24472_, new_n24473_, new_n24474_, new_n24475_, new_n24476_,
    new_n24477_, new_n24478_, new_n24479_, new_n24480_, new_n24481_,
    new_n24482_, new_n24483_, new_n24484_, new_n24485_, new_n24486_,
    new_n24487_, new_n24488_, new_n24489_, new_n24490_, new_n24491_,
    new_n24492_, new_n24493_, new_n24494_, new_n24495_, new_n24496_,
    new_n24497_, new_n24498_, new_n24499_, new_n24500_, new_n24501_,
    new_n24502_, new_n24503_, new_n24504_, new_n24505_, new_n24506_,
    new_n24507_, new_n24508_, new_n24509_, new_n24510_, new_n24511_,
    new_n24512_, new_n24513_, new_n24514_, new_n24515_, new_n24516_,
    new_n24517_, new_n24518_, new_n24519_, new_n24520_, new_n24521_,
    new_n24522_, new_n24523_, new_n24524_, new_n24525_, new_n24526_,
    new_n24527_, new_n24528_, new_n24529_, new_n24530_, new_n24531_,
    new_n24532_, new_n24533_, new_n24534_, new_n24535_, new_n24536_,
    new_n24537_, new_n24538_, new_n24539_, new_n24540_, new_n24541_,
    new_n24542_, new_n24543_, new_n24544_, new_n24545_, new_n24546_,
    new_n24547_, new_n24548_, new_n24549_, new_n24550_, new_n24551_,
    new_n24552_, new_n24553_, new_n24554_, new_n24555_, new_n24556_,
    new_n24557_, new_n24558_, new_n24559_, new_n24560_, new_n24561_,
    new_n24562_, new_n24563_, new_n24564_, new_n24565_, new_n24566_,
    new_n24567_, new_n24568_, new_n24569_, new_n24570_, new_n24571_,
    new_n24572_, new_n24573_, new_n24574_, new_n24575_, new_n24576_,
    new_n24578_, new_n24579_, new_n24580_, new_n24581_, new_n24582_,
    new_n24583_, new_n24584_, new_n24585_, new_n24586_, new_n24587_,
    new_n24588_, new_n24589_, new_n24590_, new_n24591_, new_n24592_,
    new_n24593_, new_n24594_, new_n24595_, new_n24596_, new_n24597_,
    new_n24598_, new_n24599_, new_n24600_, new_n24601_, new_n24602_,
    new_n24603_, new_n24604_, new_n24605_, new_n24606_, new_n24607_,
    new_n24608_, new_n24609_, new_n24610_, new_n24611_, new_n24612_,
    new_n24613_, new_n24614_, new_n24615_, new_n24616_, new_n24617_,
    new_n24618_, new_n24619_, new_n24620_, new_n24621_, new_n24622_,
    new_n24623_, new_n24624_, new_n24625_, new_n24626_, new_n24627_,
    new_n24628_, new_n24629_, new_n24630_, new_n24631_, new_n24633_,
    new_n24634_, new_n24635_, new_n24636_, new_n24637_, new_n24638_,
    new_n24639_, new_n24640_, new_n24641_, new_n24642_, new_n24643_,
    new_n24644_, new_n24645_, new_n24646_, new_n24647_, new_n24648_,
    new_n24649_, new_n24650_, new_n24651_, new_n24652_, new_n24653_,
    new_n24654_, new_n24655_, new_n24656_, new_n24657_, new_n24658_,
    new_n24659_, new_n24660_, new_n24661_, new_n24662_, new_n24663_,
    new_n24664_, new_n24666_, new_n24667_, new_n24668_, new_n24669_,
    new_n24670_, new_n24671_, new_n24672_, new_n24673_, new_n24674_,
    new_n24675_, new_n24676_, new_n24677_, new_n24678_, new_n24679_,
    new_n24680_, new_n24681_, new_n24682_, new_n24683_, new_n24685_,
    new_n24686_, new_n24687_, new_n24688_, new_n24689_, new_n24690_,
    new_n24691_, new_n24692_, new_n24693_, new_n24695_, new_n24696_,
    new_n24697_, new_n24698_, new_n24701_, new_n24702_, new_n24703_,
    new_n24704_, new_n24705_, new_n24706_, new_n24707_, new_n24708_,
    new_n24709_, new_n24710_, new_n24711_, new_n24712_, new_n24713_,
    new_n24714_, new_n24715_, new_n24716_, new_n24717_, new_n24718_,
    new_n24719_, new_n24720_, new_n24721_, new_n24722_, new_n24723_,
    new_n24724_, new_n24725_, new_n24726_, new_n24727_, new_n24728_,
    new_n24729_, new_n24730_, new_n24731_, new_n24732_, new_n24733_,
    new_n24734_, new_n24735_, new_n24736_, new_n24737_, new_n24738_,
    new_n24739_, new_n24740_, new_n24741_, new_n24742_, new_n24743_,
    new_n24744_, new_n24745_, new_n24746_, new_n24747_, new_n24748_,
    new_n24749_, new_n24750_, new_n24751_, new_n24752_, new_n24753_,
    new_n24754_, new_n24755_, new_n24756_, new_n24757_, new_n24758_,
    new_n24759_, new_n24760_, new_n24761_, new_n24762_, new_n24763_,
    new_n24764_, new_n24765_, new_n24766_, new_n24767_, new_n24768_,
    new_n24769_, new_n24770_, new_n24771_, new_n24772_, new_n24773_,
    new_n24774_, new_n24775_, new_n24776_, new_n24777_, new_n24778_,
    new_n24779_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24799_, new_n24800_, new_n24801_, new_n24802_, new_n24803_,
    new_n24804_, new_n24805_, new_n24806_, new_n24807_, new_n24808_,
    new_n24809_, new_n24810_, new_n24811_, new_n24812_, new_n24813_,
    new_n24814_, new_n24815_, new_n24816_, new_n24817_, new_n24818_,
    new_n24819_, new_n24820_, new_n24821_, new_n24822_, new_n24823_,
    new_n24824_, new_n24825_, new_n24826_, new_n24827_, new_n24828_,
    new_n24829_, new_n24830_, new_n24831_, new_n24832_, new_n24833_,
    new_n24834_, new_n24835_, new_n24836_, new_n24837_, new_n24838_,
    new_n24839_, new_n24840_, new_n24841_, new_n24842_, new_n24843_,
    new_n24844_, new_n24845_, new_n24846_, new_n24847_, new_n24848_,
    new_n24849_, new_n24850_, new_n24851_, new_n24852_, new_n24853_,
    new_n24854_, new_n24855_, new_n24856_, new_n24857_, new_n24858_,
    new_n24859_, new_n24860_, new_n24861_, new_n24862_, new_n24863_,
    new_n24864_, new_n24865_, new_n24866_, new_n24867_, new_n24868_,
    new_n24869_, new_n24870_, new_n24871_, new_n24872_, new_n24873_,
    new_n24874_, new_n24875_, new_n24876_, new_n24877_, new_n24878_,
    new_n24879_, new_n24880_, new_n24881_, new_n24882_, new_n24883_,
    new_n24884_, new_n24885_, new_n24886_, new_n24887_, new_n24888_,
    new_n24889_, new_n24890_, new_n24891_, new_n24892_, new_n24893_,
    new_n24894_, new_n24895_, new_n24896_, new_n24897_, new_n24898_,
    new_n24899_, new_n24900_, new_n24901_, new_n24902_, new_n24903_,
    new_n24904_, new_n24905_, new_n24906_, new_n24907_, new_n24908_,
    new_n24909_, new_n24910_, new_n24911_, new_n24912_, new_n24913_,
    new_n24914_, new_n24915_, new_n24916_, new_n24917_, new_n24918_,
    new_n24919_, new_n24920_, new_n24921_, new_n24922_, new_n24923_,
    new_n24924_, new_n24925_, new_n24926_, new_n24927_, new_n24928_,
    new_n24930_, new_n24931_, new_n24932_, new_n24933_, new_n24934_,
    new_n24938_, new_n24939_, new_n24940_, new_n24943_, new_n24944_,
    new_n24945_, new_n24946_, new_n24947_, new_n24948_, new_n24949_,
    new_n24950_, new_n24951_, new_n24952_, new_n24953_, new_n24954_,
    new_n24955_, new_n24956_, new_n24957_, new_n24958_, new_n24959_,
    new_n24960_, new_n24961_, new_n24962_, new_n24963_, new_n24964_,
    new_n24965_, new_n24966_, new_n24967_, new_n24968_, new_n24969_,
    new_n24970_, new_n24971_, new_n24972_, new_n24973_, new_n24974_,
    new_n24975_, new_n24976_, new_n24977_, new_n24978_, new_n24979_,
    new_n24980_, new_n24981_, new_n24982_, new_n24983_, new_n24984_,
    new_n24985_, new_n24986_, new_n24987_, new_n24988_, new_n24989_,
    new_n24990_, new_n24991_, new_n24992_, new_n24993_, new_n24994_,
    new_n24995_, new_n24996_, new_n24997_, new_n24998_, new_n24999_,
    new_n25000_, new_n25001_, new_n25002_, new_n25003_, new_n25004_,
    new_n25005_, new_n25006_, new_n25007_, new_n25008_, new_n25009_,
    new_n25010_, new_n25011_, new_n25012_, new_n25013_, new_n25014_,
    new_n25015_, new_n25016_, new_n25017_, new_n25018_, new_n25019_,
    new_n25020_, new_n25021_, new_n25022_, new_n25023_, new_n25024_,
    new_n25025_, new_n25026_, new_n25027_, new_n25028_, new_n25029_,
    new_n25030_, new_n25031_, new_n25032_, new_n25033_, new_n25034_,
    new_n25035_, new_n25036_, new_n25037_, new_n25038_, new_n25039_,
    new_n25040_, new_n25041_, new_n25042_, new_n25043_, new_n25044_,
    new_n25045_, new_n25046_, new_n25047_, new_n25048_, new_n25049_,
    new_n25050_, new_n25051_, new_n25052_, new_n25053_, new_n25054_,
    new_n25055_, new_n25056_, new_n25057_, new_n25058_, new_n25059_,
    new_n25060_, new_n25061_, new_n25062_, new_n25063_, new_n25064_,
    new_n25065_, new_n25066_, new_n25067_, new_n25068_, new_n25069_,
    new_n25070_, new_n25071_, new_n25072_, new_n25073_, new_n25074_,
    new_n25075_, new_n25076_, new_n25077_, new_n25078_, new_n25079_,
    new_n25080_, new_n25081_, new_n25082_, new_n25083_, new_n25084_,
    new_n25085_, new_n25086_, new_n25087_, new_n25088_, new_n25089_,
    new_n25090_, new_n25091_, new_n25092_, new_n25093_, new_n25094_,
    new_n25095_, new_n25096_, new_n25097_, new_n25098_, new_n25099_,
    new_n25100_, new_n25101_, new_n25102_, new_n25103_, new_n25104_,
    new_n25105_, new_n25106_, new_n25107_, new_n25108_, new_n25109_,
    new_n25110_, new_n25111_, new_n25112_, new_n25113_, new_n25114_,
    new_n25115_, new_n25116_, new_n25117_, new_n25118_, new_n25119_,
    new_n25120_, new_n25121_, new_n25122_, new_n25123_, new_n25124_,
    new_n25125_, new_n25126_, new_n25127_, new_n25128_, new_n25129_,
    new_n25130_, new_n25132_, new_n25133_, new_n25134_, new_n25135_,
    new_n25136_, new_n25137_, new_n25140_, new_n25141_, new_n25142_,
    new_n25143_, new_n25144_, new_n25145_, new_n25146_, new_n25147_,
    new_n25148_, new_n25149_, new_n25150_, new_n25151_, new_n25152_,
    new_n25153_, new_n25154_, new_n25155_, new_n25156_, new_n25157_,
    new_n25158_, new_n25159_, new_n25160_, new_n25161_, new_n25162_,
    new_n25163_, new_n25164_, new_n25165_, new_n25166_, new_n25167_,
    new_n25168_, new_n25169_, new_n25170_, new_n25171_, new_n25172_,
    new_n25173_, new_n25174_, new_n25175_, new_n25176_, new_n25177_,
    new_n25178_, new_n25179_, new_n25180_, new_n25181_, new_n25182_,
    new_n25183_, new_n25184_, new_n25185_, new_n25186_, new_n25187_,
    new_n25188_, new_n25189_, new_n25190_, new_n25191_, new_n25192_,
    new_n25193_, new_n25194_, new_n25195_, new_n25196_, new_n25197_,
    new_n25198_, new_n25199_, new_n25200_, new_n25201_, new_n25202_,
    new_n25203_, new_n25204_, new_n25205_, new_n25206_, new_n25207_,
    new_n25208_, new_n25209_, new_n25210_, new_n25211_, new_n25212_,
    new_n25213_, new_n25214_, new_n25215_, new_n25218_, new_n25219_,
    new_n25220_, new_n25221_, new_n25222_, new_n25223_, new_n25224_,
    new_n25225_, new_n25226_, new_n25227_, new_n25228_, new_n25229_,
    new_n25230_, new_n25231_, new_n25232_, new_n25233_, new_n25234_,
    new_n25235_, new_n25236_, new_n25237_, new_n25238_, new_n25239_,
    new_n25240_, new_n25241_, new_n25242_, new_n25243_, new_n25244_,
    new_n25245_, new_n25246_, new_n25247_, new_n25248_, new_n25249_,
    new_n25250_, new_n25251_, new_n25252_, new_n25253_, new_n25254_,
    new_n25255_, new_n25256_, new_n25257_, new_n25258_, new_n25259_,
    new_n25260_, new_n25261_, new_n25262_, new_n25263_, new_n25264_,
    new_n25265_, new_n25266_, new_n25267_, new_n25268_, new_n25269_,
    new_n25270_, new_n25271_, new_n25272_, new_n25273_, new_n25274_,
    new_n25275_, new_n25276_, new_n25277_, new_n25278_, new_n25279_,
    new_n25280_, new_n25281_, new_n25282_, new_n25283_, new_n25284_,
    new_n25285_, new_n25286_, new_n25287_, new_n25288_, new_n25289_,
    new_n25290_, new_n25291_, new_n25292_, new_n25293_, new_n25294_,
    new_n25295_, new_n25296_, new_n25297_, new_n25298_, new_n25299_,
    new_n25300_, new_n25301_, new_n25302_, new_n25303_, new_n25304_,
    new_n25305_, new_n25306_, new_n25307_, new_n25308_, new_n25309_,
    new_n25311_, new_n25312_, new_n25313_, new_n25314_, new_n25315_,
    new_n25316_, new_n25319_, new_n25320_, new_n25321_, new_n25322_,
    new_n25323_, new_n25324_, new_n25325_, new_n25326_, new_n25327_,
    new_n25328_, new_n25329_, new_n25330_, new_n25331_, new_n25332_,
    new_n25333_, new_n25334_, new_n25335_, new_n25336_, new_n25337_,
    new_n25338_, new_n25339_, new_n25340_, new_n25341_, new_n25342_,
    new_n25343_, new_n25344_, new_n25345_, new_n25346_, new_n25347_,
    new_n25348_, new_n25349_, new_n25350_, new_n25351_, new_n25352_,
    new_n25353_, new_n25354_, new_n25355_, new_n25356_, new_n25357_,
    new_n25358_, new_n25359_, new_n25360_, new_n25361_, new_n25362_,
    new_n25363_, new_n25364_, new_n25365_, new_n25366_, new_n25367_,
    new_n25368_, new_n25369_, new_n25370_, new_n25371_, new_n25372_,
    new_n25373_, new_n25374_, new_n25375_, new_n25376_, new_n25377_,
    new_n25378_, new_n25379_, new_n25380_, new_n25381_, new_n25382_,
    new_n25383_, new_n25384_, new_n25385_, new_n25386_, new_n25387_,
    new_n25388_, new_n25389_, new_n25390_, new_n25391_, new_n25392_,
    new_n25393_, new_n25394_, new_n25395_, new_n25396_, new_n25397_,
    new_n25398_, new_n25399_, new_n25400_, new_n25401_, new_n25402_,
    new_n25403_, new_n25404_, new_n25405_, new_n25406_, new_n25407_,
    new_n25408_, new_n25409_, new_n25410_, new_n25411_, new_n25412_,
    new_n25413_, new_n25414_, new_n25415_, new_n25416_, new_n25417_,
    new_n25418_, new_n25419_, new_n25420_, new_n25421_, new_n25422_,
    new_n25424_, new_n25425_, new_n25426_, new_n25427_, new_n25428_,
    new_n25429_, new_n25430_, new_n25431_, new_n25432_, new_n25433_,
    new_n25434_, new_n25435_, new_n25436_, new_n25437_, new_n25438_,
    new_n25439_, new_n25440_, new_n25441_, new_n25442_, new_n25443_,
    new_n25444_, new_n25445_, new_n25446_, new_n25447_, new_n25448_,
    new_n25449_, new_n25450_, new_n25451_, new_n25452_, new_n25453_,
    new_n25454_, new_n25455_, new_n25456_, new_n25457_, new_n25458_,
    new_n25459_, new_n25460_, new_n25461_, new_n25462_, new_n25463_,
    new_n25464_, new_n25465_, new_n25466_, new_n25467_, new_n25468_,
    new_n25469_, new_n25470_, new_n25471_, new_n25472_, new_n25473_,
    new_n25474_, new_n25475_, new_n25477_, new_n25478_, new_n25479_,
    new_n25480_, new_n25481_, new_n25482_, new_n25483_, new_n25484_,
    new_n25485_, new_n25486_, new_n25487_, new_n25488_, new_n25489_,
    new_n25490_, new_n25491_, new_n25492_, new_n25493_, new_n25494_,
    new_n25495_, new_n25496_, new_n25497_, new_n25498_, new_n25499_,
    new_n25500_, new_n25501_, new_n25502_, new_n25503_, new_n25504_,
    new_n25505_, new_n25507_, new_n25508_, new_n25509_, new_n25510_,
    new_n25511_, new_n25512_, new_n25513_, new_n25514_, new_n25515_,
    new_n25516_, new_n25517_, new_n25518_, new_n25519_, new_n25520_,
    new_n25521_, new_n25523_, new_n25524_, new_n25525_, new_n25526_,
    new_n25527_, new_n25528_, new_n25529_, new_n25530_, new_n25532_,
    new_n25533_, new_n25534_, new_n25535_, new_n25538_, new_n25539_,
    new_n25540_, new_n25541_, new_n25542_, new_n25543_, new_n25544_,
    new_n25545_, new_n25546_, new_n25547_, new_n25548_, new_n25549_,
    new_n25550_, new_n25551_, new_n25552_, new_n25553_, new_n25554_,
    new_n25555_, new_n25556_, new_n25557_, new_n25558_, new_n25559_,
    new_n25560_, new_n25561_, new_n25562_, new_n25563_, new_n25564_,
    new_n25565_, new_n25566_, new_n25567_, new_n25568_, new_n25569_,
    new_n25570_, new_n25571_, new_n25572_, new_n25573_, new_n25574_,
    new_n25575_, new_n25576_, new_n25577_, new_n25578_, new_n25579_,
    new_n25580_, new_n25581_, new_n25582_, new_n25583_, new_n25584_,
    new_n25585_, new_n25586_, new_n25587_, new_n25588_, new_n25589_,
    new_n25590_, new_n25591_, new_n25592_, new_n25593_, new_n25594_,
    new_n25595_, new_n25596_, new_n25597_, new_n25598_, new_n25599_,
    new_n25600_, new_n25601_, new_n25602_, new_n25603_, new_n25604_,
    new_n25605_, new_n25606_, new_n25607_, new_n25608_, new_n25609_,
    new_n25610_, new_n25611_, new_n25612_, new_n25613_, new_n25614_,
    new_n25615_, new_n25616_, new_n25617_, new_n25618_, new_n25619_,
    new_n25620_, new_n25621_, new_n25622_, new_n25623_, new_n25624_,
    new_n25625_, new_n25626_, new_n25627_, new_n25628_, new_n25629_,
    new_n25630_, new_n25631_, new_n25632_, new_n25633_, new_n25634_,
    new_n25635_, new_n25636_, new_n25637_, new_n25638_, new_n25639_,
    new_n25640_, new_n25641_, new_n25642_, new_n25643_, new_n25644_,
    new_n25645_, new_n25647_, new_n25648_, new_n25649_, new_n25650_,
    new_n25651_, new_n25652_, new_n25653_, new_n25654_, new_n25655_,
    new_n25656_, new_n25657_, new_n25658_, new_n25659_, new_n25660_,
    new_n25661_, new_n25662_, new_n25663_, new_n25664_, new_n25665_,
    new_n25666_, new_n25667_, new_n25668_, new_n25669_, new_n25670_,
    new_n25671_, new_n25672_, new_n25673_, new_n25674_, new_n25675_,
    new_n25676_, new_n25677_, new_n25678_, new_n25679_, new_n25680_,
    new_n25681_, new_n25682_, new_n25683_, new_n25684_, new_n25685_,
    new_n25686_, new_n25687_, new_n25688_, new_n25689_, new_n25690_,
    new_n25691_, new_n25692_, new_n25693_, new_n25694_, new_n25695_,
    new_n25696_, new_n25697_, new_n25698_, new_n25699_, new_n25700_,
    new_n25701_, new_n25702_, new_n25703_, new_n25704_, new_n25705_,
    new_n25706_, new_n25707_, new_n25708_, new_n25709_, new_n25710_,
    new_n25711_, new_n25712_, new_n25713_, new_n25714_, new_n25715_,
    new_n25716_, new_n25717_, new_n25718_, new_n25719_, new_n25720_,
    new_n25721_, new_n25722_, new_n25723_, new_n25724_, new_n25725_,
    new_n25726_, new_n25727_, new_n25728_, new_n25729_, new_n25730_,
    new_n25731_, new_n25732_, new_n25733_, new_n25734_, new_n25735_,
    new_n25736_, new_n25737_, new_n25738_, new_n25739_, new_n25740_,
    new_n25741_, new_n25742_, new_n25743_, new_n25744_, new_n25745_,
    new_n25746_, new_n25747_, new_n25748_, new_n25749_, new_n25750_,
    new_n25751_, new_n25752_, new_n25753_, new_n25754_, new_n25755_,
    new_n25756_, new_n25757_, new_n25758_, new_n25759_, new_n25760_,
    new_n25761_, new_n25762_, new_n25763_, new_n25764_, new_n25765_,
    new_n25766_, new_n25767_, new_n25768_, new_n25769_, new_n25770_,
    new_n25771_, new_n25772_, new_n25773_, new_n25774_, new_n25775_,
    new_n25776_, new_n25777_, new_n25778_, new_n25779_, new_n25780_,
    new_n25781_, new_n25782_, new_n25783_, new_n25784_, new_n25785_,
    new_n25786_, new_n25787_, new_n25788_, new_n25789_, new_n25790_,
    new_n25791_, new_n25792_, new_n25793_, new_n25794_, new_n25795_,
    new_n25796_, new_n25797_, new_n25798_, new_n25799_, new_n25800_,
    new_n25801_, new_n25802_, new_n25803_, new_n25804_, new_n25805_,
    new_n25806_, new_n25807_, new_n25808_, new_n25809_, new_n25810_,
    new_n25811_, new_n25812_, new_n25813_, new_n25814_, new_n25815_,
    new_n25816_, new_n25817_, new_n25818_, new_n25819_, new_n25820_,
    new_n25821_, new_n25822_, new_n25823_, new_n25824_, new_n25825_,
    new_n25826_, new_n25827_, new_n25828_, new_n25829_, new_n25830_,
    new_n25831_, new_n25832_, new_n25833_, new_n25834_, new_n25835_,
    new_n25836_, new_n25837_, new_n25838_, new_n25839_, new_n25840_,
    new_n25841_, new_n25842_, new_n25843_, new_n25844_, new_n25845_,
    new_n25846_, new_n25847_, new_n25848_, new_n25849_, new_n25850_,
    new_n25851_, new_n25852_, new_n25853_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25879_, new_n25880_,
    new_n25881_, new_n25882_, new_n25883_, new_n25884_, new_n25885_,
    new_n25886_, new_n25887_, new_n25888_, new_n25889_, new_n25890_,
    new_n25891_, new_n25892_, new_n25893_, new_n25894_, new_n25895_,
    new_n25896_, new_n25897_, new_n25898_, new_n25899_, new_n25900_,
    new_n25901_, new_n25902_, new_n25903_, new_n25904_, new_n25905_,
    new_n25906_, new_n25907_, new_n25908_, new_n25909_, new_n25910_,
    new_n25911_, new_n25912_, new_n25913_, new_n25914_, new_n25915_,
    new_n25916_, new_n25917_, new_n25918_, new_n25919_, new_n25920_,
    new_n25921_, new_n25922_, new_n25923_, new_n25924_, new_n25925_,
    new_n25926_, new_n25927_, new_n25928_, new_n25929_, new_n25930_,
    new_n25931_, new_n25932_, new_n25933_, new_n25934_, new_n25935_,
    new_n25936_, new_n25937_, new_n25938_, new_n25939_, new_n25940_,
    new_n25941_, new_n25942_, new_n25943_, new_n25944_, new_n25945_,
    new_n25946_, new_n25947_, new_n25948_, new_n25949_, new_n25950_,
    new_n25951_, new_n25952_, new_n25953_, new_n25954_, new_n25955_,
    new_n25956_, new_n25957_, new_n25958_, new_n25959_, new_n25960_,
    new_n25961_, new_n25962_, new_n25963_, new_n25964_, new_n25965_,
    new_n25966_, new_n25967_, new_n25968_, new_n25969_, new_n25970_,
    new_n25971_, new_n25972_, new_n25973_, new_n25974_, new_n25975_,
    new_n25976_, new_n25977_, new_n25978_, new_n25979_, new_n25980_,
    new_n25981_, new_n25982_, new_n25983_, new_n25984_, new_n25985_,
    new_n25986_, new_n25987_, new_n25988_, new_n25989_, new_n25990_,
    new_n25991_, new_n25992_, new_n25993_, new_n25994_, new_n25995_,
    new_n25996_, new_n25997_, new_n25998_, new_n25999_, new_n26000_,
    new_n26001_, new_n26002_, new_n26003_, new_n26004_, new_n26005_,
    new_n26006_, new_n26007_, new_n26008_, new_n26009_, new_n26010_,
    new_n26011_, new_n26012_, new_n26013_, new_n26014_, new_n26015_,
    new_n26016_, new_n26017_, new_n26018_, new_n26019_, new_n26020_,
    new_n26021_, new_n26022_, new_n26023_, new_n26024_, new_n26025_,
    new_n26026_, new_n26027_, new_n26028_, new_n26029_, new_n26030_,
    new_n26031_, new_n26032_, new_n26033_, new_n26034_, new_n26035_,
    new_n26036_, new_n26037_, new_n26038_, new_n26039_, new_n26040_,
    new_n26041_, new_n26042_, new_n26043_, new_n26044_, new_n26045_,
    new_n26046_, new_n26047_, new_n26048_, new_n26049_, new_n26050_,
    new_n26051_, new_n26052_, new_n26053_, new_n26054_, new_n26055_,
    new_n26056_, new_n26057_, new_n26058_, new_n26059_, new_n26060_,
    new_n26061_, new_n26062_, new_n26063_, new_n26064_, new_n26065_,
    new_n26066_, new_n26067_, new_n26068_, new_n26069_, new_n26070_,
    new_n26071_, new_n26072_, new_n26073_, new_n26074_, new_n26075_,
    new_n26076_, new_n26077_, new_n26078_, new_n26079_, new_n26080_,
    new_n26081_, new_n26082_, new_n26083_, new_n26084_, new_n26085_,
    new_n26086_, new_n26087_, new_n26088_, new_n26089_, new_n26090_,
    new_n26091_, new_n26092_, new_n26093_, new_n26094_, new_n26095_,
    new_n26096_, new_n26097_, new_n26098_, new_n26099_, new_n26100_,
    new_n26101_, new_n26102_, new_n26103_, new_n26104_, new_n26105_,
    new_n26106_, new_n26107_, new_n26108_, new_n26109_, new_n26110_,
    new_n26111_, new_n26112_, new_n26113_, new_n26114_, new_n26115_,
    new_n26116_, new_n26117_, new_n26118_, new_n26119_, new_n26120_,
    new_n26121_, new_n26122_, new_n26125_, new_n26126_, new_n26127_,
    new_n26128_, new_n26129_, new_n26130_, new_n26131_, new_n26132_,
    new_n26133_, new_n26134_, new_n26135_, new_n26136_, new_n26137_,
    new_n26138_, new_n26139_, new_n26140_, new_n26141_, new_n26142_,
    new_n26143_, new_n26144_, new_n26145_, new_n26146_, new_n26147_,
    new_n26148_, new_n26149_, new_n26150_, new_n26151_, new_n26152_,
    new_n26153_, new_n26154_, new_n26155_, new_n26156_, new_n26157_,
    new_n26158_, new_n26159_, new_n26160_, new_n26161_, new_n26162_,
    new_n26163_, new_n26164_, new_n26165_, new_n26166_, new_n26167_,
    new_n26168_, new_n26169_, new_n26170_, new_n26171_, new_n26172_,
    new_n26173_, new_n26174_, new_n26175_, new_n26176_, new_n26177_,
    new_n26178_, new_n26179_, new_n26180_, new_n26181_, new_n26182_,
    new_n26183_, new_n26184_, new_n26185_, new_n26186_, new_n26187_,
    new_n26188_, new_n26189_, new_n26190_, new_n26191_, new_n26192_,
    new_n26193_, new_n26194_, new_n26195_, new_n26196_, new_n26197_,
    new_n26198_, new_n26199_, new_n26200_, new_n26201_, new_n26202_,
    new_n26203_, new_n26204_, new_n26205_, new_n26206_, new_n26207_,
    new_n26208_, new_n26209_, new_n26210_, new_n26211_, new_n26212_,
    new_n26213_, new_n26214_, new_n26215_, new_n26216_, new_n26217_,
    new_n26218_, new_n26219_, new_n26220_, new_n26221_, new_n26222_,
    new_n26223_, new_n26224_, new_n26225_, new_n26226_, new_n26227_,
    new_n26228_, new_n26229_, new_n26230_, new_n26231_, new_n26232_,
    new_n26233_, new_n26234_, new_n26235_, new_n26236_, new_n26237_,
    new_n26238_, new_n26239_, new_n26240_, new_n26241_, new_n26242_,
    new_n26243_, new_n26244_, new_n26245_, new_n26246_, new_n26247_,
    new_n26248_, new_n26249_, new_n26250_, new_n26251_, new_n26252_,
    new_n26253_, new_n26254_, new_n26255_, new_n26256_, new_n26257_,
    new_n26258_, new_n26259_, new_n26260_, new_n26261_, new_n26262_,
    new_n26263_, new_n26264_, new_n26265_, new_n26266_, new_n26267_,
    new_n26268_, new_n26269_, new_n26270_, new_n26271_, new_n26272_,
    new_n26273_, new_n26274_, new_n26275_, new_n26276_, new_n26277_,
    new_n26278_, new_n26279_, new_n26280_, new_n26281_, new_n26282_,
    new_n26283_, new_n26284_, new_n26285_, new_n26286_, new_n26287_,
    new_n26288_, new_n26289_, new_n26290_, new_n26291_, new_n26292_,
    new_n26293_, new_n26294_, new_n26295_, new_n26296_, new_n26297_,
    new_n26298_, new_n26299_, new_n26300_, new_n26301_, new_n26302_,
    new_n26303_, new_n26304_, new_n26305_, new_n26306_, new_n26307_,
    new_n26308_, new_n26309_, new_n26310_, new_n26311_, new_n26312_,
    new_n26313_, new_n26314_, new_n26315_, new_n26316_, new_n26317_,
    new_n26318_, new_n26319_, new_n26320_, new_n26321_, new_n26322_,
    new_n26323_, new_n26324_, new_n26325_, new_n26326_, new_n26327_,
    new_n26328_, new_n26329_, new_n26330_, new_n26331_, new_n26332_,
    new_n26333_, new_n26334_, new_n26335_, new_n26336_, new_n26337_,
    new_n26338_, new_n26339_, new_n26340_, new_n26341_, new_n26342_,
    new_n26343_, new_n26344_, new_n26345_, new_n26346_, new_n26347_,
    new_n26348_, new_n26349_, new_n26350_, new_n26351_, new_n26352_,
    new_n26353_, new_n26354_, new_n26355_, new_n26356_, new_n26357_,
    new_n26358_, new_n26360_, new_n26361_, new_n26362_, new_n26363_,
    new_n26364_, new_n26365_, new_n26366_, new_n26367_, new_n26368_,
    new_n26369_, new_n26370_, new_n26371_, new_n26372_, new_n26373_,
    new_n26374_, new_n26375_, new_n26376_, new_n26377_, new_n26378_,
    new_n26379_, new_n26380_, new_n26381_, new_n26382_, new_n26383_,
    new_n26384_, new_n26385_, new_n26386_, new_n26387_, new_n26388_,
    new_n26389_, new_n26390_, new_n26391_, new_n26392_, new_n26393_,
    new_n26394_, new_n26395_, new_n26396_, new_n26397_, new_n26398_,
    new_n26399_, new_n26400_, new_n26401_, new_n26402_, new_n26403_,
    new_n26404_, new_n26405_, new_n26406_, new_n26407_, new_n26408_,
    new_n26409_, new_n26410_, new_n26411_, new_n26412_, new_n26413_,
    new_n26414_, new_n26415_, new_n26416_, new_n26417_, new_n26418_,
    new_n26419_, new_n26420_, new_n26421_, new_n26422_, new_n26423_,
    new_n26424_, new_n26425_, new_n26426_, new_n26427_, new_n26428_,
    new_n26429_, new_n26430_, new_n26431_, new_n26432_, new_n26433_,
    new_n26434_, new_n26435_, new_n26436_, new_n26438_, new_n26439_,
    new_n26440_, new_n26441_, new_n26442_, new_n26443_, new_n26444_,
    new_n26445_, new_n26446_, new_n26447_, new_n26448_, new_n26449_,
    new_n26451_, new_n26452_, new_n26453_, new_n26454_, new_n26455_,
    new_n26456_, new_n26457_, new_n26458_, new_n26459_, new_n26460_,
    new_n26461_, new_n26462_, new_n26463_, new_n26464_, new_n26465_,
    new_n26466_, new_n26467_, new_n26468_, new_n26469_, new_n26470_,
    new_n26471_, new_n26472_, new_n26473_, new_n26474_, new_n26475_,
    new_n26476_, new_n26477_, new_n26478_, new_n26479_, new_n26480_,
    new_n26481_, new_n26482_, new_n26483_, new_n26484_, new_n26485_,
    new_n26486_, new_n26487_, new_n26488_, new_n26489_, new_n26490_,
    new_n26491_, new_n26492_, new_n26493_, new_n26494_, new_n26495_,
    new_n26496_, new_n26497_, new_n26498_, new_n26499_, new_n26500_,
    new_n26501_, new_n26502_, new_n26503_, new_n26504_, new_n26505_,
    new_n26506_, new_n26507_, new_n26508_, new_n26509_, new_n26510_,
    new_n26511_, new_n26513_, new_n26514_, new_n26515_, new_n26516_,
    new_n26517_, new_n26518_, new_n26519_, new_n26520_, new_n26521_,
    new_n26522_, new_n26523_, new_n26524_, new_n26525_, new_n26526_,
    new_n26527_, new_n26528_, new_n26529_, new_n26530_, new_n26531_,
    new_n26532_, new_n26533_, new_n26534_, new_n26535_, new_n26536_,
    new_n26537_, new_n26538_, new_n26539_, new_n26540_, new_n26541_,
    new_n26542_, new_n26543_, new_n26544_, new_n26545_, new_n26546_,
    new_n26547_, new_n26549_, new_n26550_, new_n26551_, new_n26552_,
    new_n26553_, new_n26554_, new_n26555_, new_n26556_, new_n26557_,
    new_n26558_, new_n26559_, new_n26560_, new_n26561_, new_n26562_,
    new_n26563_, new_n26564_, new_n26565_, new_n26566_, new_n26567_,
    new_n26568_, new_n26570_, new_n26571_, new_n26572_, new_n26573_,
    new_n26574_, new_n26575_, new_n26576_, new_n26577_, new_n26578_,
    new_n26579_, new_n26580_, new_n26582_, new_n26583_, new_n26584_,
    new_n26585_, new_n26586_, new_n26589_, new_n26590_, new_n26591_,
    new_n26592_, new_n26593_, new_n26594_, new_n26595_, new_n26596_,
    new_n26597_, new_n26598_, new_n26599_, new_n26600_, new_n26601_,
    new_n26602_, new_n26603_, new_n26604_, new_n26605_, new_n26606_,
    new_n26607_, new_n26608_, new_n26609_, new_n26610_, new_n26611_,
    new_n26612_, new_n26613_, new_n26614_, new_n26615_, new_n26616_,
    new_n26617_, new_n26618_, new_n26619_, new_n26620_, new_n26621_,
    new_n26622_, new_n26623_, new_n26624_, new_n26625_, new_n26626_,
    new_n26627_, new_n26628_, new_n26629_, new_n26630_, new_n26631_,
    new_n26632_, new_n26633_, new_n26634_, new_n26635_, new_n26636_,
    new_n26637_, new_n26638_, new_n26639_, new_n26640_, new_n26641_,
    new_n26642_, new_n26643_, new_n26644_, new_n26645_, new_n26646_,
    new_n26647_, new_n26648_, new_n26649_, new_n26650_, new_n26651_,
    new_n26652_, new_n26653_, new_n26654_, new_n26655_, new_n26656_,
    new_n26657_, new_n26658_, new_n26659_, new_n26660_, new_n26661_,
    new_n26662_, new_n26663_, new_n26664_, new_n26665_, new_n26666_,
    new_n26667_, new_n26668_, new_n26669_, new_n26670_, new_n26671_,
    new_n26672_, new_n26673_, new_n26674_, new_n26675_, new_n26676_,
    new_n26677_, new_n26678_, new_n26679_, new_n26680_, new_n26681_,
    new_n26682_, new_n26683_, new_n26684_, new_n26685_, new_n26686_,
    new_n26687_, new_n26688_, new_n26689_, new_n26690_, new_n26691_,
    new_n26692_, new_n26693_, new_n26694_, new_n26695_, new_n26696_,
    new_n26697_, new_n26698_, new_n26699_, new_n26700_, new_n26701_,
    new_n26702_, new_n26703_, new_n26704_, new_n26705_, new_n26706_,
    new_n26707_, new_n26708_, new_n26709_, new_n26710_, new_n26711_,
    new_n26712_, new_n26713_, new_n26714_, new_n26715_, new_n26716_,
    new_n26717_, new_n26718_, new_n26719_, new_n26720_, new_n26721_,
    new_n26722_, new_n26723_, new_n26724_, new_n26725_, new_n26726_,
    new_n26727_, new_n26728_, new_n26729_, new_n26730_, new_n26731_,
    new_n26732_, new_n26733_, new_n26734_, new_n26735_, new_n26736_,
    new_n26737_, new_n26738_, new_n26739_, new_n26740_, new_n26741_,
    new_n26742_, new_n26743_, new_n26744_, new_n26745_, new_n26746_,
    new_n26747_, new_n26748_, new_n26749_, new_n26750_, new_n26751_,
    new_n26752_, new_n26753_, new_n26754_, new_n26755_, new_n26756_,
    new_n26757_, new_n26758_, new_n26759_, new_n26760_, new_n26761_,
    new_n26762_, new_n26763_, new_n26764_, new_n26765_, new_n26766_,
    new_n26767_, new_n26768_, new_n26769_, new_n26770_, new_n26771_,
    new_n26772_, new_n26773_, new_n26774_, new_n26775_, new_n26776_,
    new_n26777_, new_n26778_, new_n26779_, new_n26780_, new_n26781_,
    new_n26782_, new_n26783_, new_n26784_, new_n26785_, new_n26786_,
    new_n26787_, new_n26788_, new_n26789_, new_n26790_, new_n26791_,
    new_n26792_, new_n26793_, new_n26794_, new_n26795_, new_n26796_,
    new_n26797_, new_n26798_, new_n26799_, new_n26800_, new_n26801_,
    new_n26802_, new_n26803_, new_n26804_, new_n26805_, new_n26806_,
    new_n26807_, new_n26808_, new_n26809_, new_n26810_, new_n26811_,
    new_n26812_, new_n26813_, new_n26814_, new_n26815_, new_n26816_,
    new_n26817_, new_n26818_, new_n26819_, new_n26820_, new_n26821_,
    new_n26822_, new_n26823_, new_n26824_, new_n26825_, new_n26826_,
    new_n26827_, new_n26828_, new_n26829_, new_n26830_, new_n26831_,
    new_n26832_, new_n26833_, new_n26834_, new_n26835_, new_n26836_,
    new_n26837_, new_n26838_, new_n26839_, new_n26840_, new_n26841_,
    new_n26842_, new_n26843_, new_n26844_, new_n26845_, new_n26846_,
    new_n26847_, new_n26848_, new_n26849_, new_n26850_, new_n26851_,
    new_n26852_, new_n26853_, new_n26854_, new_n26855_, new_n26856_,
    new_n26857_, new_n26858_, new_n26859_, new_n26860_, new_n26861_,
    new_n26862_, new_n26863_, new_n26864_, new_n26865_, new_n26866_,
    new_n26867_, new_n26868_, new_n26869_, new_n26870_, new_n26871_,
    new_n26872_, new_n26873_, new_n26874_, new_n26875_, new_n26876_,
    new_n26877_, new_n26878_, new_n26879_, new_n26880_, new_n26881_,
    new_n26882_, new_n26883_, new_n26884_, new_n26885_, new_n26886_,
    new_n26887_, new_n26888_, new_n26889_, new_n26890_, new_n26891_,
    new_n26892_, new_n26893_, new_n26894_, new_n26895_, new_n26896_,
    new_n26897_, new_n26898_, new_n26899_, new_n26900_, new_n26901_,
    new_n26902_, new_n26903_, new_n26904_, new_n26905_, new_n26906_,
    new_n26907_, new_n26908_, new_n26909_, new_n26910_, new_n26911_,
    new_n26912_, new_n26913_, new_n26914_, new_n26915_, new_n26916_,
    new_n26917_, new_n26918_, new_n26919_, new_n26920_, new_n26921_,
    new_n26922_, new_n26923_, new_n26924_, new_n26925_, new_n26926_,
    new_n26927_, new_n26928_, new_n26929_, new_n26930_, new_n26931_,
    new_n26932_, new_n26933_, new_n26934_, new_n26935_, new_n26936_,
    new_n26937_, new_n26938_, new_n26939_, new_n26940_, new_n26941_,
    new_n26942_, new_n26943_, new_n26944_, new_n26945_, new_n26946_,
    new_n26947_, new_n26948_, new_n26949_, new_n26950_, new_n26951_,
    new_n26952_, new_n26953_, new_n26954_, new_n26955_, new_n26956_,
    new_n26957_, new_n26958_, new_n26959_, new_n26960_, new_n26961_,
    new_n26962_, new_n26963_, new_n26964_, new_n26965_, new_n26966_,
    new_n26967_, new_n26968_, new_n26969_, new_n26970_, new_n26971_,
    new_n26972_, new_n26973_, new_n26974_, new_n26975_, new_n26976_,
    new_n26977_, new_n26978_, new_n26979_, new_n26980_, new_n26981_,
    new_n26982_, new_n26983_, new_n26984_, new_n26985_, new_n26986_,
    new_n26987_, new_n26988_, new_n26989_, new_n26990_, new_n26991_,
    new_n26992_, new_n26993_, new_n26994_, new_n26995_, new_n26996_,
    new_n26997_, new_n26998_, new_n26999_, new_n27000_, new_n27001_,
    new_n27002_, new_n27003_, new_n27004_, new_n27005_, new_n27006_,
    new_n27007_, new_n27008_, new_n27009_, new_n27010_, new_n27011_,
    new_n27012_, new_n27013_, new_n27014_, new_n27015_, new_n27016_,
    new_n27017_, new_n27018_, new_n27019_, new_n27020_, new_n27021_,
    new_n27022_, new_n27023_, new_n27024_, new_n27025_, new_n27026_,
    new_n27027_, new_n27028_, new_n27029_, new_n27030_, new_n27031_,
    new_n27033_, new_n27034_, new_n27035_, new_n27036_, new_n27037_,
    new_n27038_, new_n27039_, new_n27040_, new_n27041_, new_n27042_,
    new_n27043_, new_n27044_, new_n27045_, new_n27046_, new_n27047_,
    new_n27048_, new_n27049_, new_n27050_, new_n27051_, new_n27052_,
    new_n27053_, new_n27054_, new_n27055_, new_n27056_, new_n27057_,
    new_n27058_, new_n27059_, new_n27060_, new_n27061_, new_n27062_,
    new_n27063_, new_n27064_, new_n27065_, new_n27066_, new_n27067_,
    new_n27068_, new_n27069_, new_n27070_, new_n27071_, new_n27072_,
    new_n27073_, new_n27074_, new_n27075_, new_n27076_, new_n27077_,
    new_n27078_, new_n27079_, new_n27080_, new_n27081_, new_n27082_,
    new_n27083_, new_n27084_, new_n27085_, new_n27086_, new_n27087_,
    new_n27088_, new_n27089_, new_n27090_, new_n27091_, new_n27092_,
    new_n27093_, new_n27095_, new_n27096_, new_n27097_, new_n27098_,
    new_n27099_, new_n27100_, new_n27101_, new_n27102_, new_n27103_,
    new_n27104_, new_n27105_, new_n27106_, new_n27107_, new_n27108_,
    new_n27109_, new_n27110_, new_n27111_, new_n27112_, new_n27113_,
    new_n27114_, new_n27115_, new_n27116_, new_n27117_, new_n27118_,
    new_n27119_, new_n27120_, new_n27121_, new_n27122_, new_n27123_,
    new_n27124_, new_n27125_, new_n27127_, new_n27128_, new_n27129_,
    new_n27130_, new_n27131_, new_n27132_, new_n27133_, new_n27134_,
    new_n27135_, new_n27136_, new_n27137_, new_n27138_, new_n27139_,
    new_n27140_, new_n27141_, new_n27142_, new_n27143_, new_n27145_,
    new_n27146_, new_n27147_, new_n27148_, new_n27149_, new_n27150_,
    new_n27151_, new_n27152_, new_n27153_, new_n27155_, new_n27156_,
    new_n27157_, new_n27158_, new_n27161_, new_n27162_, new_n27163_,
    new_n27164_, new_n27165_, new_n27166_, new_n27167_, new_n27168_,
    new_n27169_, new_n27170_, new_n27171_, new_n27172_, new_n27173_,
    new_n27174_, new_n27175_, new_n27176_, new_n27177_, new_n27178_,
    new_n27179_, new_n27180_, new_n27181_, new_n27182_, new_n27183_,
    new_n27184_, new_n27185_, new_n27186_, new_n27187_, new_n27188_,
    new_n27189_, new_n27190_, new_n27191_, new_n27192_, new_n27193_,
    new_n27194_, new_n27195_, new_n27196_, new_n27197_, new_n27198_,
    new_n27199_, new_n27200_, new_n27201_, new_n27202_, new_n27203_,
    new_n27204_, new_n27205_, new_n27206_, new_n27207_, new_n27208_,
    new_n27209_, new_n27210_, new_n27211_, new_n27212_, new_n27213_,
    new_n27214_, new_n27215_, new_n27216_, new_n27217_, new_n27218_,
    new_n27219_, new_n27220_, new_n27221_, new_n27222_, new_n27223_,
    new_n27224_, new_n27225_, new_n27226_, new_n27227_, new_n27228_,
    new_n27229_, new_n27230_, new_n27231_, new_n27232_, new_n27233_,
    new_n27234_, new_n27235_, new_n27236_, new_n27237_, new_n27238_,
    new_n27239_, new_n27240_, new_n27241_, new_n27242_, new_n27243_,
    new_n27244_, new_n27245_, new_n27246_, new_n27247_, new_n27248_,
    new_n27249_, new_n27250_, new_n27251_, new_n27252_, new_n27253_,
    new_n27254_, new_n27255_, new_n27256_, new_n27257_, new_n27258_,
    new_n27259_, new_n27260_, new_n27261_, new_n27262_, new_n27263_,
    new_n27264_, new_n27265_, new_n27266_, new_n27267_, new_n27268_,
    new_n27269_, new_n27270_, new_n27271_, new_n27272_, new_n27273_,
    new_n27274_, new_n27275_, new_n27276_, new_n27277_, new_n27278_,
    new_n27279_, new_n27280_, new_n27281_, new_n27282_, new_n27283_,
    new_n27284_, new_n27285_, new_n27286_, new_n27287_, new_n27288_,
    new_n27289_, new_n27290_, new_n27291_, new_n27292_, new_n27293_,
    new_n27294_, new_n27295_, new_n27296_, new_n27297_, new_n27298_,
    new_n27299_, new_n27300_, new_n27301_, new_n27302_, new_n27303_,
    new_n27304_, new_n27305_, new_n27306_, new_n27307_, new_n27308_,
    new_n27309_, new_n27310_, new_n27311_, new_n27312_, new_n27313_,
    new_n27314_, new_n27315_, new_n27316_, new_n27317_, new_n27318_,
    new_n27319_, new_n27320_, new_n27321_, new_n27322_, new_n27323_,
    new_n27324_, new_n27336_, new_n27337_, new_n27338_, new_n27340_,
    new_n27341_, new_n27342_, new_n27343_, new_n27344_, new_n27345_,
    new_n27346_, new_n27347_, new_n27348_, new_n27349_, new_n27350_,
    new_n27351_, new_n27352_, new_n27353_, new_n27354_, new_n27355_,
    new_n27356_, new_n27357_, new_n27358_, new_n27359_, new_n27360_,
    new_n27361_, new_n27362_, new_n27363_, new_n27364_, new_n27365_,
    new_n27366_, new_n27367_, new_n27368_, new_n27369_, new_n27370_,
    new_n27371_, new_n27372_, new_n27373_, new_n27374_, new_n27375_,
    new_n27377_, new_n27378_, new_n27379_, new_n27380_, new_n27381_,
    new_n27382_, new_n27383_, new_n27384_, new_n27385_, new_n27386_,
    new_n27387_, new_n27388_, new_n27389_, new_n27391_, new_n27392_,
    new_n27393_, new_n27394_, new_n27395_, new_n27396_, new_n27397_,
    new_n27398_, new_n27399_, new_n27400_, new_n27401_, new_n27402_,
    new_n27403_, new_n27404_, new_n27405_, new_n27406_, new_n27407_,
    new_n27408_, new_n27409_, new_n27410_, new_n27411_, new_n27412_,
    new_n27413_, new_n27414_, new_n27415_, new_n27416_, new_n27417_,
    new_n27418_, new_n27419_, new_n27420_, new_n27421_, new_n27422_,
    new_n27423_, new_n27424_, new_n27425_, new_n27426_, new_n27427_,
    new_n27428_, new_n27429_, new_n27430_, new_n27431_, new_n27432_,
    new_n27433_, new_n27434_, new_n27435_, new_n27436_, new_n27437_,
    new_n27438_, new_n27439_, new_n27440_, new_n27441_, new_n27442_,
    new_n27443_, new_n27444_, new_n27445_, new_n27446_, new_n27447_,
    new_n27448_, new_n27449_, new_n27450_, new_n27451_, new_n27452_,
    new_n27453_, new_n27454_, new_n27455_, new_n27456_, new_n27457_,
    new_n27458_, new_n27459_, new_n27460_, new_n27461_, new_n27462_,
    new_n27463_, new_n27464_, new_n27465_, new_n27466_, new_n27467_,
    new_n27468_, new_n27469_, new_n27470_, new_n27471_, new_n27472_,
    new_n27473_, new_n27474_, new_n27475_, new_n27476_, new_n27477_,
    new_n27478_, new_n27480_, new_n27481_, new_n27482_, new_n27483_,
    new_n27484_, new_n27485_, new_n27488_, new_n27489_, new_n27490_,
    new_n27491_, new_n27492_, new_n27493_, new_n27494_, new_n27495_,
    new_n27496_, new_n27497_, new_n27498_, new_n27499_, new_n27500_,
    new_n27501_, new_n27502_, new_n27503_, new_n27504_, new_n27505_,
    new_n27506_, new_n27507_, new_n27508_, new_n27509_, new_n27510_,
    new_n27511_, new_n27512_, new_n27513_, new_n27514_, new_n27515_,
    new_n27516_, new_n27517_, new_n27518_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27623_, new_n27624_, new_n27625_,
    new_n27626_, new_n27627_, new_n27628_, new_n27629_, new_n27630_,
    new_n27631_, new_n27632_, new_n27633_, new_n27634_, new_n27635_,
    new_n27636_, new_n27637_, new_n27638_, new_n27639_, new_n27640_,
    new_n27641_, new_n27642_, new_n27643_, new_n27644_, new_n27645_,
    new_n27646_, new_n27647_, new_n27648_, new_n27649_, new_n27650_,
    new_n27651_, new_n27652_, new_n27653_, new_n27654_, new_n27655_,
    new_n27656_, new_n27657_, new_n27658_, new_n27659_, new_n27660_,
    new_n27661_, new_n27662_, new_n27663_, new_n27664_, new_n27665_,
    new_n27666_, new_n27667_, new_n27668_, new_n27669_, new_n27670_,
    new_n27671_, new_n27672_, new_n27673_, new_n27674_, new_n27675_,
    new_n27676_, new_n27677_, new_n27678_, new_n27679_, new_n27680_,
    new_n27681_, new_n27682_, new_n27683_, new_n27684_, new_n27685_,
    new_n27686_, new_n27687_, new_n27688_, new_n27689_, new_n27690_,
    new_n27691_, new_n27692_, new_n27693_, new_n27694_, new_n27695_,
    new_n27696_, new_n27697_, new_n27698_, new_n27699_, new_n27700_,
    new_n27701_, new_n27702_, new_n27703_, new_n27704_, new_n27705_,
    new_n27706_, new_n27707_, new_n27708_, new_n27709_, new_n27710_,
    new_n27711_, new_n27712_, new_n27713_, new_n27714_, new_n27715_,
    new_n27716_, new_n27717_, new_n27718_, new_n27720_, new_n27721_,
    new_n27722_, new_n27723_, new_n27724_, new_n27725_, new_n27726_,
    new_n27727_, new_n27728_, new_n27729_, new_n27730_, new_n27731_,
    new_n27732_, new_n27733_, new_n27734_, new_n27735_, new_n27736_,
    new_n27737_, new_n27738_, new_n27739_, new_n27740_, new_n27741_,
    new_n27742_, new_n27743_, new_n27744_, new_n27745_, new_n27746_,
    new_n27747_, new_n27748_, new_n27749_, new_n27750_, new_n27751_,
    new_n27752_, new_n27753_, new_n27754_, new_n27755_, new_n27756_,
    new_n27757_, new_n27758_, new_n27759_, new_n27760_, new_n27761_,
    new_n27762_, new_n27763_, new_n27764_, new_n27765_, new_n27766_,
    new_n27767_, new_n27768_, new_n27769_, new_n27770_, new_n27771_,
    new_n27772_, new_n27773_, new_n27774_, new_n27775_, new_n27777_,
    new_n27778_, new_n27779_, new_n27780_, new_n27781_, new_n27782_,
    new_n27783_, new_n27784_, new_n27785_, new_n27786_, new_n27787_,
    new_n27788_, new_n27789_, new_n27790_, new_n27791_, new_n27792_,
    new_n27793_, new_n27794_, new_n27795_, new_n27796_, new_n27797_,
    new_n27798_, new_n27799_, new_n27800_, new_n27801_, new_n27802_,
    new_n27803_, new_n27804_, new_n27805_, new_n27806_, new_n27807_,
    new_n27808_, new_n27809_, new_n27810_, new_n27812_, new_n27813_,
    new_n27814_, new_n27815_, new_n27816_, new_n27817_, new_n27818_,
    new_n27819_, new_n27820_, new_n27821_, new_n27822_, new_n27823_,
    new_n27824_, new_n27825_, new_n27826_, new_n27827_, new_n27828_,
    new_n27829_, new_n27830_, new_n27831_, new_n27833_, new_n27834_,
    new_n27835_, new_n27836_, new_n27837_, new_n27838_, new_n27839_,
    new_n27840_, new_n27841_, new_n27842_, new_n27843_, new_n27845_,
    new_n27846_, new_n27847_, new_n27848_, new_n27849_;
  assign \o[0]  = new_n6345_ ^ new_n13445_;
  assign new_n6345_ = new_n6346_ ? (~new_n12722_ ^ new_n13278_) : (new_n12722_ ^ new_n13278_);
  assign new_n6346_ = new_n6347_ ? (new_n10371_ ^ new_n12451_) : (~new_n10371_ ^ new_n12451_);
  assign new_n6347_ = new_n6348_ ? (new_n8812_ ^ new_n10163_) : (~new_n8812_ ^ new_n10163_);
  assign new_n6348_ = new_n6349_ ? (new_n7594_ ^ new_n8538_) : (~new_n7594_ ^ new_n8538_);
  assign new_n6349_ = new_n6350_ ? (new_n6843_ ^ new_n7261_) : (~new_n6843_ ^ new_n7261_);
  assign new_n6350_ = new_n6767_ & (new_n6842_ | ~new_n6351_);
  assign new_n6351_ = ~new_n6601_ & new_n6352_ & (new_n6736_ | ~new_n6701_ | ~new_n6700_);
  assign new_n6352_ = (~new_n6353_ | ~new_n6567_) & (~new_n6496_ | ~new_n6459_);
  assign new_n6353_ = new_n6354_ & ~new_n6389_ & ~new_n6425_;
  assign new_n6354_ = new_n6355_ & new_n6384_;
  assign new_n6355_ = ~new_n6356_ & ~new_n6378_;
  assign new_n6356_ = ~new_n6357_ & (\all_features[3043]  | \all_features[3044]  | \all_features[3045]  | \all_features[3046]  | \all_features[3047] );
  assign new_n6357_ = ~new_n6375_ & (new_n6373_ | (~new_n6376_ & (new_n6377_ | (~new_n6358_ & ~new_n6371_))));
  assign new_n6358_ = ~new_n6368_ & (new_n6370_ | new_n6359_);
  assign new_n6359_ = \all_features[3047]  & ((new_n6360_ & (\all_features[3046]  | \all_features[3045] )) | (~\all_features[3046]  & (\all_features[3045]  ? new_n6366_ : \all_features[3044] )));
  assign new_n6360_ = new_n6361_ & (\all_features[3045]  | ~new_n6364_ | (~new_n6365_ & ~\all_features[3044]  & new_n6363_) | (\all_features[3044]  & ~new_n6363_));
  assign new_n6361_ = \all_features[3047]  & (\all_features[3046]  | (new_n6362_ & (\all_features[3042]  | \all_features[3043]  | \all_features[3041] )));
  assign new_n6362_ = \all_features[3044]  & \all_features[3045] ;
  assign new_n6363_ = ~\all_features[3042]  & ~\all_features[3043] ;
  assign new_n6364_ = \all_features[3046]  & \all_features[3047] ;
  assign new_n6365_ = \all_features[3040]  & \all_features[3041] ;
  assign new_n6366_ = new_n6363_ & ~\all_features[3044]  & new_n6367_;
  assign new_n6367_ = ~\all_features[3040]  & ~\all_features[3041] ;
  assign new_n6368_ = ~new_n6369_ & ~\all_features[3047] ;
  assign new_n6369_ = \all_features[3045]  & \all_features[3046]  & (\all_features[3044]  | (\all_features[3042]  & \all_features[3043]  & \all_features[3041] ));
  assign new_n6370_ = ~\all_features[3047]  & (~new_n6362_ | ~\all_features[3042]  | ~\all_features[3043]  | ~\all_features[3046]  | ~new_n6365_);
  assign new_n6371_ = ~\all_features[3047]  & (~\all_features[3046]  | new_n6372_);
  assign new_n6372_ = ~\all_features[3045]  & (new_n6367_ | ~\all_features[3043]  | ~\all_features[3044]  | ~\all_features[3042] );
  assign new_n6373_ = new_n6374_ & (~\all_features[3045]  | (~\all_features[3044]  & (~\all_features[3043]  | (~\all_features[3042]  & ~\all_features[3041] ))));
  assign new_n6374_ = ~\all_features[3046]  & ~\all_features[3047] ;
  assign new_n6375_ = ~\all_features[3045]  & new_n6374_ & ((~\all_features[3042]  & new_n6367_) | ~\all_features[3044]  | ~\all_features[3043] );
  assign new_n6376_ = new_n6374_ & (~\all_features[3043]  | ~new_n6362_ | (~\all_features[3042]  & ~new_n6365_));
  assign new_n6377_ = ~\all_features[3047]  & (~\all_features[3046]  | (~\all_features[3045]  & ~\all_features[3044]  & (~\all_features[3043]  | ~\all_features[3042] )));
  assign new_n6378_ = new_n6383_ & (new_n6376_ | new_n6373_ | (~new_n6379_ & ~new_n6371_ & ~new_n6377_));
  assign new_n6379_ = ~new_n6370_ & ~new_n6368_ & (~new_n6380_ | (~new_n6382_ & new_n6361_ & new_n6381_));
  assign new_n6380_ = \all_features[3047]  & (\all_features[3046]  | (~new_n6366_ & \all_features[3045] ));
  assign new_n6381_ = new_n6364_ & (new_n6365_ | \all_features[3044]  | \all_features[3045]  | ~new_n6363_);
  assign new_n6382_ = new_n6364_ & \all_features[3045]  & ((~new_n6367_ & \all_features[3042] ) | \all_features[3044]  | \all_features[3043] );
  assign new_n6383_ = ~new_n6375_ & (\all_features[3043]  | \all_features[3044]  | \all_features[3045]  | \all_features[3046]  | \all_features[3047] );
  assign new_n6384_ = ~new_n6385_ & ~new_n6388_;
  assign new_n6385_ = new_n6383_ & ~new_n6376_ & ~new_n6386_ & ~new_n6373_;
  assign new_n6386_ = ~new_n6371_ & ~new_n6370_ & new_n6387_ & (~new_n6361_ | ~new_n6381_ | ~new_n6380_);
  assign new_n6387_ = ~new_n6368_ & ~new_n6377_;
  assign new_n6388_ = new_n6387_ & new_n6383_ & ~new_n6376_ & ~new_n6373_ & ~new_n6371_ & ~new_n6370_;
  assign new_n6389_ = new_n6390_ & ~new_n6421_ & ~new_n6424_;
  assign new_n6390_ = ~new_n6391_ & ~new_n6411_;
  assign new_n6391_ = (new_n6392_ | (~new_n6410_ & ~\all_features[3701]  & new_n6406_)) & (\all_features[3699]  | \all_features[3700]  | \all_features[3701]  | ~new_n6406_);
  assign new_n6392_ = ~new_n6405_ & (new_n6407_ | (~new_n6408_ & (new_n6409_ | new_n6393_)));
  assign new_n6393_ = ~new_n6400_ & (new_n6402_ | (~new_n6394_ & new_n6404_));
  assign new_n6394_ = \all_features[3703]  & ((~new_n6399_ & ~\all_features[3701]  & \all_features[3702] ) | (~new_n6397_ & (\all_features[3702]  | (~new_n6395_ & \all_features[3701] ))));
  assign new_n6395_ = new_n6396_ & ~\all_features[3700]  & ~\all_features[3698]  & ~\all_features[3699] ;
  assign new_n6396_ = ~\all_features[3696]  & ~\all_features[3697] ;
  assign new_n6397_ = \all_features[3703]  & (\all_features[3702]  | (new_n6398_ & (\all_features[3698]  | \all_features[3699]  | \all_features[3697] )));
  assign new_n6398_ = \all_features[3700]  & \all_features[3701] ;
  assign new_n6399_ = (~\all_features[3698]  & ~\all_features[3699]  & ~\all_features[3700]  & (~\all_features[3697]  | ~\all_features[3696] )) | (\all_features[3700]  & (\all_features[3698]  | \all_features[3699] ));
  assign new_n6400_ = ~new_n6401_ & ~\all_features[3703] ;
  assign new_n6401_ = \all_features[3701]  & \all_features[3702]  & (\all_features[3700]  | (\all_features[3698]  & \all_features[3699]  & \all_features[3697] ));
  assign new_n6402_ = ~\all_features[3703]  & (~new_n6403_ | ~\all_features[3696]  | ~\all_features[3697]  | ~\all_features[3702]  | ~new_n6398_);
  assign new_n6403_ = \all_features[3698]  & \all_features[3699] ;
  assign new_n6404_ = \all_features[3703]  & (\all_features[3701]  | \all_features[3702]  | \all_features[3700] );
  assign new_n6405_ = new_n6406_ & (~\all_features[3701]  | (~\all_features[3700]  & (~\all_features[3699]  | (~\all_features[3698]  & ~\all_features[3697] ))));
  assign new_n6406_ = ~\all_features[3702]  & ~\all_features[3703] ;
  assign new_n6407_ = new_n6406_ & (~new_n6398_ | ~\all_features[3699]  | (~\all_features[3698]  & (~\all_features[3696]  | ~\all_features[3697] )));
  assign new_n6408_ = ~\all_features[3703]  & (~\all_features[3702]  | (~\all_features[3700]  & ~\all_features[3701]  & ~new_n6403_));
  assign new_n6409_ = ~\all_features[3703]  & (~\all_features[3702]  | (~\all_features[3701]  & (new_n6396_ | ~new_n6403_ | ~\all_features[3700] )));
  assign new_n6410_ = \all_features[3699]  & \all_features[3700]  & (\all_features[3698]  | ~new_n6396_);
  assign new_n6411_ = new_n6417_ & (~new_n6418_ | (new_n6419_ & (~new_n6420_ | new_n6412_)));
  assign new_n6412_ = new_n6413_ & (~new_n6414_ | (~new_n6416_ & \all_features[3701]  & \all_features[3702]  & \all_features[3703] ));
  assign new_n6413_ = \all_features[3703]  & (\all_features[3702]  | (~new_n6395_ & \all_features[3701] ));
  assign new_n6414_ = \all_features[3703]  & \all_features[3702]  & ~new_n6415_ & new_n6397_;
  assign new_n6415_ = ~\all_features[3698]  & ~\all_features[3699]  & ~\all_features[3700]  & ~\all_features[3701]  & (~\all_features[3697]  | ~\all_features[3696] );
  assign new_n6416_ = ~\all_features[3699]  & ~\all_features[3700]  & (~\all_features[3698]  | new_n6396_);
  assign new_n6417_ = \all_features[3701]  | ~new_n6406_ | (new_n6410_ & (\all_features[3699]  | \all_features[3700] ));
  assign new_n6418_ = ~new_n6405_ & ~new_n6407_;
  assign new_n6419_ = ~new_n6408_ & ~new_n6409_;
  assign new_n6420_ = ~new_n6400_ & ~new_n6402_;
  assign new_n6421_ = new_n6422_ & (new_n6409_ | new_n6400_ | ~new_n6423_ | (new_n6414_ & new_n6413_));
  assign new_n6422_ = new_n6417_ & new_n6418_;
  assign new_n6423_ = ~new_n6408_ & ~new_n6402_;
  assign new_n6424_ = new_n6420_ & new_n6422_ & new_n6419_;
  assign new_n6425_ = new_n6426_ & (new_n6456_ | new_n6450_);
  assign new_n6426_ = new_n6427_ & new_n6448_;
  assign new_n6427_ = new_n6445_ & ~new_n6428_ & new_n6442_;
  assign new_n6428_ = ~new_n6436_ & ~new_n6438_ & ~new_n6440_ & ~new_n6441_ & (~new_n6433_ | ~new_n6429_);
  assign new_n6429_ = \all_features[3103]  & \all_features[3102]  & ~new_n6432_ & new_n6430_;
  assign new_n6430_ = \all_features[3103]  & (\all_features[3102]  | (new_n6431_ & (\all_features[3098]  | \all_features[3099]  | \all_features[3097] )));
  assign new_n6431_ = \all_features[3100]  & \all_features[3101] ;
  assign new_n6432_ = ~\all_features[3098]  & ~\all_features[3099]  & ~\all_features[3100]  & ~\all_features[3101]  & (~\all_features[3097]  | ~\all_features[3096] );
  assign new_n6433_ = \all_features[3103]  & (\all_features[3102]  | (~new_n6434_ & \all_features[3101] ));
  assign new_n6434_ = new_n6435_ & ~\all_features[3100]  & ~\all_features[3098]  & ~\all_features[3099] ;
  assign new_n6435_ = ~\all_features[3096]  & ~\all_features[3097] ;
  assign new_n6436_ = ~\all_features[3103]  & (~\all_features[3102]  | (~\all_features[3101]  & (new_n6435_ | ~new_n6437_ | ~\all_features[3100] )));
  assign new_n6437_ = \all_features[3098]  & \all_features[3099] ;
  assign new_n6438_ = ~new_n6439_ & ~\all_features[3103] ;
  assign new_n6439_ = \all_features[3101]  & \all_features[3102]  & (\all_features[3100]  | (\all_features[3098]  & \all_features[3099]  & \all_features[3097] ));
  assign new_n6440_ = ~\all_features[3103]  & (~new_n6437_ | ~\all_features[3096]  | ~\all_features[3097]  | ~\all_features[3102]  | ~new_n6431_);
  assign new_n6441_ = ~\all_features[3103]  & (~\all_features[3102]  | (~\all_features[3100]  & ~\all_features[3101]  & ~new_n6437_));
  assign new_n6442_ = ~new_n6443_ | (\all_features[3099]  & \all_features[3100]  & (\all_features[3098]  | ~new_n6435_));
  assign new_n6443_ = ~\all_features[3101]  & new_n6444_;
  assign new_n6444_ = ~\all_features[3102]  & ~\all_features[3103] ;
  assign new_n6445_ = ~new_n6446_ & ~new_n6447_;
  assign new_n6446_ = new_n6444_ & (~new_n6431_ | ~\all_features[3099]  | (~\all_features[3098]  & (~\all_features[3096]  | ~\all_features[3097] )));
  assign new_n6447_ = new_n6444_ & (~\all_features[3101]  | (~\all_features[3100]  & (~\all_features[3099]  | (~\all_features[3098]  & ~\all_features[3097] ))));
  assign new_n6448_ = new_n6445_ & new_n6442_ & new_n6449_ & ~new_n6438_ & ~new_n6440_;
  assign new_n6449_ = ~new_n6436_ & ~new_n6441_;
  assign new_n6450_ = (new_n6451_ | (new_n6443_ & (~\all_features[3099]  | ~\all_features[3100]  | (~\all_features[3098]  & new_n6435_)))) & (~new_n6443_ | \all_features[3099]  | \all_features[3100] );
  assign new_n6451_ = ~new_n6447_ & (new_n6446_ | (~new_n6441_ & ~new_n6452_));
  assign new_n6452_ = ~new_n6436_ & (new_n6438_ | (~new_n6440_ & (~new_n6455_ | new_n6453_)));
  assign new_n6453_ = \all_features[3103]  & ((~new_n6454_ & ~\all_features[3101]  & \all_features[3102] ) | (~new_n6430_ & (\all_features[3102]  | (~new_n6434_ & \all_features[3101] ))));
  assign new_n6454_ = (~\all_features[3098]  & ~\all_features[3099]  & ~\all_features[3100]  & (~\all_features[3097]  | ~\all_features[3096] )) | (\all_features[3100]  & (\all_features[3098]  | \all_features[3099] ));
  assign new_n6455_ = \all_features[3103]  & (\all_features[3101]  | \all_features[3102]  | \all_features[3100] );
  assign new_n6456_ = new_n6442_ & (~new_n6445_ | (new_n6449_ & (new_n6457_ | new_n6438_ | new_n6440_)));
  assign new_n6457_ = new_n6433_ & (~new_n6429_ | (~new_n6458_ & \all_features[3101]  & \all_features[3102]  & \all_features[3103] ));
  assign new_n6458_ = ~\all_features[3099]  & ~\all_features[3100]  & (~\all_features[3098]  | new_n6435_);
  assign new_n6459_ = ~new_n6354_ & ~new_n6460_;
  assign new_n6460_ = new_n6461_ & new_n6490_;
  assign new_n6461_ = new_n6462_ & new_n6484_;
  assign new_n6462_ = ~new_n6463_ & ~new_n6483_;
  assign new_n6463_ = ~new_n6481_ & (new_n6480_ | (~new_n6478_ & (new_n6482_ | (~new_n6464_ & ~new_n6467_))));
  assign new_n6464_ = ~\all_features[2135]  & (~\all_features[2134]  | new_n6465_);
  assign new_n6465_ = ~\all_features[2133]  & (new_n6466_ | ~\all_features[2131]  | ~\all_features[2132]  | ~\all_features[2130] );
  assign new_n6466_ = ~\all_features[2128]  & ~\all_features[2129] ;
  assign new_n6467_ = ~new_n6471_ & (new_n6468_ | (new_n6477_ & (~new_n6473_ | (~new_n6476_ & new_n6475_))));
  assign new_n6468_ = ~\all_features[2135]  & (~new_n6470_ | ~\all_features[2130]  | ~\all_features[2131]  | ~\all_features[2134]  | ~new_n6469_);
  assign new_n6469_ = \all_features[2128]  & \all_features[2129] ;
  assign new_n6470_ = \all_features[2132]  & \all_features[2133] ;
  assign new_n6471_ = ~new_n6472_ & ~\all_features[2135] ;
  assign new_n6472_ = \all_features[2133]  & \all_features[2134]  & (\all_features[2132]  | (\all_features[2130]  & \all_features[2131]  & \all_features[2129] ));
  assign new_n6473_ = \all_features[2135]  & (\all_features[2134]  | (\all_features[2133]  & (\all_features[2132]  | ~new_n6474_ | ~new_n6466_)));
  assign new_n6474_ = ~\all_features[2130]  & ~\all_features[2131] ;
  assign new_n6475_ = \all_features[2135]  & (\all_features[2134]  | (new_n6470_ & (\all_features[2130]  | \all_features[2131]  | \all_features[2129] )));
  assign new_n6476_ = ~\all_features[2133]  & \all_features[2134]  & \all_features[2135]  & (\all_features[2132]  ? new_n6474_ : (new_n6469_ | ~new_n6474_));
  assign new_n6477_ = \all_features[2135]  & (\all_features[2133]  | \all_features[2134]  | \all_features[2132] );
  assign new_n6478_ = new_n6479_ & (~\all_features[2131]  | ~new_n6470_ | (~\all_features[2130]  & ~new_n6469_));
  assign new_n6479_ = ~\all_features[2134]  & ~\all_features[2135] ;
  assign new_n6480_ = new_n6479_ & (~\all_features[2133]  | (~\all_features[2132]  & (~\all_features[2131]  | (~\all_features[2130]  & ~\all_features[2129] ))));
  assign new_n6481_ = ~\all_features[2133]  & new_n6479_ & ((~\all_features[2130]  & new_n6466_) | ~\all_features[2132]  | ~\all_features[2131] );
  assign new_n6482_ = ~\all_features[2135]  & (~\all_features[2134]  | (~\all_features[2133]  & ~\all_features[2132]  & (~\all_features[2131]  | ~\all_features[2130] )));
  assign new_n6483_ = ~\all_features[2135]  & ~\all_features[2134]  & ~\all_features[2133]  & ~\all_features[2131]  & ~\all_features[2132] ;
  assign new_n6484_ = ~new_n6483_ & ~new_n6481_ & (~new_n6489_ | (~new_n6485_ & ~new_n6464_ & ~new_n6482_));
  assign new_n6485_ = ~new_n6468_ & ~new_n6471_ & (~new_n6477_ | ~new_n6473_ | new_n6486_);
  assign new_n6486_ = new_n6475_ & new_n6487_ & (new_n6488_ | ~\all_features[2133]  | ~\all_features[2134]  | ~\all_features[2135] );
  assign new_n6487_ = \all_features[2134]  & \all_features[2135]  & (\all_features[2132]  | \all_features[2133]  | new_n6469_ | ~new_n6474_);
  assign new_n6488_ = ~\all_features[2131]  & ~\all_features[2132]  & (~\all_features[2130]  | new_n6466_);
  assign new_n6489_ = ~new_n6478_ & ~new_n6480_;
  assign new_n6490_ = new_n6491_ & new_n6495_;
  assign new_n6491_ = ~new_n6483_ & ~new_n6481_ & ~new_n6480_ & ~new_n6492_ & ~new_n6478_;
  assign new_n6492_ = ~new_n6464_ & ~new_n6468_ & new_n6493_ & (~new_n6473_ | ~new_n6494_);
  assign new_n6493_ = ~new_n6471_ & ~new_n6482_;
  assign new_n6494_ = new_n6477_ & new_n6475_ & new_n6487_;
  assign new_n6495_ = new_n6489_ & new_n6493_ & ~new_n6483_ & ~new_n6468_ & ~new_n6464_ & ~new_n6481_;
  assign new_n6496_ = new_n6497_ & new_n6533_;
  assign new_n6497_ = ~new_n6498_ & new_n6528_;
  assign new_n6498_ = new_n6499_ & new_n6521_;
  assign new_n6499_ = ~new_n6500_ & (\all_features[2803]  | \all_features[2804]  | \all_features[2805]  | \all_features[2806]  | \all_features[2807] );
  assign new_n6500_ = ~new_n6515_ & (new_n6520_ | (~new_n6517_ & (new_n6518_ | (~new_n6519_ & ~new_n6501_))));
  assign new_n6501_ = ~new_n6511_ & (new_n6513_ | new_n6502_);
  assign new_n6502_ = \all_features[2807]  & ((new_n6503_ & (\all_features[2806]  | \all_features[2805] )) | (~\all_features[2806]  & (\all_features[2805]  ? new_n6509_ : \all_features[2804] )));
  assign new_n6503_ = new_n6504_ & (\all_features[2805]  | ~new_n6508_ | (~new_n6506_ & ~\all_features[2804]  & new_n6507_) | (\all_features[2804]  & ~new_n6507_));
  assign new_n6504_ = \all_features[2807]  & (\all_features[2806]  | (new_n6505_ & (\all_features[2802]  | \all_features[2803]  | \all_features[2801] )));
  assign new_n6505_ = \all_features[2804]  & \all_features[2805] ;
  assign new_n6506_ = \all_features[2800]  & \all_features[2801] ;
  assign new_n6507_ = ~\all_features[2802]  & ~\all_features[2803] ;
  assign new_n6508_ = \all_features[2806]  & \all_features[2807] ;
  assign new_n6509_ = new_n6510_ & ~\all_features[2804]  & new_n6507_;
  assign new_n6510_ = ~\all_features[2800]  & ~\all_features[2801] ;
  assign new_n6511_ = ~new_n6512_ & ~\all_features[2807] ;
  assign new_n6512_ = \all_features[2805]  & \all_features[2806]  & (\all_features[2804]  | (\all_features[2802]  & \all_features[2803]  & \all_features[2801] ));
  assign new_n6513_ = ~\all_features[2807]  & (~\all_features[2806]  | ~new_n6506_ | ~new_n6505_ | ~new_n6514_);
  assign new_n6514_ = \all_features[2802]  & \all_features[2803] ;
  assign new_n6515_ = ~\all_features[2805]  & new_n6516_ & ((~\all_features[2802]  & new_n6510_) | ~\all_features[2804]  | ~\all_features[2803] );
  assign new_n6516_ = ~\all_features[2806]  & ~\all_features[2807] ;
  assign new_n6517_ = new_n6516_ & (~\all_features[2803]  | ~new_n6505_ | (~\all_features[2802]  & ~new_n6506_));
  assign new_n6518_ = ~\all_features[2807]  & (~\all_features[2806]  | (~\all_features[2804]  & ~\all_features[2805]  & ~new_n6514_));
  assign new_n6519_ = ~\all_features[2807]  & (~\all_features[2806]  | (~\all_features[2805]  & (new_n6510_ | ~new_n6514_ | ~\all_features[2804] )));
  assign new_n6520_ = new_n6516_ & (~\all_features[2805]  | (~\all_features[2804]  & (~\all_features[2803]  | (~\all_features[2802]  & ~\all_features[2801] ))));
  assign new_n6521_ = new_n6526_ & (~new_n6527_ | (~new_n6522_ & ~new_n6518_ & ~new_n6519_));
  assign new_n6522_ = ~new_n6513_ & ~new_n6511_ & (~new_n6523_ | (~new_n6525_ & new_n6504_ & new_n6524_));
  assign new_n6523_ = \all_features[2807]  & (\all_features[2806]  | (~new_n6509_ & \all_features[2805] ));
  assign new_n6524_ = new_n6508_ & (new_n6506_ | \all_features[2804]  | \all_features[2805]  | ~new_n6507_);
  assign new_n6525_ = new_n6508_ & \all_features[2805]  & ((~new_n6510_ & \all_features[2802] ) | \all_features[2804]  | \all_features[2803] );
  assign new_n6526_ = ~new_n6515_ & (\all_features[2803]  | \all_features[2804]  | \all_features[2805]  | \all_features[2806]  | \all_features[2807] );
  assign new_n6527_ = ~new_n6517_ & ~new_n6520_;
  assign new_n6528_ = ~new_n6529_ & ~new_n6532_;
  assign new_n6529_ = new_n6527_ & ~new_n6530_ & new_n6526_;
  assign new_n6530_ = ~new_n6519_ & ~new_n6513_ & new_n6531_ & (~new_n6524_ | ~new_n6504_ | ~new_n6523_);
  assign new_n6531_ = ~new_n6518_ & ~new_n6511_;
  assign new_n6532_ = new_n6531_ & new_n6526_ & ~new_n6520_ & ~new_n6513_ & ~new_n6517_ & ~new_n6519_;
  assign new_n6533_ = new_n6534_ & ~new_n6563_ & ~new_n6566_;
  assign new_n6534_ = ~new_n6535_ & ~new_n6556_;
  assign new_n6535_ = ~new_n6536_ & (\all_features[3483]  | \all_features[3484]  | \all_features[3485]  | \all_features[3486]  | \all_features[3487] );
  assign new_n6536_ = ~new_n6550_ & (new_n6552_ | (~new_n6553_ & (new_n6554_ | (~new_n6537_ & ~new_n6555_))));
  assign new_n6537_ = ~new_n6538_ & (new_n6540_ | (new_n6549_ & (~new_n6544_ | (~new_n6548_ & new_n6547_))));
  assign new_n6538_ = ~new_n6539_ & ~\all_features[3487] ;
  assign new_n6539_ = \all_features[3485]  & \all_features[3486]  & (\all_features[3484]  | (\all_features[3482]  & \all_features[3483]  & \all_features[3481] ));
  assign new_n6540_ = ~\all_features[3487]  & (~\all_features[3486]  | ~new_n6541_ | ~new_n6542_ | ~new_n6543_);
  assign new_n6541_ = \all_features[3480]  & \all_features[3481] ;
  assign new_n6542_ = \all_features[3484]  & \all_features[3485] ;
  assign new_n6543_ = \all_features[3482]  & \all_features[3483] ;
  assign new_n6544_ = \all_features[3487]  & (\all_features[3486]  | (\all_features[3485]  & (\all_features[3484]  | ~new_n6546_ | ~new_n6545_)));
  assign new_n6545_ = ~\all_features[3480]  & ~\all_features[3481] ;
  assign new_n6546_ = ~\all_features[3482]  & ~\all_features[3483] ;
  assign new_n6547_ = \all_features[3487]  & (\all_features[3486]  | (new_n6542_ & (\all_features[3482]  | \all_features[3483]  | \all_features[3481] )));
  assign new_n6548_ = ~\all_features[3485]  & \all_features[3486]  & \all_features[3487]  & (\all_features[3484]  ? new_n6546_ : (new_n6541_ | ~new_n6546_));
  assign new_n6549_ = \all_features[3487]  & (\all_features[3485]  | \all_features[3486]  | \all_features[3484] );
  assign new_n6550_ = ~\all_features[3485]  & new_n6551_ & ((~\all_features[3482]  & new_n6545_) | ~\all_features[3484]  | ~\all_features[3483] );
  assign new_n6551_ = ~\all_features[3486]  & ~\all_features[3487] ;
  assign new_n6552_ = new_n6551_ & (~\all_features[3485]  | (~\all_features[3484]  & (~\all_features[3483]  | (~\all_features[3482]  & ~\all_features[3481] ))));
  assign new_n6553_ = new_n6551_ & (~\all_features[3483]  | ~new_n6542_ | (~\all_features[3482]  & ~new_n6541_));
  assign new_n6554_ = ~\all_features[3487]  & (~\all_features[3486]  | (~\all_features[3484]  & ~\all_features[3485]  & ~new_n6543_));
  assign new_n6555_ = ~\all_features[3487]  & (~\all_features[3486]  | (~\all_features[3485]  & (new_n6545_ | ~new_n6543_ | ~\all_features[3484] )));
  assign new_n6556_ = new_n6562_ & (~new_n6561_ | (~new_n6557_ & ~new_n6554_ & ~new_n6555_));
  assign new_n6557_ = ~new_n6538_ & ~new_n6540_ & (~new_n6549_ | ~new_n6544_ | new_n6558_);
  assign new_n6558_ = new_n6547_ & new_n6559_ & (new_n6560_ | ~\all_features[3485]  | ~\all_features[3486]  | ~\all_features[3487] );
  assign new_n6559_ = \all_features[3486]  & \all_features[3487]  & (\all_features[3484]  | \all_features[3485]  | new_n6541_ | ~new_n6546_);
  assign new_n6560_ = ~\all_features[3483]  & ~\all_features[3484]  & (~\all_features[3482]  | new_n6545_);
  assign new_n6561_ = ~new_n6552_ & ~new_n6553_;
  assign new_n6562_ = ~new_n6550_ & (\all_features[3483]  | \all_features[3484]  | \all_features[3485]  | \all_features[3486]  | \all_features[3487] );
  assign new_n6563_ = new_n6561_ & new_n6562_ & (new_n6564_ | new_n6555_ | new_n6540_ | ~new_n6565_);
  assign new_n6564_ = new_n6549_ & new_n6559_ & new_n6544_ & new_n6547_;
  assign new_n6565_ = ~new_n6554_ & ~new_n6538_;
  assign new_n6566_ = new_n6562_ & new_n6561_ & new_n6565_ & ~new_n6555_ & ~new_n6540_;
  assign new_n6567_ = new_n6568_ & new_n6592_;
  assign new_n6568_ = new_n6569_ & new_n6591_;
  assign new_n6569_ = new_n6570_ & (~new_n6579_ | (new_n6589_ & new_n6590_ & new_n6586_ & new_n6588_));
  assign new_n6570_ = new_n6571_ & ~new_n6575_ & ~new_n6576_;
  assign new_n6571_ = ~new_n6572_ & (\all_features[2787]  | \all_features[2788]  | \all_features[2789]  | \all_features[2790]  | \all_features[2791] );
  assign new_n6572_ = ~\all_features[2789]  & new_n6574_ & ((~\all_features[2786]  & new_n6573_) | ~\all_features[2788]  | ~\all_features[2787] );
  assign new_n6573_ = ~\all_features[2784]  & ~\all_features[2785] ;
  assign new_n6574_ = ~\all_features[2790]  & ~\all_features[2791] ;
  assign new_n6575_ = new_n6574_ & (~\all_features[2789]  | (~\all_features[2788]  & (~\all_features[2787]  | (~\all_features[2786]  & ~\all_features[2785] ))));
  assign new_n6576_ = new_n6574_ & (~\all_features[2787]  | ~new_n6577_ | (~\all_features[2786]  & ~new_n6578_));
  assign new_n6577_ = \all_features[2788]  & \all_features[2789] ;
  assign new_n6578_ = \all_features[2784]  & \all_features[2785] ;
  assign new_n6579_ = ~new_n6585_ & ~new_n6584_ & ~new_n6580_ & ~new_n6582_;
  assign new_n6580_ = ~\all_features[2791]  & (~\all_features[2790]  | (~\all_features[2789]  & (new_n6573_ | ~new_n6581_ | ~\all_features[2788] )));
  assign new_n6581_ = \all_features[2786]  & \all_features[2787] ;
  assign new_n6582_ = ~new_n6583_ & ~\all_features[2791] ;
  assign new_n6583_ = \all_features[2789]  & \all_features[2790]  & (\all_features[2788]  | (\all_features[2786]  & \all_features[2787]  & \all_features[2785] ));
  assign new_n6584_ = ~\all_features[2791]  & (~\all_features[2790]  | ~new_n6577_ | ~new_n6578_ | ~new_n6581_);
  assign new_n6585_ = ~\all_features[2791]  & (~\all_features[2790]  | (~\all_features[2788]  & ~\all_features[2789]  & ~new_n6581_));
  assign new_n6586_ = \all_features[2791]  & (\all_features[2790]  | (\all_features[2789]  & (\all_features[2788]  | ~new_n6573_ | ~new_n6587_)));
  assign new_n6587_ = ~\all_features[2786]  & ~\all_features[2787] ;
  assign new_n6588_ = \all_features[2791]  & (\all_features[2790]  | (new_n6577_ & (\all_features[2786]  | \all_features[2787]  | \all_features[2785] )));
  assign new_n6589_ = \all_features[2790]  & \all_features[2791]  & (\all_features[2788]  | \all_features[2789]  | new_n6578_ | ~new_n6587_);
  assign new_n6590_ = \all_features[2791]  & (\all_features[2789]  | \all_features[2790]  | \all_features[2788] );
  assign new_n6591_ = new_n6570_ & new_n6579_;
  assign new_n6592_ = new_n6593_ & new_n6597_;
  assign new_n6593_ = ~new_n6594_ & (\all_features[2787]  | \all_features[2788]  | \all_features[2789]  | \all_features[2790]  | \all_features[2791] );
  assign new_n6594_ = ~new_n6572_ & (new_n6575_ | (~new_n6576_ & (new_n6585_ | (~new_n6580_ & ~new_n6595_))));
  assign new_n6595_ = ~new_n6582_ & (new_n6584_ | (new_n6590_ & (~new_n6586_ | (~new_n6596_ & new_n6588_))));
  assign new_n6596_ = ~\all_features[2789]  & \all_features[2790]  & \all_features[2791]  & (\all_features[2788]  ? new_n6587_ : (new_n6578_ | ~new_n6587_));
  assign new_n6597_ = new_n6571_ & (new_n6576_ | new_n6575_ | (~new_n6580_ & ~new_n6585_ & ~new_n6598_));
  assign new_n6598_ = ~new_n6584_ & ~new_n6582_ & (~new_n6590_ | ~new_n6586_ | new_n6599_);
  assign new_n6599_ = new_n6588_ & new_n6589_ & (new_n6600_ | ~\all_features[2789]  | ~\all_features[2790]  | ~\all_features[2791] );
  assign new_n6600_ = ~\all_features[2787]  & ~\all_features[2788]  & (~\all_features[2786]  | new_n6573_);
  assign new_n6601_ = new_n6602_ & (new_n6603_ ? new_n6638_ : new_n6674_);
  assign new_n6602_ = new_n6354_ & new_n6389_;
  assign new_n6603_ = new_n6604_ & new_n6629_;
  assign new_n6604_ = ~new_n6605_ & ~new_n6627_;
  assign new_n6605_ = new_n6622_ & ~new_n6626_ & ~new_n6606_ & ~new_n6625_;
  assign new_n6606_ = new_n6607_ & (~new_n6620_ | ~new_n6621_ | ~new_n6617_ | ~new_n6619_);
  assign new_n6607_ = ~new_n6614_ & ~new_n6613_ & ~new_n6608_ & ~new_n6611_;
  assign new_n6608_ = ~\all_features[1719]  & (~\all_features[1718]  | (~\all_features[1717]  & (new_n6609_ | ~new_n6610_ | ~\all_features[1716] )));
  assign new_n6609_ = ~\all_features[1712]  & ~\all_features[1713] ;
  assign new_n6610_ = \all_features[1714]  & \all_features[1715] ;
  assign new_n6611_ = ~new_n6612_ & ~\all_features[1719] ;
  assign new_n6612_ = \all_features[1717]  & \all_features[1718]  & (\all_features[1716]  | (\all_features[1714]  & \all_features[1715]  & \all_features[1713] ));
  assign new_n6613_ = ~\all_features[1719]  & (~\all_features[1718]  | (~\all_features[1716]  & ~\all_features[1717]  & ~new_n6610_));
  assign new_n6614_ = ~\all_features[1719]  & (~\all_features[1718]  | ~new_n6615_ | ~new_n6616_ | ~new_n6610_);
  assign new_n6615_ = \all_features[1716]  & \all_features[1717] ;
  assign new_n6616_ = \all_features[1712]  & \all_features[1713] ;
  assign new_n6617_ = \all_features[1719]  & (\all_features[1718]  | (\all_features[1717]  & (\all_features[1716]  | ~new_n6609_ | ~new_n6618_)));
  assign new_n6618_ = ~\all_features[1714]  & ~\all_features[1715] ;
  assign new_n6619_ = \all_features[1719]  & (\all_features[1718]  | (new_n6615_ & (\all_features[1714]  | \all_features[1715]  | \all_features[1713] )));
  assign new_n6620_ = \all_features[1718]  & \all_features[1719]  & (\all_features[1716]  | \all_features[1717]  | new_n6616_ | ~new_n6618_);
  assign new_n6621_ = \all_features[1719]  & (\all_features[1717]  | \all_features[1718]  | \all_features[1716] );
  assign new_n6622_ = ~new_n6623_ & (\all_features[1715]  | \all_features[1716]  | \all_features[1717]  | \all_features[1718]  | \all_features[1719] );
  assign new_n6623_ = ~\all_features[1717]  & new_n6624_ & ((~\all_features[1714]  & new_n6609_) | ~\all_features[1716]  | ~\all_features[1715] );
  assign new_n6624_ = ~\all_features[1718]  & ~\all_features[1719] ;
  assign new_n6625_ = new_n6624_ & (~\all_features[1717]  | (~\all_features[1716]  & (~\all_features[1715]  | (~\all_features[1714]  & ~\all_features[1713] ))));
  assign new_n6626_ = new_n6624_ & (~\all_features[1715]  | ~new_n6615_ | (~\all_features[1714]  & ~new_n6616_));
  assign new_n6627_ = new_n6628_ & new_n6622_ & ~new_n6611_ & ~new_n6625_;
  assign new_n6628_ = ~new_n6626_ & ~new_n6614_ & ~new_n6608_ & ~new_n6613_;
  assign new_n6629_ = ~new_n6630_ & ~new_n6634_;
  assign new_n6630_ = new_n6622_ & (new_n6626_ | new_n6625_ | (~new_n6608_ & ~new_n6613_ & ~new_n6631_));
  assign new_n6631_ = ~new_n6614_ & ~new_n6611_ & (~new_n6621_ | ~new_n6617_ | new_n6632_);
  assign new_n6632_ = new_n6619_ & new_n6620_ & (new_n6633_ | ~\all_features[1717]  | ~\all_features[1718]  | ~\all_features[1719] );
  assign new_n6633_ = ~\all_features[1715]  & ~\all_features[1716]  & (~\all_features[1714]  | new_n6609_);
  assign new_n6634_ = ~new_n6635_ & (\all_features[1715]  | \all_features[1716]  | \all_features[1717]  | \all_features[1718]  | \all_features[1719] );
  assign new_n6635_ = ~new_n6623_ & (new_n6625_ | (~new_n6626_ & (new_n6613_ | (~new_n6608_ & ~new_n6636_))));
  assign new_n6636_ = ~new_n6611_ & (new_n6614_ | (new_n6621_ & (~new_n6617_ | (~new_n6637_ & new_n6619_))));
  assign new_n6637_ = ~\all_features[1717]  & \all_features[1718]  & \all_features[1719]  & (\all_features[1716]  ? new_n6618_ : (new_n6616_ | ~new_n6618_));
  assign new_n6638_ = new_n6639_ & new_n6665_;
  assign new_n6639_ = ~new_n6640_ & ~new_n6662_;
  assign new_n6640_ = ~new_n6661_ & ~new_n6660_ & ~new_n6659_ & ~new_n6641_ & ~new_n6657_;
  assign new_n6641_ = new_n6642_ & (~new_n6655_ | ~new_n6656_ | ~new_n6652_ | ~new_n6654_);
  assign new_n6642_ = ~new_n6649_ & ~new_n6648_ & ~new_n6643_ & ~new_n6646_;
  assign new_n6643_ = ~\all_features[2583]  & (~\all_features[2582]  | (~\all_features[2581]  & (new_n6644_ | ~new_n6645_ | ~\all_features[2580] )));
  assign new_n6644_ = ~\all_features[2576]  & ~\all_features[2577] ;
  assign new_n6645_ = \all_features[2578]  & \all_features[2579] ;
  assign new_n6646_ = ~new_n6647_ & ~\all_features[2583] ;
  assign new_n6647_ = \all_features[2581]  & \all_features[2582]  & (\all_features[2580]  | (\all_features[2578]  & \all_features[2579]  & \all_features[2577] ));
  assign new_n6648_ = ~\all_features[2583]  & (~\all_features[2582]  | (~\all_features[2580]  & ~\all_features[2581]  & ~new_n6645_));
  assign new_n6649_ = ~\all_features[2583]  & (~\all_features[2582]  | ~new_n6650_ | ~new_n6651_ | ~new_n6645_);
  assign new_n6650_ = \all_features[2580]  & \all_features[2581] ;
  assign new_n6651_ = \all_features[2576]  & \all_features[2577] ;
  assign new_n6652_ = \all_features[2583]  & (\all_features[2582]  | (\all_features[2581]  & (\all_features[2580]  | ~new_n6644_ | ~new_n6653_)));
  assign new_n6653_ = ~\all_features[2578]  & ~\all_features[2579] ;
  assign new_n6654_ = \all_features[2583]  & (\all_features[2582]  | (new_n6650_ & (\all_features[2578]  | \all_features[2579]  | \all_features[2577] )));
  assign new_n6655_ = \all_features[2582]  & \all_features[2583]  & (\all_features[2580]  | \all_features[2581]  | new_n6651_ | ~new_n6653_);
  assign new_n6656_ = \all_features[2583]  & (\all_features[2581]  | \all_features[2582]  | \all_features[2580] );
  assign new_n6657_ = new_n6658_ & (~\all_features[2581]  | (~\all_features[2580]  & (~\all_features[2579]  | (~\all_features[2578]  & ~\all_features[2577] ))));
  assign new_n6658_ = ~\all_features[2582]  & ~\all_features[2583] ;
  assign new_n6659_ = ~\all_features[2581]  & new_n6658_ & ((~\all_features[2578]  & new_n6644_) | ~\all_features[2580]  | ~\all_features[2579] );
  assign new_n6660_ = new_n6658_ & (~\all_features[2579]  | ~new_n6650_ | (~\all_features[2578]  & ~new_n6651_));
  assign new_n6661_ = ~\all_features[2583]  & ~\all_features[2582]  & ~\all_features[2581]  & ~\all_features[2579]  & ~\all_features[2580] ;
  assign new_n6662_ = new_n6664_ & new_n6663_ & ~new_n6659_ & ~new_n6649_ & ~new_n6643_ & ~new_n6646_;
  assign new_n6663_ = ~new_n6648_ & ~new_n6661_;
  assign new_n6664_ = ~new_n6657_ & ~new_n6660_;
  assign new_n6665_ = ~new_n6666_ & ~new_n6670_;
  assign new_n6666_ = ~new_n6667_ & ~new_n6661_;
  assign new_n6667_ = ~new_n6659_ & (new_n6657_ | (~new_n6660_ & (new_n6648_ | (~new_n6643_ & ~new_n6668_))));
  assign new_n6668_ = ~new_n6646_ & (new_n6649_ | (new_n6656_ & (~new_n6652_ | (~new_n6669_ & new_n6654_))));
  assign new_n6669_ = ~\all_features[2581]  & \all_features[2582]  & \all_features[2583]  & (\all_features[2580]  ? new_n6653_ : (new_n6651_ | ~new_n6653_));
  assign new_n6670_ = ~new_n6659_ & ~new_n6661_ & (~new_n6664_ | (~new_n6671_ & ~new_n6643_ & ~new_n6648_));
  assign new_n6671_ = ~new_n6649_ & ~new_n6646_ & (~new_n6656_ | ~new_n6652_ | new_n6672_);
  assign new_n6672_ = new_n6654_ & new_n6655_ & (new_n6673_ | ~\all_features[2581]  | ~\all_features[2582]  | ~\all_features[2583] );
  assign new_n6673_ = ~\all_features[2579]  & ~\all_features[2580]  & (~\all_features[2578]  | new_n6644_);
  assign new_n6674_ = new_n6675_ & new_n6698_;
  assign new_n6675_ = new_n6693_ & ~new_n6697_ & ~new_n6676_ & ~new_n6696_;
  assign new_n6676_ = ~new_n6691_ & ~new_n6692_ & new_n6684_ & (~new_n6689_ | ~new_n6677_);
  assign new_n6677_ = new_n6683_ & new_n6678_ & new_n6680_;
  assign new_n6678_ = \all_features[2599]  & (\all_features[2598]  | (new_n6679_ & (\all_features[2594]  | \all_features[2595]  | \all_features[2593] )));
  assign new_n6679_ = \all_features[2596]  & \all_features[2597] ;
  assign new_n6680_ = \all_features[2598]  & \all_features[2599]  & (\all_features[2596]  | \all_features[2597]  | new_n6682_ | ~new_n6681_);
  assign new_n6681_ = ~\all_features[2594]  & ~\all_features[2595] ;
  assign new_n6682_ = \all_features[2592]  & \all_features[2593] ;
  assign new_n6683_ = \all_features[2599]  & (\all_features[2597]  | \all_features[2598]  | \all_features[2596] );
  assign new_n6684_ = ~new_n6685_ & ~new_n6687_;
  assign new_n6685_ = ~new_n6686_ & ~\all_features[2599] ;
  assign new_n6686_ = \all_features[2597]  & \all_features[2598]  & (\all_features[2596]  | (\all_features[2594]  & \all_features[2595]  & \all_features[2593] ));
  assign new_n6687_ = ~\all_features[2599]  & (~\all_features[2598]  | (~\all_features[2596]  & ~\all_features[2597]  & ~new_n6688_));
  assign new_n6688_ = \all_features[2594]  & \all_features[2595] ;
  assign new_n6689_ = \all_features[2599]  & (\all_features[2598]  | (\all_features[2597]  & (\all_features[2596]  | ~new_n6690_ | ~new_n6681_)));
  assign new_n6690_ = ~\all_features[2592]  & ~\all_features[2593] ;
  assign new_n6691_ = ~\all_features[2599]  & (~\all_features[2598]  | (~\all_features[2597]  & (new_n6690_ | ~new_n6688_ | ~\all_features[2596] )));
  assign new_n6692_ = ~\all_features[2599]  & (~\all_features[2598]  | ~new_n6679_ | ~new_n6682_ | ~new_n6688_);
  assign new_n6693_ = ~new_n6694_ & (\all_features[2595]  | \all_features[2596]  | \all_features[2597]  | \all_features[2598]  | \all_features[2599] );
  assign new_n6694_ = ~\all_features[2597]  & new_n6695_ & ((~\all_features[2594]  & new_n6690_) | ~\all_features[2596]  | ~\all_features[2595] );
  assign new_n6695_ = ~\all_features[2598]  & ~\all_features[2599] ;
  assign new_n6696_ = new_n6695_ & (~\all_features[2597]  | (~\all_features[2596]  & (~\all_features[2595]  | (~\all_features[2594]  & ~\all_features[2593] ))));
  assign new_n6697_ = new_n6695_ & (~\all_features[2595]  | ~new_n6679_ | (~\all_features[2594]  & ~new_n6682_));
  assign new_n6698_ = new_n6693_ & new_n6684_ & new_n6699_ & ~new_n6691_ & ~new_n6692_;
  assign new_n6699_ = ~new_n6696_ & ~new_n6697_;
  assign new_n6700_ = ~new_n6354_ & new_n6460_;
  assign new_n6701_ = new_n6734_ & (new_n6732_ | ~new_n6702_);
  assign new_n6702_ = ~new_n6703_ & ~new_n6723_;
  assign new_n6703_ = ~new_n6717_ & (new_n6720_ | (~new_n6722_ & (new_n6721_ | (~new_n6719_ & ~new_n6704_))));
  assign new_n6704_ = ~new_n6715_ & (new_n6711_ | (~new_n6713_ & (~new_n6716_ | new_n6705_)));
  assign new_n6705_ = \all_features[4119]  & ((~new_n6710_ & ~\all_features[4117]  & \all_features[4118] ) | (~new_n6708_ & (\all_features[4118]  | (~new_n6706_ & \all_features[4117] ))));
  assign new_n6706_ = new_n6707_ & ~\all_features[4116]  & ~\all_features[4114]  & ~\all_features[4115] ;
  assign new_n6707_ = ~\all_features[4112]  & ~\all_features[4113] ;
  assign new_n6708_ = \all_features[4119]  & (\all_features[4118]  | (new_n6709_ & (\all_features[4114]  | \all_features[4115]  | \all_features[4113] )));
  assign new_n6709_ = \all_features[4116]  & \all_features[4117] ;
  assign new_n6710_ = (~\all_features[4114]  & ~\all_features[4115]  & ~\all_features[4116]  & (~\all_features[4113]  | ~\all_features[4112] )) | (\all_features[4116]  & (\all_features[4114]  | \all_features[4115] ));
  assign new_n6711_ = ~new_n6712_ & ~\all_features[4119] ;
  assign new_n6712_ = \all_features[4117]  & \all_features[4118]  & (\all_features[4116]  | (\all_features[4114]  & \all_features[4115]  & \all_features[4113] ));
  assign new_n6713_ = ~\all_features[4119]  & (~new_n6709_ | ~\all_features[4112]  | ~\all_features[4113]  | ~\all_features[4118]  | ~new_n6714_);
  assign new_n6714_ = \all_features[4114]  & \all_features[4115] ;
  assign new_n6715_ = ~\all_features[4119]  & (~\all_features[4118]  | (~\all_features[4117]  & (new_n6707_ | ~\all_features[4116]  | ~new_n6714_)));
  assign new_n6716_ = \all_features[4119]  & (\all_features[4117]  | \all_features[4118]  | \all_features[4116] );
  assign new_n6717_ = new_n6718_ & ~\all_features[4117]  & ~\all_features[4115]  & ~\all_features[4116] ;
  assign new_n6718_ = ~\all_features[4118]  & ~\all_features[4119] ;
  assign new_n6719_ = ~\all_features[4119]  & (~\all_features[4118]  | (~\all_features[4116]  & ~\all_features[4117]  & ~new_n6714_));
  assign new_n6720_ = ~\all_features[4117]  & new_n6718_ & ((~\all_features[4114]  & new_n6707_) | ~\all_features[4116]  | ~\all_features[4115] );
  assign new_n6721_ = new_n6718_ & (~new_n6709_ | ~\all_features[4115]  | (~\all_features[4114]  & (~\all_features[4112]  | ~\all_features[4113] )));
  assign new_n6722_ = new_n6718_ & (~\all_features[4117]  | (~\all_features[4116]  & (~\all_features[4115]  | (~\all_features[4114]  & ~\all_features[4113] ))));
  assign new_n6723_ = new_n6731_ & (~new_n6730_ | (~new_n6724_ & ~new_n6719_ & ~new_n6715_));
  assign new_n6724_ = ~new_n6711_ & ~new_n6713_ & (~new_n6725_ | (~new_n6728_ & new_n6726_));
  assign new_n6725_ = \all_features[4119]  & (\all_features[4118]  | (~new_n6706_ & \all_features[4117] ));
  assign new_n6726_ = \all_features[4119]  & \all_features[4118]  & ~new_n6727_ & new_n6708_;
  assign new_n6727_ = ~\all_features[4114]  & ~\all_features[4115]  & ~\all_features[4116]  & ~\all_features[4117]  & (~\all_features[4113]  | ~\all_features[4112] );
  assign new_n6728_ = \all_features[4119]  & \all_features[4118]  & ~new_n6729_ & \all_features[4117] ;
  assign new_n6729_ = ~\all_features[4115]  & ~\all_features[4116]  & (~\all_features[4114]  | new_n6707_);
  assign new_n6730_ = ~new_n6721_ & ~new_n6722_;
  assign new_n6731_ = ~new_n6717_ & ~new_n6720_;
  assign new_n6732_ = new_n6731_ & ~new_n6733_ & new_n6730_;
  assign new_n6733_ = ~new_n6711_ & ~new_n6719_ & ~new_n6713_ & ~new_n6715_ & (~new_n6726_ | ~new_n6725_);
  assign new_n6734_ = new_n6730_ & new_n6735_ & ~new_n6715_ & ~new_n6720_ & ~new_n6711_ & ~new_n6713_;
  assign new_n6735_ = ~new_n6717_ & ~new_n6719_;
  assign new_n6736_ = new_n6737_ & new_n6766_;
  assign new_n6737_ = new_n6738_ & new_n6760_;
  assign new_n6738_ = new_n6755_ & ~new_n6759_ & ~new_n6739_ & ~new_n6758_;
  assign new_n6739_ = new_n6740_ & ~new_n6753_ & (~new_n6748_ | ~new_n6754_ | ~new_n6751_ | ~new_n6752_);
  assign new_n6740_ = ~new_n6745_ & ~new_n6741_ & ~new_n6743_;
  assign new_n6741_ = ~new_n6742_ & ~\all_features[3871] ;
  assign new_n6742_ = \all_features[3869]  & \all_features[3870]  & (\all_features[3868]  | (\all_features[3866]  & \all_features[3867]  & \all_features[3865] ));
  assign new_n6743_ = ~\all_features[3871]  & (~\all_features[3870]  | (~\all_features[3868]  & ~\all_features[3869]  & ~new_n6744_));
  assign new_n6744_ = \all_features[3866]  & \all_features[3867] ;
  assign new_n6745_ = ~\all_features[3871]  & (~\all_features[3870]  | ~new_n6746_ | ~new_n6747_ | ~new_n6744_);
  assign new_n6746_ = \all_features[3868]  & \all_features[3869] ;
  assign new_n6747_ = \all_features[3864]  & \all_features[3865] ;
  assign new_n6748_ = \all_features[3871]  & (\all_features[3870]  | (\all_features[3869]  & (\all_features[3868]  | ~new_n6750_ | ~new_n6749_)));
  assign new_n6749_ = ~\all_features[3866]  & ~\all_features[3867] ;
  assign new_n6750_ = ~\all_features[3864]  & ~\all_features[3865] ;
  assign new_n6751_ = \all_features[3871]  & (\all_features[3870]  | (new_n6746_ & (\all_features[3866]  | \all_features[3867]  | \all_features[3865] )));
  assign new_n6752_ = \all_features[3870]  & \all_features[3871]  & (\all_features[3868]  | \all_features[3869]  | new_n6747_ | ~new_n6749_);
  assign new_n6753_ = ~\all_features[3871]  & (~\all_features[3870]  | (~\all_features[3869]  & (new_n6750_ | ~new_n6744_ | ~\all_features[3868] )));
  assign new_n6754_ = \all_features[3871]  & (\all_features[3869]  | \all_features[3870]  | \all_features[3868] );
  assign new_n6755_ = ~new_n6756_ & (\all_features[3867]  | \all_features[3868]  | \all_features[3869]  | \all_features[3870]  | \all_features[3871] );
  assign new_n6756_ = new_n6757_ & (~\all_features[3867]  | ~new_n6746_ | (~\all_features[3866]  & ~new_n6747_));
  assign new_n6757_ = ~\all_features[3870]  & ~\all_features[3871] ;
  assign new_n6758_ = new_n6757_ & (~\all_features[3869]  | (~\all_features[3868]  & (~\all_features[3867]  | (~\all_features[3866]  & ~\all_features[3865] ))));
  assign new_n6759_ = ~\all_features[3869]  & new_n6757_ & ((~\all_features[3866]  & new_n6750_) | ~\all_features[3868]  | ~\all_features[3867] );
  assign new_n6760_ = new_n6765_ & (~new_n6764_ | (~new_n6761_ & ~new_n6753_ & ~new_n6743_));
  assign new_n6761_ = ~new_n6745_ & ~new_n6741_ & (~new_n6754_ | ~new_n6748_ | new_n6762_);
  assign new_n6762_ = new_n6751_ & new_n6752_ & (new_n6763_ | ~\all_features[3869]  | ~\all_features[3870]  | ~\all_features[3871] );
  assign new_n6763_ = ~\all_features[3867]  & ~\all_features[3868]  & (~\all_features[3866]  | new_n6750_);
  assign new_n6764_ = ~new_n6758_ & ~new_n6756_;
  assign new_n6765_ = ~new_n6759_ & (\all_features[3867]  | \all_features[3868]  | \all_features[3869]  | \all_features[3870]  | \all_features[3871] );
  assign new_n6766_ = new_n6740_ & new_n6765_ & ~new_n6753_ & new_n6764_;
  assign new_n6767_ = new_n6768_ & new_n6803_ & (new_n6496_ | ~new_n6459_);
  assign new_n6768_ = (~new_n6700_ | (new_n6736_ ? new_n6769_ : new_n6701_)) & (~new_n6353_ | new_n6567_);
  assign new_n6769_ = new_n6799_ & (new_n6801_ | ~new_n6770_);
  assign new_n6770_ = ~new_n6771_ & ~new_n6795_;
  assign new_n6771_ = new_n6787_ & (~new_n6790_ | (~new_n6772_ & ~new_n6793_ & ~new_n6794_));
  assign new_n6772_ = ~new_n6781_ & ~new_n6783_ & (~new_n6786_ | ~new_n6785_ | new_n6773_);
  assign new_n6773_ = new_n6774_ & new_n6776_ & (new_n6779_ | ~\all_features[5005]  | ~\all_features[5006]  | ~\all_features[5007] );
  assign new_n6774_ = \all_features[5007]  & (\all_features[5006]  | (new_n6775_ & (\all_features[5002]  | \all_features[5003]  | \all_features[5001] )));
  assign new_n6775_ = \all_features[5004]  & \all_features[5005] ;
  assign new_n6776_ = \all_features[5006]  & \all_features[5007]  & (\all_features[5004]  | \all_features[5005]  | new_n6777_ | ~new_n6778_);
  assign new_n6777_ = \all_features[5000]  & \all_features[5001] ;
  assign new_n6778_ = ~\all_features[5002]  & ~\all_features[5003] ;
  assign new_n6779_ = ~\all_features[5003]  & ~\all_features[5004]  & (~\all_features[5002]  | new_n6780_);
  assign new_n6780_ = ~\all_features[5000]  & ~\all_features[5001] ;
  assign new_n6781_ = ~new_n6782_ & ~\all_features[5007] ;
  assign new_n6782_ = \all_features[5005]  & \all_features[5006]  & (\all_features[5004]  | (\all_features[5002]  & \all_features[5003]  & \all_features[5001] ));
  assign new_n6783_ = ~\all_features[5007]  & (~\all_features[5006]  | ~new_n6784_ | ~new_n6777_ | ~new_n6775_);
  assign new_n6784_ = \all_features[5002]  & \all_features[5003] ;
  assign new_n6785_ = \all_features[5007]  & (\all_features[5006]  | (\all_features[5005]  & (\all_features[5004]  | ~new_n6778_ | ~new_n6780_)));
  assign new_n6786_ = \all_features[5007]  & (\all_features[5005]  | \all_features[5006]  | \all_features[5004] );
  assign new_n6787_ = ~new_n6788_ & (\all_features[5003]  | \all_features[5004]  | \all_features[5005]  | \all_features[5006]  | \all_features[5007] );
  assign new_n6788_ = ~\all_features[5005]  & new_n6789_ & ((~\all_features[5002]  & new_n6780_) | ~\all_features[5004]  | ~\all_features[5003] );
  assign new_n6789_ = ~\all_features[5006]  & ~\all_features[5007] ;
  assign new_n6790_ = ~new_n6791_ & ~new_n6792_;
  assign new_n6791_ = new_n6789_ & (~\all_features[5005]  | (~\all_features[5004]  & (~\all_features[5003]  | (~\all_features[5002]  & ~\all_features[5001] ))));
  assign new_n6792_ = new_n6789_ & (~\all_features[5003]  | ~new_n6775_ | (~\all_features[5002]  & ~new_n6777_));
  assign new_n6793_ = ~\all_features[5007]  & (~\all_features[5006]  | (~\all_features[5005]  & (new_n6780_ | ~new_n6784_ | ~\all_features[5004] )));
  assign new_n6794_ = ~\all_features[5007]  & (~\all_features[5006]  | (~\all_features[5004]  & ~\all_features[5005]  & ~new_n6784_));
  assign new_n6795_ = ~new_n6796_ & (\all_features[5003]  | \all_features[5004]  | \all_features[5005]  | \all_features[5006]  | \all_features[5007] );
  assign new_n6796_ = ~new_n6788_ & (new_n6791_ | (~new_n6792_ & (new_n6794_ | (~new_n6793_ & ~new_n6797_))));
  assign new_n6797_ = ~new_n6781_ & (new_n6783_ | (new_n6786_ & (~new_n6785_ | (~new_n6798_ & new_n6774_))));
  assign new_n6798_ = ~\all_features[5005]  & \all_features[5006]  & \all_features[5007]  & (\all_features[5004]  ? new_n6778_ : (new_n6777_ | ~new_n6778_));
  assign new_n6799_ = new_n6800_ & new_n6787_ & ~new_n6792_ & ~new_n6793_ & ~new_n6781_ & ~new_n6791_;
  assign new_n6800_ = ~new_n6783_ & ~new_n6794_;
  assign new_n6801_ = new_n6787_ & new_n6790_ & (new_n6802_ | new_n6781_ | new_n6793_ | ~new_n6800_);
  assign new_n6802_ = new_n6786_ & new_n6776_ & new_n6785_ & new_n6774_;
  assign new_n6803_ = ~new_n6354_ | ((new_n6638_ | ~new_n6603_ | ~new_n6389_) & (~new_n6425_ | ~new_n6804_ | new_n6389_));
  assign new_n6804_ = ~new_n6805_ & new_n6837_;
  assign new_n6805_ = new_n6806_ & new_n6833_;
  assign new_n6806_ = new_n6830_ & (~new_n6826_ | (~new_n6807_ & new_n6823_));
  assign new_n6807_ = new_n6811_ & ((~new_n6808_ & new_n6819_ & new_n6818_) | ~new_n6822_ | ~new_n6821_);
  assign new_n6808_ = \all_features[2351]  & \all_features[2350]  & ~new_n6809_ & \all_features[2349] ;
  assign new_n6809_ = ~\all_features[2347]  & ~\all_features[2348]  & (~\all_features[2346]  | new_n6810_);
  assign new_n6810_ = ~\all_features[2344]  & ~\all_features[2345] ;
  assign new_n6811_ = ~new_n6812_ & ~new_n6814_;
  assign new_n6812_ = ~new_n6813_ & ~\all_features[2351] ;
  assign new_n6813_ = \all_features[2349]  & \all_features[2350]  & (\all_features[2348]  | (\all_features[2346]  & \all_features[2347]  & \all_features[2345] ));
  assign new_n6814_ = ~\all_features[2351]  & (~\all_features[2350]  | ~new_n6815_ | ~new_n6816_ | ~new_n6817_);
  assign new_n6815_ = \all_features[2348]  & \all_features[2349] ;
  assign new_n6816_ = \all_features[2344]  & \all_features[2345] ;
  assign new_n6817_ = \all_features[2346]  & \all_features[2347] ;
  assign new_n6818_ = \all_features[2351]  & (\all_features[2350]  | (new_n6815_ & (\all_features[2346]  | \all_features[2347]  | \all_features[2345] )));
  assign new_n6819_ = \all_features[2350]  & \all_features[2351]  & (\all_features[2348]  | \all_features[2349]  | new_n6816_ | ~new_n6820_);
  assign new_n6820_ = ~\all_features[2346]  & ~\all_features[2347] ;
  assign new_n6821_ = \all_features[2351]  & (\all_features[2350]  | (\all_features[2349]  & (\all_features[2348]  | ~new_n6820_ | ~new_n6810_)));
  assign new_n6822_ = \all_features[2351]  & (\all_features[2349]  | \all_features[2350]  | \all_features[2348] );
  assign new_n6823_ = ~new_n6824_ & ~new_n6825_;
  assign new_n6824_ = ~\all_features[2351]  & (~\all_features[2350]  | (~\all_features[2348]  & ~\all_features[2349]  & ~new_n6817_));
  assign new_n6825_ = ~\all_features[2351]  & (~\all_features[2350]  | (~\all_features[2349]  & (new_n6810_ | ~new_n6817_ | ~\all_features[2348] )));
  assign new_n6826_ = ~new_n6827_ & ~new_n6829_;
  assign new_n6827_ = new_n6828_ & (~\all_features[2349]  | (~\all_features[2348]  & (~\all_features[2347]  | (~\all_features[2346]  & ~\all_features[2345] ))));
  assign new_n6828_ = ~\all_features[2350]  & ~\all_features[2351] ;
  assign new_n6829_ = new_n6828_ & (~\all_features[2347]  | ~new_n6815_ | (~\all_features[2346]  & ~new_n6816_));
  assign new_n6830_ = ~new_n6831_ & ~new_n6832_;
  assign new_n6831_ = ~\all_features[2349]  & new_n6828_ & ((~\all_features[2346]  & new_n6810_) | ~\all_features[2348]  | ~\all_features[2347] );
  assign new_n6832_ = ~\all_features[2351]  & ~\all_features[2350]  & ~\all_features[2349]  & ~\all_features[2347]  & ~\all_features[2348] ;
  assign new_n6833_ = ~new_n6832_ & (new_n6831_ | new_n6834_);
  assign new_n6834_ = ~new_n6827_ & (new_n6829_ | (~new_n6824_ & (new_n6825_ | (~new_n6812_ & ~new_n6835_))));
  assign new_n6835_ = ~new_n6814_ & (~new_n6822_ | (new_n6821_ & (~new_n6818_ | (~new_n6836_ & new_n6819_))));
  assign new_n6836_ = \all_features[2350]  & \all_features[2351]  & (\all_features[2349]  | (~new_n6820_ & \all_features[2348] ));
  assign new_n6837_ = ~new_n6838_ & ~new_n6841_;
  assign new_n6838_ = new_n6840_ & (~new_n6839_ | (new_n6821_ & new_n6822_ & new_n6818_ & new_n6819_));
  assign new_n6839_ = new_n6811_ & new_n6823_;
  assign new_n6840_ = new_n6826_ & new_n6830_;
  assign new_n6841_ = new_n6839_ & new_n6840_;
  assign new_n6842_ = (~new_n6736_ | ~new_n6769_ | ~new_n6700_) & (new_n6603_ | new_n6674_ | ~new_n6602_);
  assign new_n6843_ = new_n6844_ & (~new_n7161_ | ~new_n7162_ | ~new_n7223_ | ~new_n7064_);
  assign new_n6844_ = ~new_n7065_ & new_n6845_ & (~new_n7064_ | (new_n7161_ & new_n7162_) | (new_n7193_ & ~new_n7162_));
  assign new_n6845_ = (~new_n6918_ | ~new_n6846_) & (new_n7002_ | new_n7040_ | ~new_n6972_);
  assign new_n6846_ = new_n6847_ & new_n6884_;
  assign new_n6847_ = new_n6848_ & new_n6879_;
  assign new_n6848_ = ~new_n6849_ & ~new_n6869_;
  assign new_n6849_ = (new_n6850_ | (new_n6868_ & (~\all_features[3035]  | ~\all_features[3036]  | (~\all_features[3034]  & new_n6854_)))) & (~new_n6868_ | \all_features[3035]  | \all_features[3036] );
  assign new_n6850_ = ~new_n6861_ & (new_n6863_ | (~new_n6864_ & (new_n6865_ | (~new_n6851_ & ~new_n6866_))));
  assign new_n6851_ = ~new_n6859_ & (~\all_features[3039]  | new_n6852_ | (~\all_features[3036]  & ~\all_features[3037]  & ~\all_features[3038] ));
  assign new_n6852_ = \all_features[3039]  & ((~new_n6855_ & ~\all_features[3037]  & \all_features[3038] ) | (~new_n6857_ & (\all_features[3038]  | (~new_n6853_ & \all_features[3037] ))));
  assign new_n6853_ = new_n6854_ & ~\all_features[3036]  & ~\all_features[3034]  & ~\all_features[3035] ;
  assign new_n6854_ = ~\all_features[3032]  & ~\all_features[3033] ;
  assign new_n6855_ = (\all_features[3036]  & (\all_features[3034]  | \all_features[3035] )) | (~new_n6856_ & ~\all_features[3034]  & ~\all_features[3035]  & ~\all_features[3036] );
  assign new_n6856_ = \all_features[3032]  & \all_features[3033] ;
  assign new_n6857_ = \all_features[3039]  & (\all_features[3038]  | (new_n6858_ & (\all_features[3034]  | \all_features[3035]  | \all_features[3033] )));
  assign new_n6858_ = \all_features[3036]  & \all_features[3037] ;
  assign new_n6859_ = ~\all_features[3039]  & (~\all_features[3038]  | ~new_n6856_ | ~new_n6858_ | ~new_n6860_);
  assign new_n6860_ = \all_features[3034]  & \all_features[3035] ;
  assign new_n6861_ = ~\all_features[3039]  & ~new_n6862_ & ~\all_features[3038] ;
  assign new_n6862_ = \all_features[3037]  & (\all_features[3036]  | (\all_features[3035]  & (\all_features[3034]  | \all_features[3033] )));
  assign new_n6863_ = ~\all_features[3038]  & ~\all_features[3039]  & (~\all_features[3035]  | ~new_n6858_ | (~\all_features[3034]  & ~new_n6856_));
  assign new_n6864_ = ~\all_features[3039]  & (~\all_features[3038]  | (~\all_features[3036]  & ~\all_features[3037]  & ~new_n6860_));
  assign new_n6865_ = ~\all_features[3039]  & (~\all_features[3038]  | (~\all_features[3037]  & (new_n6854_ | ~new_n6860_ | ~\all_features[3036] )));
  assign new_n6866_ = ~new_n6867_ & ~\all_features[3039] ;
  assign new_n6867_ = \all_features[3037]  & \all_features[3038]  & (\all_features[3036]  | (\all_features[3034]  & \all_features[3035]  & \all_features[3033] ));
  assign new_n6868_ = ~\all_features[3039]  & ~\all_features[3037]  & ~\all_features[3038] ;
  assign new_n6869_ = new_n6878_ & (~new_n6875_ | (new_n6876_ & (~new_n6877_ | new_n6870_)));
  assign new_n6870_ = new_n6871_ & (~new_n6872_ | (~new_n6874_ & \all_features[3037]  & \all_features[3038]  & \all_features[3039] ));
  assign new_n6871_ = \all_features[3039]  & (\all_features[3038]  | (~new_n6853_ & \all_features[3037] ));
  assign new_n6872_ = \all_features[3039]  & \all_features[3038]  & ~new_n6873_ & new_n6857_;
  assign new_n6873_ = ~\all_features[3037]  & ~\all_features[3036]  & ~\all_features[3035]  & ~new_n6856_ & ~\all_features[3034] ;
  assign new_n6874_ = ~\all_features[3035]  & ~\all_features[3036]  & (~\all_features[3034]  | new_n6854_);
  assign new_n6875_ = ~new_n6861_ & ~new_n6863_;
  assign new_n6876_ = ~new_n6864_ & ~new_n6865_;
  assign new_n6877_ = ~new_n6866_ & ~new_n6859_;
  assign new_n6878_ = ~new_n6868_ | (\all_features[3035]  & \all_features[3036]  & (\all_features[3034]  | ~new_n6854_));
  assign new_n6879_ = ~new_n6880_ & ~new_n6883_;
  assign new_n6880_ = new_n6881_ & (new_n6865_ | new_n6866_ | ~new_n6882_ | (new_n6872_ & new_n6871_));
  assign new_n6881_ = new_n6875_ & new_n6878_;
  assign new_n6882_ = ~new_n6864_ & ~new_n6859_;
  assign new_n6883_ = new_n6877_ & new_n6881_ & new_n6876_;
  assign new_n6884_ = new_n6885_ & new_n6909_;
  assign new_n6885_ = ~new_n6886_ & ~new_n6908_;
  assign new_n6886_ = new_n6887_ & (~new_n6896_ | (new_n6906_ & new_n6907_ & new_n6903_ & new_n6905_));
  assign new_n6887_ = new_n6888_ & ~new_n6892_ & ~new_n6893_;
  assign new_n6888_ = ~new_n6889_ & (\all_features[3475]  | \all_features[3476]  | \all_features[3477]  | \all_features[3478]  | \all_features[3479] );
  assign new_n6889_ = ~\all_features[3477]  & new_n6891_ & ((~\all_features[3474]  & new_n6890_) | ~\all_features[3476]  | ~\all_features[3475] );
  assign new_n6890_ = ~\all_features[3472]  & ~\all_features[3473] ;
  assign new_n6891_ = ~\all_features[3478]  & ~\all_features[3479] ;
  assign new_n6892_ = new_n6891_ & (~\all_features[3477]  | (~\all_features[3476]  & (~\all_features[3475]  | (~\all_features[3474]  & ~\all_features[3473] ))));
  assign new_n6893_ = new_n6891_ & (~\all_features[3475]  | ~new_n6894_ | (~\all_features[3474]  & ~new_n6895_));
  assign new_n6894_ = \all_features[3476]  & \all_features[3477] ;
  assign new_n6895_ = \all_features[3472]  & \all_features[3473] ;
  assign new_n6896_ = ~new_n6902_ & ~new_n6901_ & ~new_n6897_ & ~new_n6899_;
  assign new_n6897_ = ~\all_features[3479]  & (~\all_features[3478]  | (~\all_features[3477]  & (new_n6890_ | ~new_n6898_ | ~\all_features[3476] )));
  assign new_n6898_ = \all_features[3474]  & \all_features[3475] ;
  assign new_n6899_ = ~new_n6900_ & ~\all_features[3479] ;
  assign new_n6900_ = \all_features[3477]  & \all_features[3478]  & (\all_features[3476]  | (\all_features[3474]  & \all_features[3475]  & \all_features[3473] ));
  assign new_n6901_ = ~\all_features[3479]  & (~\all_features[3478]  | ~new_n6894_ | ~new_n6895_ | ~new_n6898_);
  assign new_n6902_ = ~\all_features[3479]  & (~\all_features[3478]  | (~\all_features[3476]  & ~\all_features[3477]  & ~new_n6898_));
  assign new_n6903_ = \all_features[3479]  & (\all_features[3478]  | (\all_features[3477]  & (\all_features[3476]  | ~new_n6890_ | ~new_n6904_)));
  assign new_n6904_ = ~\all_features[3474]  & ~\all_features[3475] ;
  assign new_n6905_ = \all_features[3479]  & (\all_features[3478]  | (new_n6894_ & (\all_features[3474]  | \all_features[3475]  | \all_features[3473] )));
  assign new_n6906_ = \all_features[3478]  & \all_features[3479]  & (\all_features[3476]  | \all_features[3477]  | new_n6895_ | ~new_n6904_);
  assign new_n6907_ = \all_features[3479]  & (\all_features[3477]  | \all_features[3478]  | \all_features[3476] );
  assign new_n6908_ = new_n6887_ & new_n6896_;
  assign new_n6909_ = ~new_n6910_ & ~new_n6914_;
  assign new_n6910_ = new_n6888_ & (new_n6893_ | new_n6892_ | (~new_n6897_ & ~new_n6902_ & ~new_n6911_));
  assign new_n6911_ = ~new_n6901_ & ~new_n6899_ & (~new_n6907_ | ~new_n6903_ | new_n6912_);
  assign new_n6912_ = new_n6905_ & new_n6906_ & (new_n6913_ | ~\all_features[3477]  | ~\all_features[3478]  | ~\all_features[3479] );
  assign new_n6913_ = ~\all_features[3475]  & ~\all_features[3476]  & (~\all_features[3474]  | new_n6890_);
  assign new_n6914_ = ~new_n6915_ & (\all_features[3475]  | \all_features[3476]  | \all_features[3477]  | \all_features[3478]  | \all_features[3479] );
  assign new_n6915_ = ~new_n6889_ & (new_n6892_ | (~new_n6893_ & (new_n6902_ | (~new_n6897_ & ~new_n6916_))));
  assign new_n6916_ = ~new_n6899_ & (new_n6901_ | (new_n6907_ & (~new_n6903_ | (~new_n6917_ & new_n6905_))));
  assign new_n6917_ = ~\all_features[3477]  & \all_features[3478]  & \all_features[3479]  & (\all_features[3476]  ? new_n6904_ : (new_n6895_ | ~new_n6904_));
  assign new_n6918_ = new_n6919_ & new_n6955_;
  assign new_n6919_ = new_n6920_ & new_n6949_;
  assign new_n6920_ = ~new_n6921_ & ~new_n6945_;
  assign new_n6921_ = new_n6936_ & (~new_n6941_ | (~new_n6939_ & ~new_n6922_ & ~new_n6944_));
  assign new_n6922_ = ~new_n6934_ & ~new_n6932_ & (~new_n6935_ | ~new_n6931_ | new_n6923_);
  assign new_n6923_ = new_n6924_ & new_n6926_ & (new_n6929_ | ~\all_features[3213]  | ~\all_features[3214]  | ~\all_features[3215] );
  assign new_n6924_ = \all_features[3215]  & (\all_features[3214]  | (new_n6925_ & (\all_features[3210]  | \all_features[3211]  | \all_features[3209] )));
  assign new_n6925_ = \all_features[3212]  & \all_features[3213] ;
  assign new_n6926_ = \all_features[3214]  & \all_features[3215]  & (\all_features[3212]  | \all_features[3213]  | new_n6928_ | ~new_n6927_);
  assign new_n6927_ = ~\all_features[3210]  & ~\all_features[3211] ;
  assign new_n6928_ = \all_features[3208]  & \all_features[3209] ;
  assign new_n6929_ = ~\all_features[3211]  & ~\all_features[3212]  & (~\all_features[3210]  | new_n6930_);
  assign new_n6930_ = ~\all_features[3208]  & ~\all_features[3209] ;
  assign new_n6931_ = \all_features[3215]  & (\all_features[3214]  | (\all_features[3213]  & (\all_features[3212]  | ~new_n6927_ | ~new_n6930_)));
  assign new_n6932_ = ~new_n6933_ & ~\all_features[3215] ;
  assign new_n6933_ = \all_features[3213]  & \all_features[3214]  & (\all_features[3212]  | (\all_features[3210]  & \all_features[3211]  & \all_features[3209] ));
  assign new_n6934_ = ~\all_features[3215]  & (~new_n6928_ | ~\all_features[3210]  | ~\all_features[3211]  | ~\all_features[3214]  | ~new_n6925_);
  assign new_n6935_ = \all_features[3215]  & (\all_features[3213]  | \all_features[3214]  | \all_features[3212] );
  assign new_n6936_ = ~new_n6937_ & (\all_features[3211]  | \all_features[3212]  | \all_features[3213]  | \all_features[3214]  | \all_features[3215] );
  assign new_n6937_ = ~\all_features[3213]  & new_n6938_ & ((~\all_features[3210]  & new_n6930_) | ~\all_features[3212]  | ~\all_features[3211] );
  assign new_n6938_ = ~\all_features[3214]  & ~\all_features[3215] ;
  assign new_n6939_ = ~\all_features[3215]  & (~\all_features[3214]  | new_n6940_);
  assign new_n6940_ = ~\all_features[3213]  & (new_n6930_ | ~\all_features[3211]  | ~\all_features[3212]  | ~\all_features[3210] );
  assign new_n6941_ = ~new_n6942_ & ~new_n6943_;
  assign new_n6942_ = new_n6938_ & (~\all_features[3213]  | (~\all_features[3212]  & (~\all_features[3211]  | (~\all_features[3210]  & ~\all_features[3209] ))));
  assign new_n6943_ = new_n6938_ & (~\all_features[3211]  | ~new_n6925_ | (~new_n6928_ & ~\all_features[3210] ));
  assign new_n6944_ = ~\all_features[3215]  & (~\all_features[3214]  | (~\all_features[3213]  & ~\all_features[3212]  & (~\all_features[3211]  | ~\all_features[3210] )));
  assign new_n6945_ = ~new_n6946_ & (\all_features[3211]  | \all_features[3212]  | \all_features[3213]  | \all_features[3214]  | \all_features[3215] );
  assign new_n6946_ = ~new_n6937_ & (new_n6942_ | (~new_n6943_ & (new_n6944_ | (~new_n6939_ & ~new_n6947_))));
  assign new_n6947_ = ~new_n6932_ & (new_n6934_ | (new_n6935_ & (~new_n6931_ | (~new_n6948_ & new_n6924_))));
  assign new_n6948_ = ~\all_features[3213]  & \all_features[3214]  & \all_features[3215]  & (\all_features[3212]  ? new_n6927_ : (new_n6928_ | ~new_n6927_));
  assign new_n6949_ = ~new_n6950_ & ~new_n6953_;
  assign new_n6950_ = new_n6941_ & ~new_n6951_ & new_n6936_;
  assign new_n6951_ = ~new_n6944_ & ~new_n6934_ & ~new_n6932_ & ~new_n6939_ & ~new_n6952_;
  assign new_n6952_ = new_n6935_ & new_n6931_ & new_n6924_ & new_n6926_;
  assign new_n6953_ = new_n6936_ & new_n6954_ & ~new_n6932_ & ~new_n6942_;
  assign new_n6954_ = ~new_n6944_ & ~new_n6943_ & ~new_n6939_ & ~new_n6934_;
  assign new_n6955_ = new_n6961_ & new_n6956_ & new_n6967_ & ~new_n6969_ & ~new_n6971_;
  assign new_n6956_ = ~new_n6957_ & ~new_n6959_;
  assign new_n6957_ = ~\all_features[4151]  & (~\all_features[4150]  | (~\all_features[4148]  & ~\all_features[4149]  & ~new_n6958_));
  assign new_n6958_ = \all_features[4146]  & \all_features[4147] ;
  assign new_n6959_ = ~\all_features[4151]  & (~\all_features[4150]  | (~\all_features[4149]  & (new_n6960_ | ~\all_features[4148]  | ~new_n6958_)));
  assign new_n6960_ = ~\all_features[4144]  & ~\all_features[4145] ;
  assign new_n6961_ = ~new_n6962_ & ~new_n6966_;
  assign new_n6962_ = new_n6963_ & (~\all_features[4147]  | ~new_n6965_ | (~\all_features[4146]  & ~new_n6964_));
  assign new_n6963_ = ~\all_features[4150]  & ~\all_features[4151] ;
  assign new_n6964_ = \all_features[4144]  & \all_features[4145] ;
  assign new_n6965_ = \all_features[4148]  & \all_features[4149] ;
  assign new_n6966_ = new_n6963_ & (~\all_features[4149]  | (~\all_features[4148]  & (~\all_features[4147]  | (~\all_features[4146]  & ~\all_features[4145] ))));
  assign new_n6967_ = ~new_n6968_ & (\all_features[4147]  | \all_features[4148]  | \all_features[4149]  | \all_features[4150]  | \all_features[4151] );
  assign new_n6968_ = ~\all_features[4151]  & (~\all_features[4150]  | ~new_n6958_ | ~new_n6964_ | ~new_n6965_);
  assign new_n6969_ = ~new_n6970_ & ~\all_features[4151] ;
  assign new_n6970_ = \all_features[4149]  & \all_features[4150]  & (\all_features[4148]  | (\all_features[4146]  & \all_features[4147]  & \all_features[4145] ));
  assign new_n6971_ = ~\all_features[4149]  & new_n6963_ & ((~\all_features[4146]  & new_n6960_) | ~\all_features[4148]  | ~\all_features[4147] );
  assign new_n6972_ = ~new_n6884_ & new_n6973_;
  assign new_n6973_ = ~new_n6998_ & (~new_n7000_ | ~new_n6974_);
  assign new_n6974_ = new_n6990_ & (~new_n6993_ | (~new_n6975_ & ~new_n6996_ & ~new_n6997_));
  assign new_n6975_ = ~new_n6984_ & ~new_n6986_ & (~new_n6989_ | ~new_n6988_ | new_n6976_);
  assign new_n6976_ = new_n6977_ & new_n6979_ & (new_n6982_ | ~\all_features[3093]  | ~\all_features[3094]  | ~\all_features[3095] );
  assign new_n6977_ = \all_features[3095]  & (\all_features[3094]  | (new_n6978_ & (\all_features[3090]  | \all_features[3091]  | \all_features[3089] )));
  assign new_n6978_ = \all_features[3092]  & \all_features[3093] ;
  assign new_n6979_ = \all_features[3094]  & \all_features[3095]  & (\all_features[3092]  | \all_features[3093]  | new_n6980_ | ~new_n6981_);
  assign new_n6980_ = \all_features[3088]  & \all_features[3089] ;
  assign new_n6981_ = ~\all_features[3090]  & ~\all_features[3091] ;
  assign new_n6982_ = ~\all_features[3091]  & ~\all_features[3092]  & (~\all_features[3090]  | new_n6983_);
  assign new_n6983_ = ~\all_features[3088]  & ~\all_features[3089] ;
  assign new_n6984_ = ~new_n6985_ & ~\all_features[3095] ;
  assign new_n6985_ = \all_features[3093]  & \all_features[3094]  & (\all_features[3092]  | (\all_features[3090]  & \all_features[3091]  & \all_features[3089] ));
  assign new_n6986_ = ~\all_features[3095]  & (~\all_features[3094]  | ~new_n6987_ | ~new_n6980_ | ~new_n6978_);
  assign new_n6987_ = \all_features[3090]  & \all_features[3091] ;
  assign new_n6988_ = \all_features[3095]  & (\all_features[3094]  | (\all_features[3093]  & (\all_features[3092]  | ~new_n6981_ | ~new_n6983_)));
  assign new_n6989_ = \all_features[3095]  & (\all_features[3093]  | \all_features[3094]  | \all_features[3092] );
  assign new_n6990_ = ~new_n6991_ & (\all_features[3091]  | \all_features[3092]  | \all_features[3093]  | \all_features[3094]  | \all_features[3095] );
  assign new_n6991_ = ~\all_features[3093]  & new_n6992_ & ((~\all_features[3090]  & new_n6983_) | ~\all_features[3092]  | ~\all_features[3091] );
  assign new_n6992_ = ~\all_features[3094]  & ~\all_features[3095] ;
  assign new_n6993_ = ~new_n6994_ & ~new_n6995_;
  assign new_n6994_ = new_n6992_ & (~\all_features[3093]  | (~\all_features[3092]  & (~\all_features[3091]  | (~\all_features[3090]  & ~\all_features[3089] ))));
  assign new_n6995_ = new_n6992_ & (~\all_features[3091]  | ~new_n6978_ | (~\all_features[3090]  & ~new_n6980_));
  assign new_n6996_ = ~\all_features[3095]  & (~\all_features[3094]  | (~\all_features[3093]  & (new_n6983_ | ~new_n6987_ | ~\all_features[3092] )));
  assign new_n6997_ = ~\all_features[3095]  & (~\all_features[3094]  | (~\all_features[3092]  & ~\all_features[3093]  & ~new_n6987_));
  assign new_n6998_ = new_n6999_ & new_n6990_ & ~new_n6995_ & ~new_n6996_ & ~new_n6984_ & ~new_n6994_;
  assign new_n6999_ = ~new_n6986_ & ~new_n6997_;
  assign new_n7000_ = new_n6990_ & new_n6993_ & (new_n7001_ | new_n6984_ | new_n6996_ | ~new_n6999_);
  assign new_n7001_ = new_n6989_ & new_n6988_ & new_n6977_ & new_n6979_;
  assign new_n7002_ = new_n7003_ & new_n7035_;
  assign new_n7003_ = new_n7004_ & new_n7025_;
  assign new_n7004_ = ~new_n7005_ & (\all_features[2883]  | \all_features[2884]  | \all_features[2885]  | \all_features[2886]  | \all_features[2887] );
  assign new_n7005_ = ~new_n7019_ & (new_n7021_ | (~new_n7022_ & (new_n7023_ | (~new_n7006_ & ~new_n7024_))));
  assign new_n7006_ = ~new_n7014_ & (new_n7016_ | (~new_n7007_ & new_n7018_));
  assign new_n7007_ = \all_features[2887]  & ((~new_n7012_ & ~\all_features[2885]  & \all_features[2886] ) | (~new_n7010_ & (\all_features[2886]  | (~new_n7008_ & \all_features[2885] ))));
  assign new_n7008_ = new_n7009_ & ~\all_features[2884]  & ~\all_features[2882]  & ~\all_features[2883] ;
  assign new_n7009_ = ~\all_features[2880]  & ~\all_features[2881] ;
  assign new_n7010_ = \all_features[2887]  & (\all_features[2886]  | (new_n7011_ & (\all_features[2882]  | \all_features[2883]  | \all_features[2881] )));
  assign new_n7011_ = \all_features[2884]  & \all_features[2885] ;
  assign new_n7012_ = (\all_features[2884]  & (\all_features[2882]  | \all_features[2883] )) | (~new_n7013_ & ~\all_features[2882]  & ~\all_features[2883]  & ~\all_features[2884] );
  assign new_n7013_ = \all_features[2880]  & \all_features[2881] ;
  assign new_n7014_ = ~new_n7015_ & ~\all_features[2887] ;
  assign new_n7015_ = \all_features[2885]  & \all_features[2886]  & (\all_features[2884]  | (\all_features[2882]  & \all_features[2883]  & \all_features[2881] ));
  assign new_n7016_ = ~\all_features[2887]  & (~\all_features[2886]  | ~new_n7013_ | ~new_n7011_ | ~new_n7017_);
  assign new_n7017_ = \all_features[2882]  & \all_features[2883] ;
  assign new_n7018_ = \all_features[2887]  & (\all_features[2885]  | \all_features[2886]  | \all_features[2884] );
  assign new_n7019_ = ~\all_features[2885]  & new_n7020_ & ((~\all_features[2882]  & new_n7009_) | ~\all_features[2884]  | ~\all_features[2883] );
  assign new_n7020_ = ~\all_features[2886]  & ~\all_features[2887] ;
  assign new_n7021_ = new_n7020_ & (~\all_features[2885]  | (~\all_features[2884]  & (~\all_features[2883]  | (~\all_features[2882]  & ~\all_features[2881] ))));
  assign new_n7022_ = new_n7020_ & (~\all_features[2883]  | ~new_n7011_ | (~\all_features[2882]  & ~new_n7013_));
  assign new_n7023_ = ~\all_features[2887]  & (~\all_features[2886]  | (~\all_features[2884]  & ~\all_features[2885]  & ~new_n7017_));
  assign new_n7024_ = ~\all_features[2887]  & (~\all_features[2886]  | (~\all_features[2885]  & (new_n7009_ | ~new_n7017_ | ~\all_features[2884] )));
  assign new_n7025_ = new_n7031_ & (~new_n7032_ | (new_n7033_ & (~new_n7034_ | new_n7026_)));
  assign new_n7026_ = new_n7027_ & (~new_n7028_ | (~new_n7030_ & \all_features[2885]  & \all_features[2886]  & \all_features[2887] ));
  assign new_n7027_ = \all_features[2887]  & (\all_features[2886]  | (~new_n7008_ & \all_features[2885] ));
  assign new_n7028_ = \all_features[2887]  & \all_features[2886]  & ~new_n7029_ & new_n7010_;
  assign new_n7029_ = ~\all_features[2885]  & ~\all_features[2884]  & ~\all_features[2883]  & ~new_n7013_ & ~\all_features[2882] ;
  assign new_n7030_ = ~\all_features[2883]  & ~\all_features[2884]  & (~\all_features[2882]  | new_n7009_);
  assign new_n7031_ = ~new_n7019_ & (\all_features[2883]  | \all_features[2884]  | \all_features[2885]  | \all_features[2886]  | \all_features[2887] );
  assign new_n7032_ = ~new_n7021_ & ~new_n7022_;
  assign new_n7033_ = ~new_n7023_ & ~new_n7024_;
  assign new_n7034_ = ~new_n7014_ & ~new_n7016_;
  assign new_n7035_ = new_n7036_ & new_n7039_;
  assign new_n7036_ = new_n7037_ & (new_n7024_ | new_n7014_ | ~new_n7038_ | (new_n7028_ & new_n7027_));
  assign new_n7037_ = new_n7031_ & new_n7032_;
  assign new_n7038_ = ~new_n7023_ & ~new_n7016_;
  assign new_n7039_ = new_n7034_ & new_n7037_ & new_n7033_;
  assign new_n7040_ = new_n7041_ & new_n7063_;
  assign new_n7041_ = new_n7042_ & (~new_n7051_ | (new_n7061_ & new_n7062_ & new_n7058_ & new_n7060_));
  assign new_n7042_ = new_n7043_ & ~new_n7047_ & ~new_n7048_;
  assign new_n7043_ = ~new_n7044_ & (\all_features[3075]  | \all_features[3076]  | \all_features[3077]  | \all_features[3078]  | \all_features[3079] );
  assign new_n7044_ = ~\all_features[3077]  & new_n7046_ & ((~\all_features[3074]  & new_n7045_) | ~\all_features[3076]  | ~\all_features[3075] );
  assign new_n7045_ = ~\all_features[3072]  & ~\all_features[3073] ;
  assign new_n7046_ = ~\all_features[3078]  & ~\all_features[3079] ;
  assign new_n7047_ = new_n7046_ & (~\all_features[3077]  | (~\all_features[3076]  & (~\all_features[3075]  | (~\all_features[3074]  & ~\all_features[3073] ))));
  assign new_n7048_ = new_n7046_ & (~\all_features[3075]  | ~new_n7049_ | (~\all_features[3074]  & ~new_n7050_));
  assign new_n7049_ = \all_features[3076]  & \all_features[3077] ;
  assign new_n7050_ = \all_features[3072]  & \all_features[3073] ;
  assign new_n7051_ = ~new_n7057_ & ~new_n7056_ & ~new_n7052_ & ~new_n7054_;
  assign new_n7052_ = ~\all_features[3079]  & (~\all_features[3078]  | (~\all_features[3077]  & (new_n7045_ | ~new_n7053_ | ~\all_features[3076] )));
  assign new_n7053_ = \all_features[3074]  & \all_features[3075] ;
  assign new_n7054_ = ~new_n7055_ & ~\all_features[3079] ;
  assign new_n7055_ = \all_features[3077]  & \all_features[3078]  & (\all_features[3076]  | (\all_features[3074]  & \all_features[3075]  & \all_features[3073] ));
  assign new_n7056_ = ~\all_features[3079]  & (~\all_features[3078]  | ~new_n7049_ | ~new_n7050_ | ~new_n7053_);
  assign new_n7057_ = ~\all_features[3079]  & (~\all_features[3078]  | (~\all_features[3076]  & ~\all_features[3077]  & ~new_n7053_));
  assign new_n7058_ = \all_features[3079]  & (\all_features[3078]  | (\all_features[3077]  & (\all_features[3076]  | ~new_n7045_ | ~new_n7059_)));
  assign new_n7059_ = ~\all_features[3074]  & ~\all_features[3075] ;
  assign new_n7060_ = \all_features[3079]  & (\all_features[3078]  | (new_n7049_ & (\all_features[3074]  | \all_features[3075]  | \all_features[3073] )));
  assign new_n7061_ = \all_features[3078]  & \all_features[3079]  & (\all_features[3076]  | \all_features[3077]  | new_n7050_ | ~new_n7059_);
  assign new_n7062_ = \all_features[3079]  & (\all_features[3077]  | \all_features[3078]  | \all_features[3076] );
  assign new_n7063_ = new_n7042_ & new_n7051_;
  assign new_n7064_ = ~new_n6847_ & new_n6884_;
  assign new_n7065_ = ~new_n6884_ & ((~new_n7136_ & new_n7040_ & new_n6973_) | (~new_n7066_ & ~new_n7102_ & ~new_n6973_));
  assign new_n7066_ = ~new_n7067_ & new_n7097_;
  assign new_n7067_ = new_n7068_ & new_n7089_;
  assign new_n7068_ = ~new_n7069_ & (\all_features[3051]  | \all_features[3052]  | \all_features[3053]  | \all_features[3054]  | \all_features[3055] );
  assign new_n7069_ = ~new_n7083_ & (new_n7088_ | (~new_n7085_ & (new_n7086_ | (~new_n7087_ & ~new_n7070_))));
  assign new_n7070_ = ~new_n7071_ & (new_n7080_ | (new_n7082_ & (~new_n7073_ | (~new_n7078_ & new_n7076_))));
  assign new_n7071_ = ~new_n7072_ & ~\all_features[3055] ;
  assign new_n7072_ = \all_features[3053]  & \all_features[3054]  & (\all_features[3052]  | (\all_features[3050]  & \all_features[3051]  & \all_features[3049] ));
  assign new_n7073_ = \all_features[3055]  & (\all_features[3054]  | (\all_features[3053]  & (\all_features[3052]  | ~new_n7075_ | ~new_n7074_)));
  assign new_n7074_ = ~\all_features[3048]  & ~\all_features[3049] ;
  assign new_n7075_ = ~\all_features[3050]  & ~\all_features[3051] ;
  assign new_n7076_ = \all_features[3055]  & (\all_features[3054]  | (new_n7077_ & (\all_features[3050]  | \all_features[3051]  | \all_features[3049] )));
  assign new_n7077_ = \all_features[3052]  & \all_features[3053] ;
  assign new_n7078_ = ~\all_features[3053]  & \all_features[3054]  & \all_features[3055]  & (\all_features[3052]  ? new_n7075_ : (new_n7079_ | ~new_n7075_));
  assign new_n7079_ = \all_features[3048]  & \all_features[3049] ;
  assign new_n7080_ = ~\all_features[3055]  & (~\all_features[3054]  | ~new_n7079_ | ~new_n7077_ | ~new_n7081_);
  assign new_n7081_ = \all_features[3050]  & \all_features[3051] ;
  assign new_n7082_ = \all_features[3055]  & (\all_features[3053]  | \all_features[3054]  | \all_features[3052] );
  assign new_n7083_ = ~\all_features[3053]  & new_n7084_ & ((~\all_features[3050]  & new_n7074_) | ~\all_features[3052]  | ~\all_features[3051] );
  assign new_n7084_ = ~\all_features[3054]  & ~\all_features[3055] ;
  assign new_n7085_ = new_n7084_ & (~\all_features[3051]  | ~new_n7077_ | (~\all_features[3050]  & ~new_n7079_));
  assign new_n7086_ = ~\all_features[3055]  & (~\all_features[3054]  | (~\all_features[3052]  & ~\all_features[3053]  & ~new_n7081_));
  assign new_n7087_ = ~\all_features[3055]  & (~\all_features[3054]  | (~\all_features[3053]  & (new_n7074_ | ~new_n7081_ | ~\all_features[3052] )));
  assign new_n7088_ = new_n7084_ & (~\all_features[3053]  | (~\all_features[3052]  & (~\all_features[3051]  | (~\all_features[3050]  & ~\all_features[3049] ))));
  assign new_n7089_ = new_n7095_ & (~new_n7096_ | (~new_n7090_ & ~new_n7086_ & ~new_n7087_));
  assign new_n7090_ = new_n7093_ & ((~new_n7091_ & new_n7076_ & new_n7094_) | ~new_n7082_ | ~new_n7073_);
  assign new_n7091_ = \all_features[3055]  & \all_features[3054]  & ~new_n7092_ & \all_features[3053] ;
  assign new_n7092_ = ~\all_features[3051]  & ~\all_features[3052]  & (~\all_features[3050]  | new_n7074_);
  assign new_n7093_ = ~new_n7071_ & ~new_n7080_;
  assign new_n7094_ = \all_features[3054]  & \all_features[3055]  & (\all_features[3052]  | \all_features[3053]  | new_n7079_ | ~new_n7075_);
  assign new_n7095_ = ~new_n7083_ & (\all_features[3051]  | \all_features[3052]  | \all_features[3053]  | \all_features[3054]  | \all_features[3055] );
  assign new_n7096_ = ~new_n7085_ & ~new_n7088_;
  assign new_n7097_ = ~new_n7098_ & ~new_n7101_;
  assign new_n7098_ = new_n7096_ & ~new_n7099_ & new_n7095_;
  assign new_n7099_ = new_n7100_ & (~new_n7094_ | ~new_n7082_ | ~new_n7073_ | ~new_n7076_);
  assign new_n7100_ = ~new_n7080_ & ~new_n7071_ & ~new_n7086_ & ~new_n7087_;
  assign new_n7101_ = new_n7093_ & new_n7095_ & ~new_n7088_ & ~new_n7087_ & ~new_n7085_ & ~new_n7086_;
  assign new_n7102_ = new_n7103_ & (new_n7131_ | new_n7128_);
  assign new_n7103_ = new_n7104_ & new_n7126_;
  assign new_n7104_ = new_n7123_ & ~new_n7105_ & new_n7119_;
  assign new_n7105_ = ~new_n7113_ & ~new_n7115_ & ~new_n7117_ & ~new_n7118_ & (~new_n7110_ | ~new_n7106_);
  assign new_n7106_ = \all_features[1495]  & \all_features[1494]  & ~new_n7109_ & new_n7107_;
  assign new_n7107_ = \all_features[1495]  & (\all_features[1494]  | (new_n7108_ & (\all_features[1490]  | \all_features[1491]  | \all_features[1489] )));
  assign new_n7108_ = \all_features[1492]  & \all_features[1493] ;
  assign new_n7109_ = ~\all_features[1490]  & ~\all_features[1491]  & ~\all_features[1492]  & ~\all_features[1493]  & (~\all_features[1489]  | ~\all_features[1488] );
  assign new_n7110_ = \all_features[1495]  & (\all_features[1494]  | (~new_n7111_ & \all_features[1493] ));
  assign new_n7111_ = new_n7112_ & ~\all_features[1492]  & ~\all_features[1490]  & ~\all_features[1491] ;
  assign new_n7112_ = ~\all_features[1488]  & ~\all_features[1489] ;
  assign new_n7113_ = ~\all_features[1495]  & (~\all_features[1494]  | (~\all_features[1493]  & (new_n7112_ | ~new_n7114_ | ~\all_features[1492] )));
  assign new_n7114_ = \all_features[1490]  & \all_features[1491] ;
  assign new_n7115_ = ~new_n7116_ & ~\all_features[1495] ;
  assign new_n7116_ = \all_features[1493]  & \all_features[1494]  & (\all_features[1492]  | (\all_features[1490]  & \all_features[1491]  & \all_features[1489] ));
  assign new_n7117_ = ~\all_features[1495]  & (~\all_features[1494]  | (~\all_features[1492]  & ~\all_features[1493]  & ~new_n7114_));
  assign new_n7118_ = ~\all_features[1495]  & (~new_n7114_ | ~\all_features[1488]  | ~\all_features[1489]  | ~\all_features[1494]  | ~new_n7108_);
  assign new_n7119_ = ~new_n7120_ & ~new_n7122_;
  assign new_n7120_ = ~\all_features[1493]  & new_n7121_ & ((~\all_features[1490]  & new_n7112_) | ~\all_features[1492]  | ~\all_features[1491] );
  assign new_n7121_ = ~\all_features[1494]  & ~\all_features[1495] ;
  assign new_n7122_ = ~\all_features[1495]  & ~\all_features[1494]  & ~\all_features[1493]  & ~\all_features[1491]  & ~\all_features[1492] ;
  assign new_n7123_ = ~new_n7124_ & ~new_n7125_;
  assign new_n7124_ = new_n7121_ & (~new_n7108_ | ~\all_features[1491]  | (~\all_features[1490]  & (~\all_features[1488]  | ~\all_features[1489] )));
  assign new_n7125_ = new_n7121_ & (~\all_features[1493]  | (~\all_features[1492]  & (~\all_features[1491]  | (~\all_features[1490]  & ~\all_features[1489] ))));
  assign new_n7126_ = new_n7123_ & new_n7119_ & new_n7127_ & ~new_n7115_ & ~new_n7118_;
  assign new_n7127_ = ~new_n7113_ & ~new_n7117_;
  assign new_n7128_ = new_n7119_ & (~new_n7123_ | (new_n7127_ & (new_n7129_ | new_n7115_ | new_n7118_)));
  assign new_n7129_ = new_n7110_ & (~new_n7106_ | (~new_n7130_ & \all_features[1493]  & \all_features[1494]  & \all_features[1495] ));
  assign new_n7130_ = ~\all_features[1491]  & ~\all_features[1492]  & (~\all_features[1490]  | new_n7112_);
  assign new_n7131_ = ~new_n7122_ & (new_n7120_ | (~new_n7125_ & (new_n7124_ | (~new_n7132_ & ~new_n7117_))));
  assign new_n7132_ = ~new_n7113_ & (new_n7115_ | (~new_n7118_ & (~new_n7135_ | new_n7133_)));
  assign new_n7133_ = \all_features[1495]  & ((~new_n7134_ & ~\all_features[1493]  & \all_features[1494] ) | (~new_n7107_ & (\all_features[1494]  | (~new_n7111_ & \all_features[1493] ))));
  assign new_n7134_ = (~\all_features[1490]  & ~\all_features[1491]  & ~\all_features[1492]  & (~\all_features[1489]  | ~\all_features[1488] )) | (\all_features[1492]  & (\all_features[1490]  | \all_features[1491] ));
  assign new_n7135_ = \all_features[1495]  & (\all_features[1493]  | \all_features[1494]  | \all_features[1492] );
  assign new_n7136_ = new_n7137_ & new_n7159_;
  assign new_n7137_ = new_n7154_ & ~new_n7158_ & ~new_n7138_ & ~new_n7157_;
  assign new_n7138_ = new_n7139_ & ~new_n7152_ & (~new_n7147_ | ~new_n7153_ | ~new_n7150_ | ~new_n7151_);
  assign new_n7139_ = ~new_n7144_ & ~new_n7140_ & ~new_n7142_;
  assign new_n7140_ = ~new_n7141_ & ~\all_features[4335] ;
  assign new_n7141_ = \all_features[4333]  & \all_features[4334]  & (\all_features[4332]  | (\all_features[4330]  & \all_features[4331]  & \all_features[4329] ));
  assign new_n7142_ = ~\all_features[4335]  & (~\all_features[4334]  | (~\all_features[4332]  & ~\all_features[4333]  & ~new_n7143_));
  assign new_n7143_ = \all_features[4330]  & \all_features[4331] ;
  assign new_n7144_ = ~\all_features[4335]  & (~\all_features[4334]  | ~new_n7145_ | ~new_n7146_ | ~new_n7143_);
  assign new_n7145_ = \all_features[4332]  & \all_features[4333] ;
  assign new_n7146_ = \all_features[4328]  & \all_features[4329] ;
  assign new_n7147_ = \all_features[4335]  & (\all_features[4334]  | (\all_features[4333]  & (\all_features[4332]  | ~new_n7149_ | ~new_n7148_)));
  assign new_n7148_ = ~\all_features[4330]  & ~\all_features[4331] ;
  assign new_n7149_ = ~\all_features[4328]  & ~\all_features[4329] ;
  assign new_n7150_ = \all_features[4335]  & (\all_features[4334]  | (new_n7145_ & (\all_features[4330]  | \all_features[4331]  | \all_features[4329] )));
  assign new_n7151_ = \all_features[4334]  & \all_features[4335]  & (\all_features[4332]  | \all_features[4333]  | new_n7146_ | ~new_n7148_);
  assign new_n7152_ = ~\all_features[4335]  & (~\all_features[4334]  | (~\all_features[4333]  & (new_n7149_ | ~new_n7143_ | ~\all_features[4332] )));
  assign new_n7153_ = \all_features[4335]  & (\all_features[4333]  | \all_features[4334]  | \all_features[4332] );
  assign new_n7154_ = ~new_n7155_ & (\all_features[4331]  | \all_features[4332]  | \all_features[4333]  | \all_features[4334]  | \all_features[4335] );
  assign new_n7155_ = ~\all_features[4333]  & new_n7156_ & ((~\all_features[4330]  & new_n7149_) | ~\all_features[4332]  | ~\all_features[4331] );
  assign new_n7156_ = ~\all_features[4334]  & ~\all_features[4335] ;
  assign new_n7157_ = new_n7156_ & (~\all_features[4333]  | (~\all_features[4332]  & (~\all_features[4331]  | (~\all_features[4330]  & ~\all_features[4329] ))));
  assign new_n7158_ = new_n7156_ & (~\all_features[4331]  | ~new_n7145_ | (~\all_features[4330]  & ~new_n7146_));
  assign new_n7159_ = new_n7139_ & new_n7160_ & ~new_n7152_ & new_n7154_;
  assign new_n7160_ = ~new_n7157_ & ~new_n7158_;
  assign new_n7161_ = new_n6495_ & (new_n6491_ | new_n6461_);
  assign new_n7162_ = ~new_n7163_ & new_n7192_;
  assign new_n7163_ = ~new_n7164_ & ~new_n7188_;
  assign new_n7164_ = new_n7165_ & (~new_n7179_ | (new_n7175_ & new_n7186_ & new_n7187_));
  assign new_n7165_ = new_n7166_ & ~new_n7171_ & ~new_n7172_;
  assign new_n7166_ = ~new_n7167_ & ~new_n7170_;
  assign new_n7167_ = ~\all_features[3645]  & new_n7169_ & ((~\all_features[3642]  & new_n7168_) | ~\all_features[3644]  | ~\all_features[3643] );
  assign new_n7168_ = ~\all_features[3640]  & ~\all_features[3641] ;
  assign new_n7169_ = ~\all_features[3646]  & ~\all_features[3647] ;
  assign new_n7170_ = ~\all_features[3647]  & ~\all_features[3646]  & ~\all_features[3645]  & ~\all_features[3643]  & ~\all_features[3644] ;
  assign new_n7171_ = new_n7169_ & (~\all_features[3645]  | (~\all_features[3644]  & (~\all_features[3643]  | (~\all_features[3642]  & ~\all_features[3641] ))));
  assign new_n7172_ = new_n7169_ & (~\all_features[3643]  | ~new_n7174_ | (~\all_features[3642]  & ~new_n7173_));
  assign new_n7173_ = \all_features[3640]  & \all_features[3641] ;
  assign new_n7174_ = \all_features[3644]  & \all_features[3645] ;
  assign new_n7175_ = new_n7176_ & new_n7178_;
  assign new_n7176_ = \all_features[3647]  & (\all_features[3646]  | (\all_features[3645]  & (\all_features[3644]  | ~new_n7168_ | ~new_n7177_)));
  assign new_n7177_ = ~\all_features[3642]  & ~\all_features[3643] ;
  assign new_n7178_ = \all_features[3647]  & (\all_features[3645]  | \all_features[3646]  | \all_features[3644] );
  assign new_n7179_ = ~new_n7185_ & ~new_n7184_ & ~new_n7180_ & ~new_n7182_;
  assign new_n7180_ = ~\all_features[3647]  & (~\all_features[3646]  | (~\all_features[3645]  & (new_n7168_ | ~new_n7181_ | ~\all_features[3644] )));
  assign new_n7181_ = \all_features[3642]  & \all_features[3643] ;
  assign new_n7182_ = ~new_n7183_ & ~\all_features[3647] ;
  assign new_n7183_ = \all_features[3645]  & \all_features[3646]  & (\all_features[3644]  | (\all_features[3642]  & \all_features[3643]  & \all_features[3641] ));
  assign new_n7184_ = ~\all_features[3647]  & (~\all_features[3646]  | ~new_n7173_ | ~new_n7174_ | ~new_n7181_);
  assign new_n7185_ = ~\all_features[3647]  & (~\all_features[3646]  | (~\all_features[3644]  & ~\all_features[3645]  & ~new_n7181_));
  assign new_n7186_ = \all_features[3646]  & \all_features[3647]  & (\all_features[3644]  | \all_features[3645]  | new_n7173_ | ~new_n7177_);
  assign new_n7187_ = \all_features[3647]  & (\all_features[3646]  | (new_n7174_ & (\all_features[3642]  | \all_features[3643]  | \all_features[3641] )));
  assign new_n7188_ = new_n7166_ & (new_n7172_ | new_n7171_ | (~new_n7180_ & ~new_n7185_ & ~new_n7189_));
  assign new_n7189_ = ~new_n7182_ & ~new_n7184_ & (~new_n7175_ | (~new_n7190_ & new_n7186_ & new_n7187_));
  assign new_n7190_ = \all_features[3647]  & \all_features[3646]  & ~new_n7191_ & \all_features[3645] ;
  assign new_n7191_ = ~\all_features[3643]  & ~\all_features[3644]  & (~\all_features[3642]  | new_n7168_);
  assign new_n7192_ = new_n7165_ & new_n7179_;
  assign new_n7193_ = new_n7221_ & (new_n7218_ | new_n7194_);
  assign new_n7194_ = new_n7215_ & ~new_n7195_ & new_n7211_;
  assign new_n7195_ = ~new_n7196_ & ~new_n7207_ & ~new_n7209_ & ~new_n7210_ & (~new_n7202_ | ~new_n7199_);
  assign new_n7196_ = ~\all_features[1959]  & (~\all_features[1958]  | new_n7197_);
  assign new_n7197_ = ~\all_features[1957]  & (new_n7198_ | ~\all_features[1955]  | ~\all_features[1956]  | ~\all_features[1954] );
  assign new_n7198_ = ~\all_features[1952]  & ~\all_features[1953] ;
  assign new_n7199_ = \all_features[1959]  & (\all_features[1958]  | (~new_n7200_ & \all_features[1957] ));
  assign new_n7200_ = new_n7198_ & ~\all_features[1956]  & new_n7201_;
  assign new_n7201_ = ~\all_features[1954]  & ~\all_features[1955] ;
  assign new_n7202_ = new_n7203_ & new_n7206_ & (new_n7205_ | \all_features[1956]  | \all_features[1957]  | ~new_n7201_);
  assign new_n7203_ = \all_features[1959]  & (\all_features[1958]  | (new_n7204_ & (\all_features[1954]  | \all_features[1955]  | \all_features[1953] )));
  assign new_n7204_ = \all_features[1956]  & \all_features[1957] ;
  assign new_n7205_ = \all_features[1952]  & \all_features[1953] ;
  assign new_n7206_ = \all_features[1958]  & \all_features[1959] ;
  assign new_n7207_ = ~new_n7208_ & ~\all_features[1959] ;
  assign new_n7208_ = \all_features[1957]  & \all_features[1958]  & (\all_features[1956]  | (\all_features[1954]  & \all_features[1955]  & \all_features[1953] ));
  assign new_n7209_ = ~\all_features[1959]  & (~new_n7204_ | ~\all_features[1954]  | ~\all_features[1955]  | ~\all_features[1958]  | ~new_n7205_);
  assign new_n7210_ = ~\all_features[1959]  & (~\all_features[1958]  | (~\all_features[1957]  & ~\all_features[1956]  & (~\all_features[1955]  | ~\all_features[1954] )));
  assign new_n7211_ = ~new_n7212_ & ~new_n7214_;
  assign new_n7212_ = new_n7213_ & (~\all_features[1955]  | ~new_n7204_ | (~\all_features[1954]  & ~new_n7205_));
  assign new_n7213_ = ~\all_features[1958]  & ~\all_features[1959] ;
  assign new_n7214_ = new_n7213_ & (~\all_features[1957]  | (~\all_features[1956]  & (~\all_features[1955]  | (~\all_features[1954]  & ~\all_features[1953] ))));
  assign new_n7215_ = ~new_n7216_ & ~new_n7217_;
  assign new_n7216_ = ~\all_features[1957]  & new_n7213_ & ((~\all_features[1954]  & new_n7198_) | ~\all_features[1956]  | ~\all_features[1955] );
  assign new_n7217_ = ~\all_features[1959]  & ~\all_features[1958]  & ~\all_features[1957]  & ~\all_features[1955]  & ~\all_features[1956] ;
  assign new_n7218_ = new_n7215_ & (~new_n7211_ | (~new_n7196_ & ~new_n7219_ & ~new_n7210_));
  assign new_n7219_ = ~new_n7209_ & ~new_n7207_ & (~new_n7199_ | (~new_n7220_ & new_n7202_));
  assign new_n7220_ = new_n7206_ & \all_features[1957]  & ((~new_n7198_ & \all_features[1954] ) | \all_features[1956]  | \all_features[1955] );
  assign new_n7221_ = new_n7222_ & new_n7211_ & ~new_n7216_ & ~new_n7209_ & ~new_n7196_ & ~new_n7207_;
  assign new_n7222_ = ~new_n7217_ & ~new_n7210_;
  assign new_n7223_ = ~new_n7225_ & new_n7224_ & (~new_n7193_ | new_n7162_ | ~new_n7064_);
  assign new_n7224_ = (~new_n6846_ | new_n6918_) & (~new_n6972_ | (new_n7040_ ? ~new_n7136_ : ~new_n7002_));
  assign new_n7225_ = ~new_n6884_ & ~new_n6973_ & (new_n7102_ ? ~new_n7226_ : new_n7066_);
  assign new_n7226_ = ~new_n7257_ & new_n7227_;
  assign new_n7227_ = ~new_n7253_ & new_n7228_;
  assign new_n7228_ = ~new_n7229_ & ~new_n7251_;
  assign new_n7229_ = new_n7246_ & ~new_n7250_ & ~new_n7230_ & ~new_n7249_;
  assign new_n7230_ = new_n7231_ & (~new_n7244_ | ~new_n7245_ | ~new_n7241_ | ~new_n7243_);
  assign new_n7231_ = ~new_n7238_ & ~new_n7236_ & ~new_n7232_ & ~new_n7234_;
  assign new_n7232_ = ~\all_features[3295]  & (~\all_features[3294]  | (~\all_features[3292]  & ~\all_features[3293]  & ~new_n7233_));
  assign new_n7233_ = \all_features[3290]  & \all_features[3291] ;
  assign new_n7234_ = ~\all_features[3295]  & (~\all_features[3294]  | (~\all_features[3293]  & (new_n7235_ | ~new_n7233_ | ~\all_features[3292] )));
  assign new_n7235_ = ~\all_features[3288]  & ~\all_features[3289] ;
  assign new_n7236_ = ~new_n7237_ & ~\all_features[3295] ;
  assign new_n7237_ = \all_features[3293]  & \all_features[3294]  & (\all_features[3292]  | (\all_features[3290]  & \all_features[3291]  & \all_features[3289] ));
  assign new_n7238_ = ~\all_features[3295]  & (~\all_features[3294]  | ~new_n7239_ | ~new_n7240_ | ~new_n7233_);
  assign new_n7239_ = \all_features[3288]  & \all_features[3289] ;
  assign new_n7240_ = \all_features[3292]  & \all_features[3293] ;
  assign new_n7241_ = \all_features[3295]  & (\all_features[3294]  | (\all_features[3293]  & (\all_features[3292]  | ~new_n7242_ | ~new_n7235_)));
  assign new_n7242_ = ~\all_features[3290]  & ~\all_features[3291] ;
  assign new_n7243_ = \all_features[3295]  & (\all_features[3294]  | (new_n7240_ & (\all_features[3290]  | \all_features[3291]  | \all_features[3289] )));
  assign new_n7244_ = \all_features[3294]  & \all_features[3295]  & (\all_features[3292]  | \all_features[3293]  | new_n7239_ | ~new_n7242_);
  assign new_n7245_ = \all_features[3295]  & (\all_features[3293]  | \all_features[3294]  | \all_features[3292] );
  assign new_n7246_ = ~new_n7247_ & (\all_features[3291]  | \all_features[3292]  | \all_features[3293]  | \all_features[3294]  | \all_features[3295] );
  assign new_n7247_ = ~\all_features[3293]  & new_n7248_ & ((~\all_features[3290]  & new_n7235_) | ~\all_features[3292]  | ~\all_features[3291] );
  assign new_n7248_ = ~\all_features[3294]  & ~\all_features[3295] ;
  assign new_n7249_ = new_n7248_ & (~\all_features[3293]  | (~\all_features[3292]  & (~\all_features[3291]  | (~\all_features[3290]  & ~\all_features[3289] ))));
  assign new_n7250_ = new_n7248_ & (~\all_features[3291]  | ~new_n7240_ | (~\all_features[3290]  & ~new_n7239_));
  assign new_n7251_ = new_n7252_ & new_n7246_ & ~new_n7249_ & ~new_n7236_;
  assign new_n7252_ = ~new_n7238_ & ~new_n7234_ & ~new_n7250_ & ~new_n7232_;
  assign new_n7253_ = new_n7246_ & (new_n7250_ | new_n7249_ | (~new_n7254_ & ~new_n7232_ & ~new_n7234_));
  assign new_n7254_ = ~new_n7236_ & ~new_n7238_ & (~new_n7245_ | ~new_n7241_ | new_n7255_);
  assign new_n7255_ = new_n7243_ & new_n7244_ & (new_n7256_ | ~\all_features[3293]  | ~\all_features[3294]  | ~\all_features[3295] );
  assign new_n7256_ = ~\all_features[3291]  & ~\all_features[3292]  & (~\all_features[3290]  | new_n7235_);
  assign new_n7257_ = ~new_n7258_ & (\all_features[3291]  | \all_features[3292]  | \all_features[3293]  | \all_features[3294]  | \all_features[3295] );
  assign new_n7258_ = ~new_n7247_ & (new_n7249_ | (~new_n7250_ & (new_n7232_ | (~new_n7259_ & ~new_n7234_))));
  assign new_n7259_ = ~new_n7236_ & (new_n7238_ | (new_n7245_ & (~new_n7241_ | (~new_n7260_ & new_n7243_))));
  assign new_n7260_ = ~\all_features[3293]  & \all_features[3294]  & \all_features[3295]  & (\all_features[3292]  ? new_n7242_ : (new_n7239_ | ~new_n7242_));
  assign new_n7261_ = new_n7551_ & (~new_n7262_ | (~new_n7592_ & ~new_n7593_));
  assign new_n7262_ = ~new_n7514_ & new_n7263_;
  assign new_n7263_ = new_n7264_ & (new_n7268_ | new_n7442_);
  assign new_n7264_ = (new_n7374_ | ~new_n7265_ | ~new_n7267_) & (~new_n7408_ | ~new_n7338_);
  assign new_n7265_ = ~new_n7266_ & new_n7035_;
  assign new_n7266_ = ~new_n7004_ & ~new_n7025_;
  assign new_n7267_ = ~new_n7303_ & new_n7268_;
  assign new_n7268_ = new_n7269_ & (~new_n7299_ | ~new_n7295_);
  assign new_n7269_ = ~new_n7270_ & ~new_n7293_;
  assign new_n7270_ = new_n7288_ & ~new_n7292_ & ~new_n7271_ & ~new_n7291_;
  assign new_n7271_ = ~new_n7286_ & ~new_n7287_ & new_n7279_ & (~new_n7284_ | ~new_n7272_);
  assign new_n7272_ = new_n7278_ & new_n7273_ & new_n7275_;
  assign new_n7273_ = \all_features[2871]  & (\all_features[2870]  | (new_n7274_ & (\all_features[2866]  | \all_features[2867]  | \all_features[2865] )));
  assign new_n7274_ = \all_features[2868]  & \all_features[2869] ;
  assign new_n7275_ = \all_features[2870]  & \all_features[2871]  & (\all_features[2868]  | \all_features[2869]  | new_n7277_ | ~new_n7276_);
  assign new_n7276_ = ~\all_features[2866]  & ~\all_features[2867] ;
  assign new_n7277_ = \all_features[2864]  & \all_features[2865] ;
  assign new_n7278_ = \all_features[2871]  & (\all_features[2869]  | \all_features[2870]  | \all_features[2868] );
  assign new_n7279_ = ~new_n7280_ & ~new_n7282_;
  assign new_n7280_ = ~new_n7281_ & ~\all_features[2871] ;
  assign new_n7281_ = \all_features[2869]  & \all_features[2870]  & (\all_features[2868]  | (\all_features[2866]  & \all_features[2867]  & \all_features[2865] ));
  assign new_n7282_ = ~\all_features[2871]  & (~\all_features[2870]  | (~\all_features[2868]  & ~\all_features[2869]  & ~new_n7283_));
  assign new_n7283_ = \all_features[2866]  & \all_features[2867] ;
  assign new_n7284_ = \all_features[2871]  & (\all_features[2870]  | (\all_features[2869]  & (\all_features[2868]  | ~new_n7285_ | ~new_n7276_)));
  assign new_n7285_ = ~\all_features[2864]  & ~\all_features[2865] ;
  assign new_n7286_ = ~\all_features[2871]  & (~\all_features[2870]  | (~\all_features[2869]  & (new_n7285_ | ~new_n7283_ | ~\all_features[2868] )));
  assign new_n7287_ = ~\all_features[2871]  & (~\all_features[2870]  | ~new_n7274_ | ~new_n7277_ | ~new_n7283_);
  assign new_n7288_ = ~new_n7289_ & (\all_features[2867]  | \all_features[2868]  | \all_features[2869]  | \all_features[2870]  | \all_features[2871] );
  assign new_n7289_ = ~\all_features[2869]  & new_n7290_ & ((~\all_features[2866]  & new_n7285_) | ~\all_features[2868]  | ~\all_features[2867] );
  assign new_n7290_ = ~\all_features[2870]  & ~\all_features[2871] ;
  assign new_n7291_ = new_n7290_ & (~\all_features[2869]  | (~\all_features[2868]  & (~\all_features[2867]  | (~\all_features[2866]  & ~\all_features[2865] ))));
  assign new_n7292_ = new_n7290_ & (~\all_features[2867]  | ~new_n7274_ | (~\all_features[2866]  & ~new_n7277_));
  assign new_n7293_ = new_n7288_ & new_n7279_ & new_n7294_ & ~new_n7286_ & ~new_n7287_;
  assign new_n7294_ = ~new_n7291_ & ~new_n7292_;
  assign new_n7295_ = new_n7288_ & (~new_n7294_ | (~new_n7296_ & ~new_n7282_ & ~new_n7286_));
  assign new_n7296_ = ~new_n7287_ & ~new_n7280_ & (~new_n7278_ | ~new_n7284_ | new_n7297_);
  assign new_n7297_ = new_n7273_ & new_n7275_ & (new_n7298_ | ~\all_features[2869]  | ~\all_features[2870]  | ~\all_features[2871] );
  assign new_n7298_ = ~\all_features[2867]  & ~\all_features[2868]  & (~\all_features[2866]  | new_n7285_);
  assign new_n7299_ = ~new_n7300_ & (\all_features[2867]  | \all_features[2868]  | \all_features[2869]  | \all_features[2870]  | \all_features[2871] );
  assign new_n7300_ = ~new_n7289_ & (new_n7291_ | (~new_n7292_ & (new_n7282_ | (~new_n7286_ & ~new_n7301_))));
  assign new_n7301_ = ~new_n7280_ & (new_n7287_ | (new_n7278_ & (~new_n7284_ | (~new_n7302_ & new_n7273_))));
  assign new_n7302_ = ~\all_features[2869]  & \all_features[2870]  & \all_features[2871]  & (\all_features[2868]  ? new_n7276_ : (new_n7277_ | ~new_n7276_));
  assign new_n7303_ = new_n7304_ & ~new_n7330_ & ~new_n7334_;
  assign new_n7304_ = ~new_n7305_ & ~new_n7327_;
  assign new_n7305_ = new_n7322_ & ~new_n7326_ & ~new_n7306_ & ~new_n7325_;
  assign new_n7306_ = new_n7307_ & ~new_n7315_ & (~new_n7320_ | ~new_n7321_ | ~new_n7317_ | ~new_n7319_);
  assign new_n7307_ = ~new_n7312_ & ~new_n7308_ & ~new_n7310_;
  assign new_n7308_ = ~\all_features[3263]  & (~\all_features[3262]  | (~\all_features[3260]  & ~\all_features[3261]  & ~new_n7309_));
  assign new_n7309_ = \all_features[3258]  & \all_features[3259] ;
  assign new_n7310_ = ~new_n7311_ & ~\all_features[3263] ;
  assign new_n7311_ = \all_features[3261]  & \all_features[3262]  & (\all_features[3260]  | (\all_features[3258]  & \all_features[3259]  & \all_features[3257] ));
  assign new_n7312_ = ~\all_features[3263]  & (~\all_features[3262]  | ~new_n7313_ | ~new_n7314_ | ~new_n7309_);
  assign new_n7313_ = \all_features[3256]  & \all_features[3257] ;
  assign new_n7314_ = \all_features[3260]  & \all_features[3261] ;
  assign new_n7315_ = ~\all_features[3263]  & (~\all_features[3262]  | (~\all_features[3261]  & (new_n7316_ | ~new_n7309_ | ~\all_features[3260] )));
  assign new_n7316_ = ~\all_features[3256]  & ~\all_features[3257] ;
  assign new_n7317_ = \all_features[3263]  & (\all_features[3262]  | (\all_features[3261]  & (\all_features[3260]  | ~new_n7318_ | ~new_n7316_)));
  assign new_n7318_ = ~\all_features[3258]  & ~\all_features[3259] ;
  assign new_n7319_ = \all_features[3263]  & (\all_features[3262]  | (new_n7314_ & (\all_features[3258]  | \all_features[3259]  | \all_features[3257] )));
  assign new_n7320_ = \all_features[3262]  & \all_features[3263]  & (\all_features[3260]  | \all_features[3261]  | new_n7313_ | ~new_n7318_);
  assign new_n7321_ = \all_features[3263]  & (\all_features[3261]  | \all_features[3262]  | \all_features[3260] );
  assign new_n7322_ = ~new_n7323_ & (\all_features[3259]  | \all_features[3260]  | \all_features[3261]  | \all_features[3262]  | \all_features[3263] );
  assign new_n7323_ = new_n7324_ & (~\all_features[3259]  | ~new_n7314_ | (~\all_features[3258]  & ~new_n7313_));
  assign new_n7324_ = ~\all_features[3262]  & ~\all_features[3263] ;
  assign new_n7325_ = ~\all_features[3261]  & new_n7324_ & ((~\all_features[3258]  & new_n7316_) | ~\all_features[3260]  | ~\all_features[3259] );
  assign new_n7326_ = new_n7324_ & (~\all_features[3261]  | (~\all_features[3260]  & (~\all_features[3259]  | (~\all_features[3258]  & ~\all_features[3257] ))));
  assign new_n7327_ = new_n7307_ & new_n7329_ & ~new_n7315_ & new_n7328_;
  assign new_n7328_ = ~new_n7325_ & (\all_features[3259]  | \all_features[3260]  | \all_features[3261]  | \all_features[3262]  | \all_features[3263] );
  assign new_n7329_ = ~new_n7326_ & ~new_n7323_;
  assign new_n7330_ = ~new_n7331_ & (\all_features[3259]  | \all_features[3260]  | \all_features[3261]  | \all_features[3262]  | \all_features[3263] );
  assign new_n7331_ = ~new_n7325_ & (new_n7326_ | (~new_n7323_ & (new_n7308_ | (~new_n7332_ & ~new_n7315_))));
  assign new_n7332_ = ~new_n7310_ & (new_n7312_ | (new_n7321_ & (~new_n7317_ | (~new_n7333_ & new_n7319_))));
  assign new_n7333_ = ~\all_features[3261]  & \all_features[3262]  & \all_features[3263]  & (\all_features[3260]  ? new_n7318_ : (new_n7313_ | ~new_n7318_));
  assign new_n7334_ = new_n7328_ & (~new_n7329_ | (~new_n7335_ & ~new_n7308_ & ~new_n7315_));
  assign new_n7335_ = ~new_n7310_ & ~new_n7312_ & (~new_n7321_ | ~new_n7317_ | new_n7336_);
  assign new_n7336_ = new_n7319_ & new_n7320_ & (new_n7337_ | ~\all_features[3261]  | ~\all_features[3262]  | ~\all_features[3263] );
  assign new_n7337_ = ~\all_features[3259]  & ~\all_features[3260]  & (~\all_features[3258]  | new_n7316_);
  assign new_n7338_ = new_n7339_ & ~new_n7268_ & new_n6533_;
  assign new_n7339_ = new_n7340_ & new_n7366_;
  assign new_n7340_ = ~new_n7341_ & ~new_n7363_;
  assign new_n7341_ = ~new_n7362_ & ~new_n7361_ & ~new_n7360_ & ~new_n7342_ & ~new_n7358_;
  assign new_n7342_ = new_n7346_ & (~new_n7355_ | ~new_n7357_ | ~new_n7343_ | ~new_n7354_);
  assign new_n7343_ = \all_features[4319]  & (\all_features[4318]  | new_n7344_);
  assign new_n7344_ = \all_features[4317]  & (\all_features[4314]  | \all_features[4315]  | \all_features[4316]  | ~new_n7345_);
  assign new_n7345_ = ~\all_features[4312]  & ~\all_features[4313] ;
  assign new_n7346_ = ~new_n7352_ & ~new_n7351_ & ~new_n7347_ & ~new_n7349_;
  assign new_n7347_ = ~\all_features[4319]  & (~\all_features[4318]  | (~\all_features[4317]  & (new_n7345_ | ~new_n7348_ | ~\all_features[4316] )));
  assign new_n7348_ = \all_features[4314]  & \all_features[4315] ;
  assign new_n7349_ = ~new_n7350_ & ~\all_features[4319] ;
  assign new_n7350_ = \all_features[4317]  & \all_features[4318]  & (\all_features[4316]  | (\all_features[4314]  & \all_features[4315]  & \all_features[4313] ));
  assign new_n7351_ = ~\all_features[4319]  & (~\all_features[4318]  | (~\all_features[4316]  & ~\all_features[4317]  & ~new_n7348_));
  assign new_n7352_ = ~\all_features[4319]  & (~new_n7348_ | ~\all_features[4312]  | ~\all_features[4313]  | ~\all_features[4318]  | ~new_n7353_);
  assign new_n7353_ = \all_features[4316]  & \all_features[4317] ;
  assign new_n7354_ = \all_features[4319]  & (\all_features[4318]  | (new_n7353_ & (\all_features[4314]  | \all_features[4315]  | \all_features[4313] )));
  assign new_n7355_ = \all_features[4319]  & ~new_n7356_ & \all_features[4318] ;
  assign new_n7356_ = ~\all_features[4314]  & ~\all_features[4315]  & ~\all_features[4316]  & ~\all_features[4317]  & (~\all_features[4313]  | ~\all_features[4312] );
  assign new_n7357_ = \all_features[4319]  & (\all_features[4317]  | \all_features[4318]  | \all_features[4316] );
  assign new_n7358_ = new_n7359_ & (~\all_features[4317]  | (~\all_features[4316]  & (~\all_features[4315]  | (~\all_features[4314]  & ~\all_features[4313] ))));
  assign new_n7359_ = ~\all_features[4318]  & ~\all_features[4319] ;
  assign new_n7360_ = ~\all_features[4317]  & new_n7359_ & ((~\all_features[4314]  & new_n7345_) | ~\all_features[4316]  | ~\all_features[4315] );
  assign new_n7361_ = new_n7359_ & (~new_n7353_ | ~\all_features[4315]  | (~\all_features[4314]  & (~\all_features[4312]  | ~\all_features[4313] )));
  assign new_n7362_ = ~\all_features[4319]  & ~\all_features[4318]  & ~\all_features[4317]  & ~\all_features[4315]  & ~\all_features[4316] ;
  assign new_n7363_ = new_n7365_ & new_n7364_ & ~new_n7360_ & ~new_n7352_ & ~new_n7347_ & ~new_n7349_;
  assign new_n7364_ = ~new_n7351_ & ~new_n7362_;
  assign new_n7365_ = ~new_n7358_ & ~new_n7361_;
  assign new_n7366_ = ~new_n7367_ & (new_n7362_ | (~new_n7371_ & ~new_n7360_));
  assign new_n7367_ = ~new_n7360_ & ~new_n7362_ & (~new_n7365_ | (~new_n7368_ & ~new_n7347_ & ~new_n7351_));
  assign new_n7368_ = ~new_n7352_ & ~new_n7349_ & (~new_n7357_ | new_n7369_ | ~new_n7343_);
  assign new_n7369_ = ~new_n7356_ & new_n7354_ & \all_features[4318]  & \all_features[4319]  & (~\all_features[4317]  | new_n7370_);
  assign new_n7370_ = ~\all_features[4315]  & ~\all_features[4316]  & (~\all_features[4314]  | new_n7345_);
  assign new_n7371_ = ~new_n7358_ & (new_n7361_ | (~new_n7351_ & (new_n7347_ | (~new_n7349_ & ~new_n7372_))));
  assign new_n7372_ = ~new_n7352_ & (~new_n7357_ | (new_n7343_ & (~new_n7354_ | (~new_n7373_ & new_n7355_))));
  assign new_n7373_ = \all_features[4318]  & \all_features[4319]  & (\all_features[4317]  | (\all_features[4316]  & (\all_features[4315]  | \all_features[4314] )));
  assign new_n7374_ = new_n7407_ & (new_n7405_ | new_n7375_);
  assign new_n7375_ = new_n7376_ & new_n7396_;
  assign new_n7376_ = ~new_n7395_ & (new_n7394_ | (~new_n7393_ & (new_n7391_ | (~new_n7390_ & ~new_n7377_))));
  assign new_n7377_ = ~new_n7384_ & (new_n7386_ | (~new_n7388_ & (~new_n7389_ | new_n7378_)));
  assign new_n7378_ = \all_features[4103]  & ((~new_n7383_ & ~\all_features[4101]  & \all_features[4102] ) | (~new_n7381_ & (\all_features[4102]  | (~new_n7379_ & \all_features[4101] ))));
  assign new_n7379_ = new_n7380_ & ~\all_features[4100]  & ~\all_features[4098]  & ~\all_features[4099] ;
  assign new_n7380_ = ~\all_features[4096]  & ~\all_features[4097] ;
  assign new_n7381_ = \all_features[4103]  & (\all_features[4102]  | (new_n7382_ & (\all_features[4098]  | \all_features[4099]  | \all_features[4097] )));
  assign new_n7382_ = \all_features[4100]  & \all_features[4101] ;
  assign new_n7383_ = (~\all_features[4098]  & ~\all_features[4099]  & ~\all_features[4100]  & (~\all_features[4097]  | ~\all_features[4096] )) | (\all_features[4100]  & (\all_features[4098]  | \all_features[4099] ));
  assign new_n7384_ = ~\all_features[4103]  & (~\all_features[4102]  | (~\all_features[4101]  & (new_n7380_ | ~\all_features[4100]  | ~new_n7385_)));
  assign new_n7385_ = \all_features[4098]  & \all_features[4099] ;
  assign new_n7386_ = ~new_n7387_ & ~\all_features[4103] ;
  assign new_n7387_ = \all_features[4101]  & \all_features[4102]  & (\all_features[4100]  | (\all_features[4098]  & \all_features[4099]  & \all_features[4097] ));
  assign new_n7388_ = ~\all_features[4103]  & (~new_n7382_ | ~\all_features[4096]  | ~\all_features[4097]  | ~\all_features[4102]  | ~new_n7385_);
  assign new_n7389_ = \all_features[4103]  & (\all_features[4101]  | \all_features[4102]  | \all_features[4100] );
  assign new_n7390_ = ~\all_features[4103]  & (~\all_features[4102]  | (~\all_features[4100]  & ~\all_features[4101]  & ~new_n7385_));
  assign new_n7391_ = new_n7392_ & (~new_n7382_ | ~\all_features[4099]  | (~\all_features[4098]  & (~\all_features[4096]  | ~\all_features[4097] )));
  assign new_n7392_ = ~\all_features[4102]  & ~\all_features[4103] ;
  assign new_n7393_ = new_n7392_ & (~\all_features[4101]  | (~\all_features[4100]  & (~\all_features[4099]  | (~\all_features[4098]  & ~\all_features[4097] ))));
  assign new_n7394_ = ~\all_features[4101]  & new_n7392_ & ((~\all_features[4098]  & new_n7380_) | ~\all_features[4100]  | ~\all_features[4099] );
  assign new_n7395_ = ~\all_features[4103]  & ~\all_features[4102]  & ~\all_features[4101]  & ~\all_features[4099]  & ~\all_features[4100] ;
  assign new_n7396_ = new_n7404_ & (~new_n7403_ | (new_n7402_ & (new_n7397_ | new_n7386_ | new_n7388_)));
  assign new_n7397_ = new_n7398_ & (~new_n7399_ | (~new_n7401_ & \all_features[4101]  & \all_features[4102]  & \all_features[4103] ));
  assign new_n7398_ = \all_features[4103]  & (\all_features[4102]  | (~new_n7379_ & \all_features[4101] ));
  assign new_n7399_ = \all_features[4103]  & \all_features[4102]  & ~new_n7400_ & new_n7381_;
  assign new_n7400_ = ~\all_features[4098]  & ~\all_features[4099]  & ~\all_features[4100]  & ~\all_features[4101]  & (~\all_features[4097]  | ~\all_features[4096] );
  assign new_n7401_ = ~\all_features[4099]  & ~\all_features[4100]  & (~\all_features[4098]  | new_n7380_);
  assign new_n7402_ = ~new_n7390_ & ~new_n7384_;
  assign new_n7403_ = ~new_n7391_ & ~new_n7393_;
  assign new_n7404_ = ~new_n7394_ & ~new_n7395_;
  assign new_n7405_ = new_n7404_ & ~new_n7406_ & new_n7403_;
  assign new_n7406_ = ~new_n7390_ & ~new_n7384_ & ~new_n7386_ & ~new_n7388_ & (~new_n7399_ | ~new_n7398_);
  assign new_n7407_ = new_n7403_ & new_n7402_ & new_n7404_ & ~new_n7386_ & ~new_n7388_;
  assign new_n7408_ = new_n7409_ & ~new_n7434_ & ~new_n7438_;
  assign new_n7409_ = ~new_n7410_ & ~new_n7432_;
  assign new_n7410_ = new_n7427_ & ~new_n7431_ & ~new_n7411_ & ~new_n7430_;
  assign new_n7411_ = new_n7412_ & (~new_n7425_ | ~new_n7426_ | ~new_n7422_ | ~new_n7424_);
  assign new_n7412_ = ~new_n7419_ & ~new_n7417_ & ~new_n7413_ & ~new_n7415_;
  assign new_n7413_ = ~\all_features[1487]  & (~\all_features[1486]  | (~\all_features[1484]  & ~\all_features[1485]  & ~new_n7414_));
  assign new_n7414_ = \all_features[1482]  & \all_features[1483] ;
  assign new_n7415_ = ~\all_features[1487]  & (~\all_features[1486]  | (~\all_features[1485]  & (new_n7416_ | ~new_n7414_ | ~\all_features[1484] )));
  assign new_n7416_ = ~\all_features[1480]  & ~\all_features[1481] ;
  assign new_n7417_ = ~new_n7418_ & ~\all_features[1487] ;
  assign new_n7418_ = \all_features[1485]  & \all_features[1486]  & (\all_features[1484]  | (\all_features[1482]  & \all_features[1483]  & \all_features[1481] ));
  assign new_n7419_ = ~\all_features[1487]  & (~\all_features[1486]  | ~new_n7420_ | ~new_n7421_ | ~new_n7414_);
  assign new_n7420_ = \all_features[1480]  & \all_features[1481] ;
  assign new_n7421_ = \all_features[1484]  & \all_features[1485] ;
  assign new_n7422_ = \all_features[1487]  & (\all_features[1486]  | (\all_features[1485]  & (\all_features[1484]  | ~new_n7423_ | ~new_n7416_)));
  assign new_n7423_ = ~\all_features[1482]  & ~\all_features[1483] ;
  assign new_n7424_ = \all_features[1487]  & (\all_features[1486]  | (new_n7421_ & (\all_features[1482]  | \all_features[1483]  | \all_features[1481] )));
  assign new_n7425_ = \all_features[1486]  & \all_features[1487]  & (\all_features[1484]  | \all_features[1485]  | new_n7420_ | ~new_n7423_);
  assign new_n7426_ = \all_features[1487]  & (\all_features[1485]  | \all_features[1486]  | \all_features[1484] );
  assign new_n7427_ = ~new_n7428_ & (\all_features[1483]  | \all_features[1484]  | \all_features[1485]  | \all_features[1486]  | \all_features[1487] );
  assign new_n7428_ = ~\all_features[1485]  & new_n7429_ & ((~\all_features[1482]  & new_n7416_) | ~\all_features[1484]  | ~\all_features[1483] );
  assign new_n7429_ = ~\all_features[1486]  & ~\all_features[1487] ;
  assign new_n7430_ = new_n7429_ & (~\all_features[1485]  | (~\all_features[1484]  & (~\all_features[1483]  | (~\all_features[1482]  & ~\all_features[1481] ))));
  assign new_n7431_ = new_n7429_ & (~\all_features[1483]  | ~new_n7421_ | (~\all_features[1482]  & ~new_n7420_));
  assign new_n7432_ = new_n7433_ & new_n7427_ & ~new_n7430_ & ~new_n7417_;
  assign new_n7433_ = ~new_n7419_ & ~new_n7415_ & ~new_n7431_ & ~new_n7413_;
  assign new_n7434_ = ~new_n7435_ & (\all_features[1483]  | \all_features[1484]  | \all_features[1485]  | \all_features[1486]  | \all_features[1487] );
  assign new_n7435_ = ~new_n7428_ & (new_n7430_ | (~new_n7431_ & (new_n7413_ | (~new_n7436_ & ~new_n7415_))));
  assign new_n7436_ = ~new_n7417_ & (new_n7419_ | (new_n7426_ & (~new_n7422_ | (~new_n7437_ & new_n7424_))));
  assign new_n7437_ = ~\all_features[1485]  & \all_features[1486]  & \all_features[1487]  & (\all_features[1484]  ? new_n7423_ : (new_n7420_ | ~new_n7423_));
  assign new_n7438_ = new_n7427_ & (new_n7431_ | new_n7430_ | (~new_n7439_ & ~new_n7413_ & ~new_n7415_));
  assign new_n7439_ = ~new_n7417_ & ~new_n7419_ & (~new_n7426_ | ~new_n7422_ | new_n7440_);
  assign new_n7440_ = new_n7424_ & new_n7425_ & (new_n7441_ | ~\all_features[1485]  | ~\all_features[1486]  | ~\all_features[1487] );
  assign new_n7441_ = ~\all_features[1483]  & ~\all_features[1484]  & (~\all_features[1482]  | new_n7416_);
  assign new_n7442_ = (new_n7339_ | ~new_n6533_ | (new_n7509_ & ~new_n7479_)) & (new_n7443_ | ~new_n7445_ | new_n6533_);
  assign new_n7443_ = new_n7444_ & new_n6662_;
  assign new_n7444_ = new_n6640_ & new_n6670_;
  assign new_n7445_ = new_n7475_ & (new_n7477_ | new_n7446_);
  assign new_n7446_ = new_n7447_ & new_n7471_;
  assign new_n7447_ = new_n7463_ & (~new_n7466_ | (~new_n7448_ & ~new_n7469_ & ~new_n7470_));
  assign new_n7448_ = ~new_n7457_ & ~new_n7459_ & (~new_n7462_ | ~new_n7461_ | new_n7449_);
  assign new_n7449_ = new_n7450_ & new_n7452_ & (new_n7455_ | ~\all_features[2573]  | ~\all_features[2574]  | ~\all_features[2575] );
  assign new_n7450_ = \all_features[2575]  & (\all_features[2574]  | (new_n7451_ & (\all_features[2570]  | \all_features[2571]  | \all_features[2569] )));
  assign new_n7451_ = \all_features[2572]  & \all_features[2573] ;
  assign new_n7452_ = \all_features[2574]  & \all_features[2575]  & (\all_features[2572]  | \all_features[2573]  | new_n7453_ | ~new_n7454_);
  assign new_n7453_ = \all_features[2568]  & \all_features[2569] ;
  assign new_n7454_ = ~\all_features[2570]  & ~\all_features[2571] ;
  assign new_n7455_ = ~\all_features[2571]  & ~\all_features[2572]  & (~\all_features[2570]  | new_n7456_);
  assign new_n7456_ = ~\all_features[2568]  & ~\all_features[2569] ;
  assign new_n7457_ = ~new_n7458_ & ~\all_features[2575] ;
  assign new_n7458_ = \all_features[2573]  & \all_features[2574]  & (\all_features[2572]  | (\all_features[2570]  & \all_features[2571]  & \all_features[2569] ));
  assign new_n7459_ = ~\all_features[2575]  & (~\all_features[2574]  | ~new_n7460_ | ~new_n7453_ | ~new_n7451_);
  assign new_n7460_ = \all_features[2570]  & \all_features[2571] ;
  assign new_n7461_ = \all_features[2575]  & (\all_features[2574]  | (\all_features[2573]  & (\all_features[2572]  | ~new_n7454_ | ~new_n7456_)));
  assign new_n7462_ = \all_features[2575]  & (\all_features[2573]  | \all_features[2574]  | \all_features[2572] );
  assign new_n7463_ = ~new_n7464_ & (\all_features[2571]  | \all_features[2572]  | \all_features[2573]  | \all_features[2574]  | \all_features[2575] );
  assign new_n7464_ = ~\all_features[2573]  & new_n7465_ & ((~\all_features[2570]  & new_n7456_) | ~\all_features[2572]  | ~\all_features[2571] );
  assign new_n7465_ = ~\all_features[2574]  & ~\all_features[2575] ;
  assign new_n7466_ = ~new_n7467_ & ~new_n7468_;
  assign new_n7467_ = new_n7465_ & (~\all_features[2573]  | (~\all_features[2572]  & (~\all_features[2571]  | (~\all_features[2570]  & ~\all_features[2569] ))));
  assign new_n7468_ = new_n7465_ & (~\all_features[2571]  | ~new_n7451_ | (~\all_features[2570]  & ~new_n7453_));
  assign new_n7469_ = ~\all_features[2575]  & (~\all_features[2574]  | (~\all_features[2573]  & (new_n7456_ | ~new_n7460_ | ~\all_features[2572] )));
  assign new_n7470_ = ~\all_features[2575]  & (~\all_features[2574]  | (~\all_features[2572]  & ~\all_features[2573]  & ~new_n7460_));
  assign new_n7471_ = ~new_n7472_ & (\all_features[2571]  | \all_features[2572]  | \all_features[2573]  | \all_features[2574]  | \all_features[2575] );
  assign new_n7472_ = ~new_n7464_ & (new_n7467_ | (~new_n7468_ & (new_n7470_ | (~new_n7469_ & ~new_n7473_))));
  assign new_n7473_ = ~new_n7457_ & (new_n7459_ | (new_n7462_ & (~new_n7461_ | (~new_n7474_ & new_n7450_))));
  assign new_n7474_ = ~\all_features[2573]  & \all_features[2574]  & \all_features[2575]  & (\all_features[2572]  ? new_n7454_ : (new_n7453_ | ~new_n7454_));
  assign new_n7475_ = new_n7476_ & new_n7463_ & ~new_n7468_ & ~new_n7469_ & ~new_n7457_ & ~new_n7467_;
  assign new_n7476_ = ~new_n7459_ & ~new_n7470_;
  assign new_n7477_ = new_n7463_ & new_n7466_ & (new_n7478_ | new_n7457_ | new_n7469_ | ~new_n7476_);
  assign new_n7478_ = new_n7462_ & new_n7452_ & new_n7461_ & new_n7450_;
  assign new_n7479_ = new_n7480_ & new_n7501_;
  assign new_n7480_ = ~new_n7481_ & (\all_features[3691]  | \all_features[3692]  | \all_features[3693]  | \all_features[3694]  | \all_features[3695] );
  assign new_n7481_ = ~new_n7495_ & (new_n7500_ | (~new_n7497_ & (new_n7498_ | (~new_n7499_ & ~new_n7482_))));
  assign new_n7482_ = ~new_n7483_ & (new_n7492_ | (new_n7494_ & (~new_n7485_ | (~new_n7490_ & new_n7488_))));
  assign new_n7483_ = ~new_n7484_ & ~\all_features[3695] ;
  assign new_n7484_ = \all_features[3693]  & \all_features[3694]  & (\all_features[3692]  | (\all_features[3690]  & \all_features[3691]  & \all_features[3689] ));
  assign new_n7485_ = \all_features[3695]  & (\all_features[3694]  | (\all_features[3693]  & (\all_features[3692]  | ~new_n7487_ | ~new_n7486_)));
  assign new_n7486_ = ~\all_features[3688]  & ~\all_features[3689] ;
  assign new_n7487_ = ~\all_features[3690]  & ~\all_features[3691] ;
  assign new_n7488_ = \all_features[3695]  & (\all_features[3694]  | (new_n7489_ & (\all_features[3690]  | \all_features[3691]  | \all_features[3689] )));
  assign new_n7489_ = \all_features[3692]  & \all_features[3693] ;
  assign new_n7490_ = ~\all_features[3693]  & \all_features[3694]  & \all_features[3695]  & (\all_features[3692]  ? new_n7487_ : (new_n7491_ | ~new_n7487_));
  assign new_n7491_ = \all_features[3688]  & \all_features[3689] ;
  assign new_n7492_ = ~\all_features[3695]  & (~\all_features[3694]  | ~new_n7491_ | ~new_n7489_ | ~new_n7493_);
  assign new_n7493_ = \all_features[3690]  & \all_features[3691] ;
  assign new_n7494_ = \all_features[3695]  & (\all_features[3693]  | \all_features[3694]  | \all_features[3692] );
  assign new_n7495_ = ~\all_features[3693]  & new_n7496_ & ((~\all_features[3690]  & new_n7486_) | ~\all_features[3692]  | ~\all_features[3691] );
  assign new_n7496_ = ~\all_features[3694]  & ~\all_features[3695] ;
  assign new_n7497_ = new_n7496_ & (~\all_features[3691]  | ~new_n7489_ | (~\all_features[3690]  & ~new_n7491_));
  assign new_n7498_ = ~\all_features[3695]  & (~\all_features[3694]  | (~\all_features[3692]  & ~\all_features[3693]  & ~new_n7493_));
  assign new_n7499_ = ~\all_features[3695]  & (~\all_features[3694]  | (~\all_features[3693]  & (new_n7486_ | ~new_n7493_ | ~\all_features[3692] )));
  assign new_n7500_ = new_n7496_ & (~\all_features[3693]  | (~\all_features[3692]  & (~\all_features[3691]  | (~\all_features[3690]  & ~\all_features[3689] ))));
  assign new_n7501_ = new_n7507_ & (~new_n7508_ | (~new_n7502_ & ~new_n7498_ & ~new_n7499_));
  assign new_n7502_ = new_n7505_ & ((~new_n7503_ & new_n7488_ & new_n7506_) | ~new_n7494_ | ~new_n7485_);
  assign new_n7503_ = \all_features[3695]  & \all_features[3694]  & ~new_n7504_ & \all_features[3693] ;
  assign new_n7504_ = ~\all_features[3691]  & ~\all_features[3692]  & (~\all_features[3690]  | new_n7486_);
  assign new_n7505_ = ~new_n7483_ & ~new_n7492_;
  assign new_n7506_ = \all_features[3694]  & \all_features[3695]  & (\all_features[3692]  | \all_features[3693]  | new_n7491_ | ~new_n7487_);
  assign new_n7507_ = ~new_n7495_ & (\all_features[3691]  | \all_features[3692]  | \all_features[3693]  | \all_features[3694]  | \all_features[3695] );
  assign new_n7508_ = ~new_n7497_ & ~new_n7500_;
  assign new_n7509_ = ~new_n7510_ & ~new_n7513_;
  assign new_n7510_ = new_n7508_ & ~new_n7511_ & new_n7507_;
  assign new_n7511_ = new_n7512_ & (~new_n7506_ | ~new_n7494_ | ~new_n7485_ | ~new_n7488_);
  assign new_n7512_ = ~new_n7492_ & ~new_n7483_ & ~new_n7498_ & ~new_n7499_;
  assign new_n7513_ = new_n7505_ & new_n7507_ & ~new_n7500_ & ~new_n7499_ & ~new_n7497_ & ~new_n7498_;
  assign new_n7514_ = new_n7443_ & ~new_n7516_ & new_n7515_;
  assign new_n7515_ = ~new_n6533_ & ~new_n7268_;
  assign new_n7516_ = ~new_n7550_ & (~new_n7547_ | new_n7517_);
  assign new_n7517_ = ~new_n7518_ & (new_n7537_ | (~new_n7543_ & ~new_n7535_));
  assign new_n7518_ = new_n7534_ & (~new_n7538_ | (~new_n7519_ & ~new_n7541_ & ~new_n7542_));
  assign new_n7519_ = ~new_n7531_ & ~new_n7529_ & (~new_n7533_ | new_n7523_ | ~new_n7520_);
  assign new_n7520_ = \all_features[4311]  & (\all_features[4310]  | new_n7521_);
  assign new_n7521_ = \all_features[4309]  & (\all_features[4306]  | \all_features[4307]  | \all_features[4308]  | ~new_n7522_);
  assign new_n7522_ = ~\all_features[4304]  & ~\all_features[4305] ;
  assign new_n7523_ = ~new_n7526_ & new_n7524_ & \all_features[4310]  & \all_features[4311]  & (~\all_features[4309]  | new_n7528_);
  assign new_n7524_ = \all_features[4311]  & (\all_features[4310]  | (new_n7525_ & (\all_features[4306]  | \all_features[4307]  | \all_features[4305] )));
  assign new_n7525_ = \all_features[4308]  & \all_features[4309] ;
  assign new_n7526_ = ~\all_features[4309]  & ~\all_features[4308]  & ~\all_features[4307]  & ~new_n7527_ & ~\all_features[4306] ;
  assign new_n7527_ = \all_features[4304]  & \all_features[4305] ;
  assign new_n7528_ = ~\all_features[4307]  & ~\all_features[4308]  & (~\all_features[4306]  | new_n7522_);
  assign new_n7529_ = ~new_n7530_ & ~\all_features[4311] ;
  assign new_n7530_ = \all_features[4309]  & \all_features[4310]  & (\all_features[4308]  | (\all_features[4306]  & \all_features[4307]  & \all_features[4305] ));
  assign new_n7531_ = ~\all_features[4311]  & (~\all_features[4310]  | ~new_n7532_ | ~new_n7527_ | ~new_n7525_);
  assign new_n7532_ = \all_features[4306]  & \all_features[4307] ;
  assign new_n7533_ = \all_features[4311]  & (\all_features[4309]  | \all_features[4310]  | \all_features[4308] );
  assign new_n7534_ = ~new_n7535_ & ~new_n7537_;
  assign new_n7535_ = ~\all_features[4309]  & new_n7536_ & ((~\all_features[4306]  & new_n7522_) | ~\all_features[4308]  | ~\all_features[4307] );
  assign new_n7536_ = ~\all_features[4310]  & ~\all_features[4311] ;
  assign new_n7537_ = ~\all_features[4311]  & ~\all_features[4310]  & ~\all_features[4309]  & ~\all_features[4307]  & ~\all_features[4308] ;
  assign new_n7538_ = ~new_n7539_ & ~new_n7540_;
  assign new_n7539_ = new_n7536_ & (~\all_features[4309]  | (~\all_features[4308]  & (~\all_features[4307]  | (~\all_features[4306]  & ~\all_features[4305] ))));
  assign new_n7540_ = new_n7536_ & (~\all_features[4307]  | ~new_n7525_ | (~\all_features[4306]  & ~new_n7527_));
  assign new_n7541_ = ~\all_features[4311]  & (~\all_features[4310]  | (~\all_features[4309]  & (new_n7522_ | ~new_n7532_ | ~\all_features[4308] )));
  assign new_n7542_ = ~\all_features[4311]  & (~\all_features[4310]  | (~\all_features[4308]  & ~\all_features[4309]  & ~new_n7532_));
  assign new_n7543_ = ~new_n7539_ & (new_n7540_ | (~new_n7542_ & (new_n7541_ | (~new_n7529_ & ~new_n7544_))));
  assign new_n7544_ = ~new_n7531_ & (~new_n7533_ | (new_n7520_ & (~new_n7524_ | (~new_n7546_ & new_n7545_))));
  assign new_n7545_ = \all_features[4311]  & ~new_n7526_ & \all_features[4310] ;
  assign new_n7546_ = \all_features[4310]  & \all_features[4311]  & (\all_features[4309]  | (\all_features[4308]  & (\all_features[4307]  | \all_features[4306] )));
  assign new_n7547_ = new_n7534_ & new_n7538_ & (new_n7548_ | new_n7529_ | new_n7541_ | ~new_n7549_);
  assign new_n7548_ = new_n7533_ & new_n7524_ & new_n7520_ & new_n7545_;
  assign new_n7549_ = ~new_n7531_ & ~new_n7542_;
  assign new_n7550_ = new_n7549_ & new_n7534_ & ~new_n7540_ & ~new_n7541_ & ~new_n7529_ & ~new_n7539_;
  assign new_n7551_ = ~new_n7552_ & ~new_n7553_ & (~new_n7267_ | (~new_n7374_ & new_n7265_));
  assign new_n7552_ = new_n7515_ & (new_n7443_ ? new_n7516_ : ~new_n7445_);
  assign new_n7553_ = new_n7554_ & (new_n7591_ ? new_n7555_ : ~new_n7556_);
  assign new_n7554_ = new_n7268_ & new_n7303_;
  assign new_n7555_ = new_n7266_ & ~new_n7036_ & ~new_n7039_;
  assign new_n7556_ = ~new_n7587_ & new_n7557_;
  assign new_n7557_ = ~new_n7583_ & new_n7558_;
  assign new_n7558_ = ~new_n7559_ & ~new_n7581_;
  assign new_n7559_ = new_n7576_ & ~new_n7580_ & ~new_n7560_ & ~new_n7579_;
  assign new_n7560_ = new_n7561_ & (~new_n7574_ | ~new_n7575_ | ~new_n7571_ | ~new_n7573_);
  assign new_n7561_ = ~new_n7568_ & ~new_n7566_ & ~new_n7562_ & ~new_n7564_;
  assign new_n7562_ = ~\all_features[3919]  & (~\all_features[3918]  | (~\all_features[3916]  & ~\all_features[3917]  & ~new_n7563_));
  assign new_n7563_ = \all_features[3914]  & \all_features[3915] ;
  assign new_n7564_ = ~\all_features[3919]  & (~\all_features[3918]  | (~\all_features[3917]  & (new_n7565_ | ~new_n7563_ | ~\all_features[3916] )));
  assign new_n7565_ = ~\all_features[3912]  & ~\all_features[3913] ;
  assign new_n7566_ = ~new_n7567_ & ~\all_features[3919] ;
  assign new_n7567_ = \all_features[3917]  & \all_features[3918]  & (\all_features[3916]  | (\all_features[3914]  & \all_features[3915]  & \all_features[3913] ));
  assign new_n7568_ = ~\all_features[3919]  & (~\all_features[3918]  | ~new_n7569_ | ~new_n7570_ | ~new_n7563_);
  assign new_n7569_ = \all_features[3912]  & \all_features[3913] ;
  assign new_n7570_ = \all_features[3916]  & \all_features[3917] ;
  assign new_n7571_ = \all_features[3919]  & (\all_features[3918]  | (\all_features[3917]  & (\all_features[3916]  | ~new_n7572_ | ~new_n7565_)));
  assign new_n7572_ = ~\all_features[3914]  & ~\all_features[3915] ;
  assign new_n7573_ = \all_features[3919]  & (\all_features[3918]  | (new_n7570_ & (\all_features[3914]  | \all_features[3915]  | \all_features[3913] )));
  assign new_n7574_ = \all_features[3918]  & \all_features[3919]  & (\all_features[3916]  | \all_features[3917]  | new_n7569_ | ~new_n7572_);
  assign new_n7575_ = \all_features[3919]  & (\all_features[3917]  | \all_features[3918]  | \all_features[3916] );
  assign new_n7576_ = ~new_n7577_ & (\all_features[3915]  | \all_features[3916]  | \all_features[3917]  | \all_features[3918]  | \all_features[3919] );
  assign new_n7577_ = ~\all_features[3917]  & new_n7578_ & ((~\all_features[3914]  & new_n7565_) | ~\all_features[3916]  | ~\all_features[3915] );
  assign new_n7578_ = ~\all_features[3918]  & ~\all_features[3919] ;
  assign new_n7579_ = new_n7578_ & (~\all_features[3917]  | (~\all_features[3916]  & (~\all_features[3915]  | (~\all_features[3914]  & ~\all_features[3913] ))));
  assign new_n7580_ = new_n7578_ & (~\all_features[3915]  | ~new_n7570_ | (~\all_features[3914]  & ~new_n7569_));
  assign new_n7581_ = new_n7582_ & new_n7576_ & ~new_n7579_ & ~new_n7566_;
  assign new_n7582_ = ~new_n7568_ & ~new_n7564_ & ~new_n7580_ & ~new_n7562_;
  assign new_n7583_ = new_n7576_ & (new_n7580_ | new_n7579_ | (~new_n7584_ & ~new_n7562_ & ~new_n7564_));
  assign new_n7584_ = ~new_n7566_ & ~new_n7568_ & (~new_n7575_ | ~new_n7571_ | new_n7585_);
  assign new_n7585_ = new_n7573_ & new_n7574_ & (new_n7586_ | ~\all_features[3917]  | ~\all_features[3918]  | ~\all_features[3919] );
  assign new_n7586_ = ~\all_features[3915]  & ~\all_features[3916]  & (~\all_features[3914]  | new_n7565_);
  assign new_n7587_ = ~new_n7588_ & (\all_features[3915]  | \all_features[3916]  | \all_features[3917]  | \all_features[3918]  | \all_features[3919] );
  assign new_n7588_ = ~new_n7577_ & (new_n7579_ | (~new_n7580_ & (new_n7562_ | (~new_n7589_ & ~new_n7564_))));
  assign new_n7589_ = ~new_n7566_ & (new_n7568_ | (new_n7575_ & (~new_n7571_ | (~new_n7590_ & new_n7573_))));
  assign new_n7590_ = ~\all_features[3917]  & \all_features[3918]  & \all_features[3919]  & (\all_features[3916]  ? new_n7572_ : (new_n7569_ | ~new_n7572_));
  assign new_n7591_ = ~new_n7405_ & ~new_n7407_;
  assign new_n7592_ = new_n7554_ & ~new_n7591_ & new_n7556_;
  assign new_n7593_ = (new_n7555_ | ~new_n7554_ | ~new_n7591_) & (~new_n7338_ | new_n7408_);
  assign new_n7594_ = new_n7595_ ? (new_n7951_ ^ new_n8350_) : (~new_n7951_ ^ new_n8350_);
  assign new_n7595_ = ~new_n7947_ & new_n7596_;
  assign new_n7596_ = new_n7597_ & (new_n7867_ | new_n7635_ | ~new_n7600_);
  assign new_n7597_ = new_n7598_ & (new_n7600_ | new_n7698_ | ~new_n7803_ | (new_n7866_ & new_n7833_));
  assign new_n7598_ = ~new_n7669_ & (~new_n7599_ | (~new_n7799_ & new_n7771_ & new_n7737_) | (new_n7699_ & ~new_n7737_));
  assign new_n7599_ = new_n7600_ & new_n7635_;
  assign new_n7600_ = ~new_n7631_ & new_n7601_;
  assign new_n7601_ = ~new_n7627_ & new_n7602_;
  assign new_n7602_ = ~new_n7603_ & ~new_n7625_;
  assign new_n7603_ = new_n7620_ & ~new_n7624_ & ~new_n7604_ & ~new_n7623_;
  assign new_n7604_ = new_n7605_ & (~new_n7618_ | ~new_n7619_ | ~new_n7615_ | ~new_n7617_);
  assign new_n7605_ = ~new_n7612_ & ~new_n7610_ & ~new_n7606_ & ~new_n7608_;
  assign new_n7606_ = ~\all_features[5255]  & (~\all_features[5254]  | (~\all_features[5252]  & ~\all_features[5253]  & ~new_n7607_));
  assign new_n7607_ = \all_features[5250]  & \all_features[5251] ;
  assign new_n7608_ = ~\all_features[5255]  & (~\all_features[5254]  | (~\all_features[5253]  & (new_n7609_ | ~new_n7607_ | ~\all_features[5252] )));
  assign new_n7609_ = ~\all_features[5248]  & ~\all_features[5249] ;
  assign new_n7610_ = ~new_n7611_ & ~\all_features[5255] ;
  assign new_n7611_ = \all_features[5253]  & \all_features[5254]  & (\all_features[5252]  | (\all_features[5250]  & \all_features[5251]  & \all_features[5249] ));
  assign new_n7612_ = ~\all_features[5255]  & (~\all_features[5254]  | ~new_n7613_ | ~new_n7614_ | ~new_n7607_);
  assign new_n7613_ = \all_features[5248]  & \all_features[5249] ;
  assign new_n7614_ = \all_features[5252]  & \all_features[5253] ;
  assign new_n7615_ = \all_features[5255]  & (\all_features[5254]  | (\all_features[5253]  & (\all_features[5252]  | ~new_n7616_ | ~new_n7609_)));
  assign new_n7616_ = ~\all_features[5250]  & ~\all_features[5251] ;
  assign new_n7617_ = \all_features[5255]  & (\all_features[5254]  | (new_n7614_ & (\all_features[5250]  | \all_features[5251]  | \all_features[5249] )));
  assign new_n7618_ = \all_features[5254]  & \all_features[5255]  & (\all_features[5252]  | \all_features[5253]  | new_n7613_ | ~new_n7616_);
  assign new_n7619_ = \all_features[5255]  & (\all_features[5253]  | \all_features[5254]  | \all_features[5252] );
  assign new_n7620_ = ~new_n7621_ & (\all_features[5251]  | \all_features[5252]  | \all_features[5253]  | \all_features[5254]  | \all_features[5255] );
  assign new_n7621_ = ~\all_features[5253]  & new_n7622_ & ((~\all_features[5250]  & new_n7609_) | ~\all_features[5252]  | ~\all_features[5251] );
  assign new_n7622_ = ~\all_features[5254]  & ~\all_features[5255] ;
  assign new_n7623_ = new_n7622_ & (~\all_features[5253]  | (~\all_features[5252]  & (~\all_features[5251]  | (~\all_features[5250]  & ~\all_features[5249] ))));
  assign new_n7624_ = new_n7622_ & (~\all_features[5251]  | ~new_n7614_ | (~\all_features[5250]  & ~new_n7613_));
  assign new_n7625_ = new_n7626_ & new_n7620_ & ~new_n7623_ & ~new_n7610_;
  assign new_n7626_ = ~new_n7612_ & ~new_n7608_ & ~new_n7624_ & ~new_n7606_;
  assign new_n7627_ = new_n7620_ & (new_n7624_ | new_n7623_ | (~new_n7628_ & ~new_n7606_ & ~new_n7608_));
  assign new_n7628_ = ~new_n7610_ & ~new_n7612_ & (~new_n7619_ | ~new_n7615_ | new_n7629_);
  assign new_n7629_ = new_n7617_ & new_n7618_ & (new_n7630_ | ~\all_features[5253]  | ~\all_features[5254]  | ~\all_features[5255] );
  assign new_n7630_ = ~\all_features[5251]  & ~\all_features[5252]  & (~\all_features[5250]  | new_n7609_);
  assign new_n7631_ = ~new_n7632_ & (\all_features[5251]  | \all_features[5252]  | \all_features[5253]  | \all_features[5254]  | \all_features[5255] );
  assign new_n7632_ = ~new_n7621_ & (new_n7623_ | (~new_n7624_ & (new_n7606_ | (~new_n7633_ & ~new_n7608_))));
  assign new_n7633_ = ~new_n7610_ & (new_n7612_ | (new_n7619_ & (~new_n7615_ | (~new_n7634_ & new_n7617_))));
  assign new_n7634_ = ~\all_features[5253]  & \all_features[5254]  & \all_features[5255]  & (\all_features[5252]  ? new_n7616_ : (new_n7613_ | ~new_n7616_));
  assign new_n7635_ = new_n7636_ & ~new_n7661_ & ~new_n7665_;
  assign new_n7636_ = ~new_n7637_ & ~new_n7659_;
  assign new_n7637_ = new_n7654_ & ~new_n7658_ & ~new_n7638_ & ~new_n7657_;
  assign new_n7638_ = new_n7639_ & (~new_n7652_ | ~new_n7653_ | ~new_n7649_ | ~new_n7651_);
  assign new_n7639_ = ~new_n7646_ & ~new_n7644_ & ~new_n7640_ & ~new_n7642_;
  assign new_n7640_ = ~\all_features[2431]  & (~\all_features[2430]  | (~\all_features[2428]  & ~\all_features[2429]  & ~new_n7641_));
  assign new_n7641_ = \all_features[2426]  & \all_features[2427] ;
  assign new_n7642_ = ~\all_features[2431]  & (~\all_features[2430]  | (~\all_features[2429]  & (new_n7643_ | ~new_n7641_ | ~\all_features[2428] )));
  assign new_n7643_ = ~\all_features[2424]  & ~\all_features[2425] ;
  assign new_n7644_ = ~new_n7645_ & ~\all_features[2431] ;
  assign new_n7645_ = \all_features[2429]  & \all_features[2430]  & (\all_features[2428]  | (\all_features[2426]  & \all_features[2427]  & \all_features[2425] ));
  assign new_n7646_ = ~\all_features[2431]  & (~\all_features[2430]  | ~new_n7647_ | ~new_n7648_ | ~new_n7641_);
  assign new_n7647_ = \all_features[2424]  & \all_features[2425] ;
  assign new_n7648_ = \all_features[2428]  & \all_features[2429] ;
  assign new_n7649_ = \all_features[2431]  & (\all_features[2430]  | (\all_features[2429]  & (\all_features[2428]  | ~new_n7650_ | ~new_n7643_)));
  assign new_n7650_ = ~\all_features[2426]  & ~\all_features[2427] ;
  assign new_n7651_ = \all_features[2431]  & (\all_features[2430]  | (new_n7648_ & (\all_features[2426]  | \all_features[2427]  | \all_features[2425] )));
  assign new_n7652_ = \all_features[2430]  & \all_features[2431]  & (\all_features[2428]  | \all_features[2429]  | new_n7647_ | ~new_n7650_);
  assign new_n7653_ = \all_features[2431]  & (\all_features[2429]  | \all_features[2430]  | \all_features[2428] );
  assign new_n7654_ = ~new_n7655_ & (\all_features[2427]  | \all_features[2428]  | \all_features[2429]  | \all_features[2430]  | \all_features[2431] );
  assign new_n7655_ = ~\all_features[2429]  & new_n7656_ & ((~\all_features[2426]  & new_n7643_) | ~\all_features[2428]  | ~\all_features[2427] );
  assign new_n7656_ = ~\all_features[2430]  & ~\all_features[2431] ;
  assign new_n7657_ = new_n7656_ & (~\all_features[2429]  | (~\all_features[2428]  & (~\all_features[2427]  | (~\all_features[2426]  & ~\all_features[2425] ))));
  assign new_n7658_ = new_n7656_ & (~\all_features[2427]  | ~new_n7648_ | (~\all_features[2426]  & ~new_n7647_));
  assign new_n7659_ = new_n7660_ & new_n7654_ & ~new_n7657_ & ~new_n7644_;
  assign new_n7660_ = ~new_n7646_ & ~new_n7642_ & ~new_n7658_ & ~new_n7640_;
  assign new_n7661_ = ~new_n7662_ & (\all_features[2427]  | \all_features[2428]  | \all_features[2429]  | \all_features[2430]  | \all_features[2431] );
  assign new_n7662_ = ~new_n7655_ & (new_n7657_ | (~new_n7658_ & (new_n7640_ | (~new_n7663_ & ~new_n7642_))));
  assign new_n7663_ = ~new_n7644_ & (new_n7646_ | (new_n7653_ & (~new_n7649_ | (~new_n7664_ & new_n7651_))));
  assign new_n7664_ = ~\all_features[2429]  & \all_features[2430]  & \all_features[2431]  & (\all_features[2428]  ? new_n7650_ : (new_n7647_ | ~new_n7650_));
  assign new_n7665_ = new_n7654_ & (new_n7658_ | new_n7657_ | (~new_n7666_ & ~new_n7640_ & ~new_n7642_));
  assign new_n7666_ = ~new_n7644_ & ~new_n7646_ & (~new_n7653_ | ~new_n7649_ | new_n7667_);
  assign new_n7667_ = new_n7651_ & new_n7652_ & (new_n7668_ | ~\all_features[2429]  | ~\all_features[2430]  | ~\all_features[2431] );
  assign new_n7668_ = ~\all_features[2427]  & ~\all_features[2428]  & (~\all_features[2426]  | new_n7643_);
  assign new_n7669_ = new_n7698_ & ~new_n7600_ & new_n7670_;
  assign new_n7670_ = ~new_n7672_ & new_n7671_;
  assign new_n7671_ = ~new_n7192_ & new_n7163_;
  assign new_n7672_ = new_n7673_ & new_n7696_;
  assign new_n7673_ = ~new_n7695_ & ~new_n7694_ & ~new_n7693_ & ~new_n7674_ & ~new_n7691_;
  assign new_n7674_ = ~new_n7675_ & ~new_n7689_ & new_n7678_ & (~new_n7690_ | ~new_n7682_);
  assign new_n7675_ = ~\all_features[3631]  & (~\all_features[3630]  | new_n7676_);
  assign new_n7676_ = ~\all_features[3629]  & (new_n7677_ | ~\all_features[3627]  | ~\all_features[3628]  | ~\all_features[3626] );
  assign new_n7677_ = ~\all_features[3624]  & ~\all_features[3625] ;
  assign new_n7678_ = ~new_n7679_ & ~new_n7681_;
  assign new_n7679_ = ~new_n7680_ & ~\all_features[3631] ;
  assign new_n7680_ = \all_features[3629]  & \all_features[3630]  & (\all_features[3628]  | (\all_features[3626]  & \all_features[3627]  & \all_features[3625] ));
  assign new_n7681_ = ~\all_features[3631]  & (~\all_features[3630]  | (~\all_features[3629]  & ~\all_features[3628]  & (~\all_features[3627]  | ~\all_features[3626] )));
  assign new_n7682_ = new_n7688_ & new_n7683_ & new_n7685_;
  assign new_n7683_ = \all_features[3631]  & (\all_features[3630]  | (new_n7684_ & (\all_features[3626]  | \all_features[3627]  | \all_features[3625] )));
  assign new_n7684_ = \all_features[3628]  & \all_features[3629] ;
  assign new_n7685_ = \all_features[3630]  & \all_features[3631]  & (\all_features[3628]  | \all_features[3629]  | new_n7686_ | ~new_n7687_);
  assign new_n7686_ = \all_features[3624]  & \all_features[3625] ;
  assign new_n7687_ = ~\all_features[3626]  & ~\all_features[3627] ;
  assign new_n7688_ = \all_features[3631]  & (\all_features[3629]  | \all_features[3630]  | \all_features[3628] );
  assign new_n7689_ = ~\all_features[3631]  & (~new_n7684_ | ~\all_features[3626]  | ~\all_features[3627]  | ~\all_features[3630]  | ~new_n7686_);
  assign new_n7690_ = \all_features[3631]  & (\all_features[3630]  | (\all_features[3629]  & (\all_features[3628]  | ~new_n7687_ | ~new_n7677_)));
  assign new_n7691_ = new_n7692_ & (~\all_features[3627]  | ~new_n7684_ | (~\all_features[3626]  & ~new_n7686_));
  assign new_n7692_ = ~\all_features[3630]  & ~\all_features[3631] ;
  assign new_n7693_ = new_n7692_ & (~\all_features[3629]  | (~\all_features[3628]  & (~\all_features[3627]  | (~\all_features[3626]  & ~\all_features[3625] ))));
  assign new_n7694_ = ~\all_features[3629]  & new_n7692_ & ((~\all_features[3626]  & new_n7677_) | ~\all_features[3628]  | ~\all_features[3627] );
  assign new_n7695_ = ~\all_features[3631]  & ~\all_features[3630]  & ~\all_features[3629]  & ~\all_features[3627]  & ~\all_features[3628] ;
  assign new_n7696_ = new_n7697_ & new_n7678_ & ~new_n7695_ & ~new_n7689_ & ~new_n7675_ & ~new_n7694_;
  assign new_n7697_ = ~new_n7691_ & ~new_n7693_;
  assign new_n7698_ = ~new_n6734_ & (~new_n6723_ | ~new_n6732_);
  assign new_n7699_ = ~new_n7700_ & new_n7732_;
  assign new_n7700_ = ~new_n7701_ & ~new_n7722_;
  assign new_n7701_ = ~new_n7702_ & (\all_features[3219]  | \all_features[3220]  | \all_features[3221]  | \all_features[3222]  | \all_features[3223] );
  assign new_n7702_ = ~new_n7716_ & (new_n7718_ | (~new_n7719_ & (new_n7720_ | (~new_n7703_ & ~new_n7721_))));
  assign new_n7703_ = ~new_n7711_ & (new_n7713_ | (~new_n7704_ & new_n7715_));
  assign new_n7704_ = \all_features[3223]  & ((~new_n7709_ & ~\all_features[3221]  & \all_features[3222] ) | (~new_n7707_ & (\all_features[3222]  | (~new_n7705_ & \all_features[3221] ))));
  assign new_n7705_ = new_n7706_ & ~\all_features[3220]  & ~\all_features[3218]  & ~\all_features[3219] ;
  assign new_n7706_ = ~\all_features[3216]  & ~\all_features[3217] ;
  assign new_n7707_ = \all_features[3223]  & (\all_features[3222]  | (new_n7708_ & (\all_features[3218]  | \all_features[3219]  | \all_features[3217] )));
  assign new_n7708_ = \all_features[3220]  & \all_features[3221] ;
  assign new_n7709_ = (\all_features[3220]  & (\all_features[3218]  | \all_features[3219] )) | (~new_n7710_ & ~\all_features[3218]  & ~\all_features[3219]  & ~\all_features[3220] );
  assign new_n7710_ = \all_features[3216]  & \all_features[3217] ;
  assign new_n7711_ = ~new_n7712_ & ~\all_features[3223] ;
  assign new_n7712_ = \all_features[3221]  & \all_features[3222]  & (\all_features[3220]  | (\all_features[3218]  & \all_features[3219]  & \all_features[3217] ));
  assign new_n7713_ = ~\all_features[3223]  & (~\all_features[3222]  | ~new_n7710_ | ~new_n7708_ | ~new_n7714_);
  assign new_n7714_ = \all_features[3218]  & \all_features[3219] ;
  assign new_n7715_ = \all_features[3223]  & (\all_features[3221]  | \all_features[3222]  | \all_features[3220] );
  assign new_n7716_ = ~\all_features[3221]  & new_n7717_ & ((~\all_features[3218]  & new_n7706_) | ~\all_features[3220]  | ~\all_features[3219] );
  assign new_n7717_ = ~\all_features[3222]  & ~\all_features[3223] ;
  assign new_n7718_ = new_n7717_ & (~\all_features[3221]  | (~\all_features[3220]  & (~\all_features[3219]  | (~\all_features[3218]  & ~\all_features[3217] ))));
  assign new_n7719_ = new_n7717_ & (~\all_features[3219]  | ~new_n7708_ | (~\all_features[3218]  & ~new_n7710_));
  assign new_n7720_ = ~\all_features[3223]  & (~\all_features[3222]  | (~\all_features[3220]  & ~\all_features[3221]  & ~new_n7714_));
  assign new_n7721_ = ~\all_features[3223]  & (~\all_features[3222]  | (~\all_features[3221]  & (new_n7706_ | ~new_n7714_ | ~\all_features[3220] )));
  assign new_n7722_ = new_n7728_ & (~new_n7729_ | (new_n7730_ & (~new_n7731_ | new_n7723_)));
  assign new_n7723_ = new_n7724_ & (~new_n7725_ | (~new_n7727_ & \all_features[3221]  & \all_features[3222]  & \all_features[3223] ));
  assign new_n7724_ = \all_features[3223]  & (\all_features[3222]  | (~new_n7705_ & \all_features[3221] ));
  assign new_n7725_ = \all_features[3223]  & \all_features[3222]  & ~new_n7726_ & new_n7707_;
  assign new_n7726_ = ~\all_features[3221]  & ~\all_features[3220]  & ~\all_features[3219]  & ~new_n7710_ & ~\all_features[3218] ;
  assign new_n7727_ = ~\all_features[3219]  & ~\all_features[3220]  & (~\all_features[3218]  | new_n7706_);
  assign new_n7728_ = ~new_n7716_ & (\all_features[3219]  | \all_features[3220]  | \all_features[3221]  | \all_features[3222]  | \all_features[3223] );
  assign new_n7729_ = ~new_n7718_ & ~new_n7719_;
  assign new_n7730_ = ~new_n7720_ & ~new_n7721_;
  assign new_n7731_ = ~new_n7711_ & ~new_n7713_;
  assign new_n7732_ = new_n7733_ & new_n7736_;
  assign new_n7733_ = new_n7734_ & (new_n7721_ | new_n7711_ | ~new_n7735_ | (new_n7725_ & new_n7724_));
  assign new_n7734_ = new_n7728_ & new_n7729_;
  assign new_n7735_ = ~new_n7720_ & ~new_n7713_;
  assign new_n7736_ = new_n7731_ & new_n7734_ & new_n7730_;
  assign new_n7737_ = new_n7769_ & new_n7767_ & new_n7738_ & new_n7760_;
  assign new_n7738_ = ~new_n7759_ & (new_n7754_ | (~new_n7756_ & (new_n7757_ | (~new_n7739_ & ~new_n7758_))));
  assign new_n7739_ = ~new_n7746_ & (new_n7749_ | (~new_n7751_ & (~new_n7753_ | (~new_n7740_ & new_n7752_))));
  assign new_n7740_ = new_n7741_ & (\all_features[4005]  | ~new_n7745_ | (~new_n7743_ & ~\all_features[4004]  & new_n7744_) | (\all_features[4004]  & ~new_n7744_));
  assign new_n7741_ = \all_features[4007]  & (\all_features[4006]  | (new_n7742_ & (\all_features[4002]  | \all_features[4003]  | \all_features[4001] )));
  assign new_n7742_ = \all_features[4004]  & \all_features[4005] ;
  assign new_n7743_ = \all_features[4000]  & \all_features[4001] ;
  assign new_n7744_ = ~\all_features[4002]  & ~\all_features[4003] ;
  assign new_n7745_ = \all_features[4006]  & \all_features[4007] ;
  assign new_n7746_ = ~\all_features[4007]  & (~\all_features[4006]  | (~\all_features[4005]  & (new_n7747_ | ~new_n7748_ | ~\all_features[4004] )));
  assign new_n7747_ = ~\all_features[4000]  & ~\all_features[4001] ;
  assign new_n7748_ = \all_features[4002]  & \all_features[4003] ;
  assign new_n7749_ = ~new_n7750_ & ~\all_features[4007] ;
  assign new_n7750_ = \all_features[4005]  & \all_features[4006]  & (\all_features[4004]  | (\all_features[4002]  & \all_features[4003]  & \all_features[4001] ));
  assign new_n7751_ = ~\all_features[4007]  & (~\all_features[4006]  | ~new_n7743_ | ~new_n7742_ | ~new_n7748_);
  assign new_n7752_ = \all_features[4007]  & (\all_features[4006]  | (\all_features[4005]  & (\all_features[4004]  | ~new_n7744_ | ~new_n7747_)));
  assign new_n7753_ = \all_features[4007]  & (\all_features[4005]  | \all_features[4006]  | \all_features[4004] );
  assign new_n7754_ = ~\all_features[4005]  & new_n7755_ & ((~\all_features[4002]  & new_n7747_) | ~\all_features[4004]  | ~\all_features[4003] );
  assign new_n7755_ = ~\all_features[4006]  & ~\all_features[4007] ;
  assign new_n7756_ = new_n7755_ & (~\all_features[4005]  | (~\all_features[4004]  & (~\all_features[4003]  | (~\all_features[4002]  & ~\all_features[4001] ))));
  assign new_n7757_ = new_n7755_ & (~\all_features[4003]  | ~new_n7742_ | (~\all_features[4002]  & ~new_n7743_));
  assign new_n7758_ = ~\all_features[4007]  & (~\all_features[4006]  | (~\all_features[4004]  & ~\all_features[4005]  & ~new_n7748_));
  assign new_n7759_ = ~\all_features[4007]  & ~\all_features[4006]  & ~\all_features[4005]  & ~\all_features[4003]  & ~\all_features[4004] ;
  assign new_n7760_ = ~new_n7754_ & ~new_n7759_ & (~new_n7765_ | (~new_n7761_ & new_n7766_));
  assign new_n7761_ = new_n7762_ & ((~new_n7764_ & new_n7763_ & new_n7741_) | ~new_n7753_ | ~new_n7752_);
  assign new_n7762_ = ~new_n7749_ & ~new_n7751_;
  assign new_n7763_ = new_n7745_ & (new_n7743_ | \all_features[4004]  | \all_features[4005]  | ~new_n7744_);
  assign new_n7764_ = new_n7745_ & \all_features[4005]  & ((~new_n7747_ & \all_features[4002] ) | \all_features[4004]  | \all_features[4003] );
  assign new_n7765_ = ~new_n7756_ & ~new_n7757_;
  assign new_n7766_ = ~new_n7758_ & ~new_n7746_;
  assign new_n7767_ = ~new_n7759_ & ~new_n7757_ & ~new_n7756_ & ~new_n7768_ & ~new_n7754_;
  assign new_n7768_ = new_n7766_ & new_n7762_ & (~new_n7763_ | ~new_n7753_ | ~new_n7752_ | ~new_n7741_);
  assign new_n7769_ = new_n7770_ & new_n7765_ & ~new_n7749_ & ~new_n7746_ & ~new_n7754_ & ~new_n7758_;
  assign new_n7770_ = ~new_n7751_ & ~new_n7759_;
  assign new_n7771_ = ~new_n7772_ & ~new_n7798_;
  assign new_n7772_ = new_n7785_ & (~new_n7773_ | (new_n7796_ & new_n7797_ & new_n7793_ & new_n7794_));
  assign new_n7773_ = new_n7774_ & new_n7781_;
  assign new_n7774_ = ~new_n7775_ & ~new_n7777_;
  assign new_n7775_ = ~new_n7776_ & ~\all_features[3687] ;
  assign new_n7776_ = \all_features[3685]  & \all_features[3686]  & (\all_features[3684]  | (\all_features[3682]  & \all_features[3683]  & \all_features[3681] ));
  assign new_n7777_ = ~\all_features[3687]  & (~\all_features[3686]  | ~new_n7778_ | ~new_n7779_ | ~new_n7780_);
  assign new_n7778_ = \all_features[3684]  & \all_features[3685] ;
  assign new_n7779_ = \all_features[3680]  & \all_features[3681] ;
  assign new_n7780_ = \all_features[3682]  & \all_features[3683] ;
  assign new_n7781_ = ~new_n7782_ & ~new_n7783_;
  assign new_n7782_ = ~\all_features[3687]  & (~\all_features[3686]  | (~\all_features[3684]  & ~\all_features[3685]  & ~new_n7780_));
  assign new_n7783_ = ~\all_features[3687]  & (~\all_features[3686]  | (~\all_features[3685]  & (new_n7784_ | ~new_n7780_ | ~\all_features[3684] )));
  assign new_n7784_ = ~\all_features[3680]  & ~\all_features[3681] ;
  assign new_n7785_ = new_n7786_ & new_n7790_;
  assign new_n7786_ = ~new_n7787_ & ~new_n7789_;
  assign new_n7787_ = new_n7788_ & (~\all_features[3685]  | (~\all_features[3684]  & (~\all_features[3683]  | (~\all_features[3682]  & ~\all_features[3681] ))));
  assign new_n7788_ = ~\all_features[3686]  & ~\all_features[3687] ;
  assign new_n7789_ = new_n7788_ & (~\all_features[3683]  | ~new_n7778_ | (~\all_features[3682]  & ~new_n7779_));
  assign new_n7790_ = ~new_n7791_ & ~new_n7792_;
  assign new_n7791_ = ~\all_features[3685]  & new_n7788_ & ((~\all_features[3682]  & new_n7784_) | ~\all_features[3684]  | ~\all_features[3683] );
  assign new_n7792_ = ~\all_features[3687]  & ~\all_features[3686]  & ~\all_features[3685]  & ~\all_features[3683]  & ~\all_features[3684] ;
  assign new_n7793_ = \all_features[3687]  & (\all_features[3686]  | (new_n7778_ & (\all_features[3682]  | \all_features[3683]  | \all_features[3681] )));
  assign new_n7794_ = \all_features[3686]  & \all_features[3687]  & (\all_features[3684]  | \all_features[3685]  | new_n7779_ | ~new_n7795_);
  assign new_n7795_ = ~\all_features[3682]  & ~\all_features[3683] ;
  assign new_n7796_ = \all_features[3687]  & (\all_features[3686]  | (\all_features[3685]  & (\all_features[3684]  | ~new_n7795_ | ~new_n7784_)));
  assign new_n7797_ = \all_features[3687]  & (\all_features[3685]  | \all_features[3686]  | \all_features[3684] );
  assign new_n7798_ = new_n7773_ & new_n7785_;
  assign new_n7799_ = new_n7790_ & (~new_n7786_ | (~new_n7800_ & new_n7781_));
  assign new_n7800_ = new_n7774_ & ((~new_n7801_ & new_n7794_ & new_n7793_) | ~new_n7797_ | ~new_n7796_);
  assign new_n7801_ = \all_features[3687]  & \all_features[3686]  & ~new_n7802_ & \all_features[3685] ;
  assign new_n7802_ = ~\all_features[3683]  & ~\all_features[3684]  & (~\all_features[3682]  | new_n7784_);
  assign new_n7803_ = ~new_n7832_ & new_n7804_;
  assign new_n7804_ = ~new_n7805_ & ~new_n7830_;
  assign new_n7805_ = new_n7806_ & (~new_n7824_ | (new_n7820_ & (new_n7812_ | new_n7827_ | new_n7829_)));
  assign new_n7806_ = ~new_n7807_ & ~new_n7811_;
  assign new_n7807_ = new_n7808_ & ((~\all_features[3442]  & new_n7810_) | ~\all_features[3444]  | ~\all_features[3443] );
  assign new_n7808_ = ~\all_features[3445]  & new_n7809_;
  assign new_n7809_ = ~\all_features[3446]  & ~\all_features[3447] ;
  assign new_n7810_ = ~\all_features[3440]  & ~\all_features[3441] ;
  assign new_n7811_ = new_n7808_ & ~\all_features[3443]  & ~\all_features[3444] ;
  assign new_n7812_ = new_n7813_ & (~new_n7815_ | (~new_n7819_ & \all_features[3445]  & \all_features[3446]  & \all_features[3447] ));
  assign new_n7813_ = \all_features[3447]  & (\all_features[3446]  | (~new_n7814_ & \all_features[3445] ));
  assign new_n7814_ = new_n7810_ & ~\all_features[3444]  & ~\all_features[3442]  & ~\all_features[3443] ;
  assign new_n7815_ = \all_features[3447]  & \all_features[3446]  & ~new_n7818_ & new_n7816_;
  assign new_n7816_ = \all_features[3447]  & (\all_features[3446]  | (new_n7817_ & (\all_features[3442]  | \all_features[3443]  | \all_features[3441] )));
  assign new_n7817_ = \all_features[3444]  & \all_features[3445] ;
  assign new_n7818_ = ~\all_features[3442]  & ~\all_features[3443]  & ~\all_features[3444]  & ~\all_features[3445]  & (~\all_features[3441]  | ~\all_features[3440] );
  assign new_n7819_ = ~\all_features[3443]  & ~\all_features[3444]  & (~\all_features[3442]  | new_n7810_);
  assign new_n7820_ = ~new_n7821_ & ~new_n7823_;
  assign new_n7821_ = ~\all_features[3447]  & (~\all_features[3446]  | (~\all_features[3444]  & ~\all_features[3445]  & ~new_n7822_));
  assign new_n7822_ = \all_features[3442]  & \all_features[3443] ;
  assign new_n7823_ = ~\all_features[3447]  & (~\all_features[3446]  | (~\all_features[3445]  & (new_n7810_ | ~\all_features[3444]  | ~new_n7822_)));
  assign new_n7824_ = ~new_n7825_ & ~new_n7826_;
  assign new_n7825_ = new_n7809_ & (~new_n7817_ | ~\all_features[3443]  | (~\all_features[3442]  & (~\all_features[3440]  | ~\all_features[3441] )));
  assign new_n7826_ = new_n7809_ & (~\all_features[3445]  | (~\all_features[3444]  & (~\all_features[3443]  | (~\all_features[3442]  & ~\all_features[3441] ))));
  assign new_n7827_ = ~new_n7828_ & ~\all_features[3447] ;
  assign new_n7828_ = \all_features[3445]  & \all_features[3446]  & (\all_features[3444]  | (\all_features[3442]  & \all_features[3443]  & \all_features[3441] ));
  assign new_n7829_ = ~\all_features[3447]  & (~new_n7817_ | ~\all_features[3440]  | ~\all_features[3441]  | ~\all_features[3446]  | ~new_n7822_);
  assign new_n7830_ = new_n7824_ & ~new_n7831_ & new_n7806_;
  assign new_n7831_ = ~new_n7821_ & ~new_n7823_ & ~new_n7827_ & ~new_n7829_ & (~new_n7815_ | ~new_n7813_);
  assign new_n7832_ = new_n7824_ & new_n7820_ & ~new_n7829_ & ~new_n7827_ & ~new_n7807_ & ~new_n7811_;
  assign new_n7833_ = new_n7834_ & new_n7863_;
  assign new_n7834_ = new_n7835_ & new_n7859_;
  assign new_n7835_ = new_n7851_ & (~new_n7854_ | (~new_n7836_ & ~new_n7857_ & ~new_n7858_));
  assign new_n7836_ = ~new_n7845_ & ~new_n7847_ & (~new_n7850_ | ~new_n7849_ | new_n7837_);
  assign new_n7837_ = new_n7838_ & new_n7840_ & (new_n7843_ | ~\all_features[3653]  | ~\all_features[3654]  | ~\all_features[3655] );
  assign new_n7838_ = \all_features[3655]  & (\all_features[3654]  | (new_n7839_ & (\all_features[3650]  | \all_features[3651]  | \all_features[3649] )));
  assign new_n7839_ = \all_features[3652]  & \all_features[3653] ;
  assign new_n7840_ = \all_features[3654]  & \all_features[3655]  & (\all_features[3652]  | \all_features[3653]  | new_n7841_ | ~new_n7842_);
  assign new_n7841_ = \all_features[3648]  & \all_features[3649] ;
  assign new_n7842_ = ~\all_features[3650]  & ~\all_features[3651] ;
  assign new_n7843_ = ~\all_features[3651]  & ~\all_features[3652]  & (~\all_features[3650]  | new_n7844_);
  assign new_n7844_ = ~\all_features[3648]  & ~\all_features[3649] ;
  assign new_n7845_ = ~new_n7846_ & ~\all_features[3655] ;
  assign new_n7846_ = \all_features[3653]  & \all_features[3654]  & (\all_features[3652]  | (\all_features[3650]  & \all_features[3651]  & \all_features[3649] ));
  assign new_n7847_ = ~\all_features[3655]  & (~\all_features[3654]  | ~new_n7848_ | ~new_n7841_ | ~new_n7839_);
  assign new_n7848_ = \all_features[3650]  & \all_features[3651] ;
  assign new_n7849_ = \all_features[3655]  & (\all_features[3654]  | (\all_features[3653]  & (\all_features[3652]  | ~new_n7842_ | ~new_n7844_)));
  assign new_n7850_ = \all_features[3655]  & (\all_features[3653]  | \all_features[3654]  | \all_features[3652] );
  assign new_n7851_ = ~new_n7852_ & (\all_features[3651]  | \all_features[3652]  | \all_features[3653]  | \all_features[3654]  | \all_features[3655] );
  assign new_n7852_ = ~\all_features[3653]  & new_n7853_ & ((~\all_features[3650]  & new_n7844_) | ~\all_features[3652]  | ~\all_features[3651] );
  assign new_n7853_ = ~\all_features[3654]  & ~\all_features[3655] ;
  assign new_n7854_ = ~new_n7855_ & ~new_n7856_;
  assign new_n7855_ = new_n7853_ & (~\all_features[3653]  | (~\all_features[3652]  & (~\all_features[3651]  | (~\all_features[3650]  & ~\all_features[3649] ))));
  assign new_n7856_ = new_n7853_ & (~\all_features[3651]  | ~new_n7839_ | (~\all_features[3650]  & ~new_n7841_));
  assign new_n7857_ = ~\all_features[3655]  & (~\all_features[3654]  | (~\all_features[3653]  & (new_n7844_ | ~new_n7848_ | ~\all_features[3652] )));
  assign new_n7858_ = ~\all_features[3655]  & (~\all_features[3654]  | (~\all_features[3652]  & ~\all_features[3653]  & ~new_n7848_));
  assign new_n7859_ = ~new_n7860_ & (\all_features[3651]  | \all_features[3652]  | \all_features[3653]  | \all_features[3654]  | \all_features[3655] );
  assign new_n7860_ = ~new_n7852_ & (new_n7855_ | (~new_n7856_ & (new_n7858_ | (~new_n7857_ & ~new_n7861_))));
  assign new_n7861_ = ~new_n7845_ & (new_n7847_ | (new_n7850_ & (~new_n7849_ | (~new_n7862_ & new_n7838_))));
  assign new_n7862_ = ~\all_features[3653]  & \all_features[3654]  & \all_features[3655]  & (\all_features[3652]  ? new_n7842_ : (new_n7841_ | ~new_n7842_));
  assign new_n7863_ = new_n7851_ & new_n7854_ & (new_n7865_ | new_n7845_ | new_n7857_ | ~new_n7864_);
  assign new_n7864_ = ~new_n7847_ & ~new_n7858_;
  assign new_n7865_ = new_n7850_ & new_n7840_ & new_n7849_ & new_n7838_;
  assign new_n7866_ = new_n7864_ & new_n7851_ & ~new_n7856_ & ~new_n7857_ & ~new_n7845_ & ~new_n7855_;
  assign new_n7867_ = (~new_n7904_ & new_n7868_) | (~new_n7913_ & new_n7942_ & ~new_n7868_);
  assign new_n7868_ = ~new_n7902_ & (~new_n7899_ | new_n7869_);
  assign new_n7869_ = ~new_n7870_ & ~new_n7895_;
  assign new_n7870_ = new_n7890_ & (~new_n7886_ | (new_n7882_ & (new_n7871_ | new_n7892_ | new_n7894_)));
  assign new_n7871_ = new_n7875_ & new_n7881_ & (~new_n7879_ | ~new_n7877_ | new_n7872_);
  assign new_n7872_ = \all_features[1927]  & \all_features[1926]  & ~new_n7873_ & \all_features[1925] ;
  assign new_n7873_ = ~\all_features[1923]  & ~\all_features[1924]  & (~\all_features[1922]  | new_n7874_);
  assign new_n7874_ = ~\all_features[1920]  & ~\all_features[1921] ;
  assign new_n7875_ = \all_features[1927]  & (\all_features[1926]  | (\all_features[1925]  & (\all_features[1924]  | ~new_n7876_ | ~new_n7874_)));
  assign new_n7876_ = ~\all_features[1922]  & ~\all_features[1923] ;
  assign new_n7877_ = \all_features[1927]  & (\all_features[1926]  | (new_n7878_ & (\all_features[1922]  | \all_features[1923]  | \all_features[1921] )));
  assign new_n7878_ = \all_features[1924]  & \all_features[1925] ;
  assign new_n7879_ = \all_features[1926]  & \all_features[1927]  & (\all_features[1924]  | \all_features[1925]  | new_n7880_ | ~new_n7876_);
  assign new_n7880_ = \all_features[1920]  & \all_features[1921] ;
  assign new_n7881_ = \all_features[1927]  & (\all_features[1925]  | \all_features[1926]  | \all_features[1924] );
  assign new_n7882_ = ~new_n7883_ & ~new_n7885_;
  assign new_n7883_ = ~\all_features[1927]  & (~\all_features[1926]  | (~\all_features[1924]  & ~\all_features[1925]  & ~new_n7884_));
  assign new_n7884_ = \all_features[1922]  & \all_features[1923] ;
  assign new_n7885_ = ~\all_features[1927]  & (~\all_features[1926]  | (~\all_features[1925]  & (new_n7874_ | ~\all_features[1924]  | ~new_n7884_)));
  assign new_n7886_ = ~new_n7887_ & ~new_n7889_;
  assign new_n7887_ = new_n7888_ & (~\all_features[1923]  | ~new_n7878_ | (~\all_features[1922]  & ~new_n7880_));
  assign new_n7888_ = ~\all_features[1926]  & ~\all_features[1927] ;
  assign new_n7889_ = new_n7888_ & (~\all_features[1925]  | (~\all_features[1924]  & (~\all_features[1923]  | (~\all_features[1922]  & ~\all_features[1921] ))));
  assign new_n7890_ = ~new_n7891_ & (\all_features[1923]  | \all_features[1924]  | \all_features[1925]  | \all_features[1926]  | \all_features[1927] );
  assign new_n7891_ = ~\all_features[1925]  & new_n7888_ & ((~\all_features[1922]  & new_n7874_) | ~\all_features[1924]  | ~\all_features[1923] );
  assign new_n7892_ = ~new_n7893_ & ~\all_features[1927] ;
  assign new_n7893_ = \all_features[1925]  & \all_features[1926]  & (\all_features[1924]  | (\all_features[1922]  & \all_features[1923]  & \all_features[1921] ));
  assign new_n7894_ = ~\all_features[1927]  & (~\all_features[1926]  | ~new_n7884_ | ~new_n7880_ | ~new_n7878_);
  assign new_n7895_ = ~new_n7896_ & (\all_features[1923]  | \all_features[1924]  | \all_features[1925]  | \all_features[1926]  | \all_features[1927] );
  assign new_n7896_ = ~new_n7891_ & (new_n7889_ | (~new_n7887_ & (new_n7883_ | (~new_n7885_ & ~new_n7897_))));
  assign new_n7897_ = ~new_n7892_ & (new_n7894_ | (new_n7881_ & (~new_n7875_ | (~new_n7898_ & new_n7877_))));
  assign new_n7898_ = ~\all_features[1925]  & \all_features[1926]  & \all_features[1927]  & (\all_features[1924]  ? new_n7876_ : (new_n7880_ | ~new_n7876_));
  assign new_n7899_ = new_n7890_ & ~new_n7900_ & new_n7886_;
  assign new_n7900_ = new_n7901_ & (~new_n7879_ | ~new_n7881_ | ~new_n7875_ | ~new_n7877_);
  assign new_n7901_ = ~new_n7894_ & ~new_n7892_ & ~new_n7883_ & ~new_n7885_;
  assign new_n7902_ = new_n7886_ & new_n7882_ & new_n7903_ & ~new_n7892_ & ~new_n7891_;
  assign new_n7903_ = ~new_n7894_ & (\all_features[1923]  | \all_features[1924]  | \all_features[1925]  | \all_features[1926]  | \all_features[1927] );
  assign new_n7904_ = ~new_n7696_ & (~new_n7673_ | (~new_n7905_ & ~new_n7909_));
  assign new_n7905_ = ~new_n7695_ & ~new_n7694_ & (~new_n7697_ | (~new_n7906_ & ~new_n7675_ & ~new_n7681_));
  assign new_n7906_ = ~new_n7689_ & ~new_n7679_ & (~new_n7688_ | ~new_n7690_ | new_n7907_);
  assign new_n7907_ = new_n7683_ & new_n7685_ & (new_n7908_ | ~\all_features[3629]  | ~\all_features[3630]  | ~\all_features[3631] );
  assign new_n7908_ = ~\all_features[3627]  & ~\all_features[3628]  & (~\all_features[3626]  | new_n7677_);
  assign new_n7909_ = ~new_n7910_ & ~new_n7695_;
  assign new_n7910_ = ~new_n7694_ & (new_n7693_ | (~new_n7691_ & (new_n7681_ | (~new_n7675_ & ~new_n7911_))));
  assign new_n7911_ = ~new_n7679_ & (new_n7689_ | (new_n7688_ & (~new_n7690_ | (~new_n7912_ & new_n7683_))));
  assign new_n7912_ = ~\all_features[3629]  & \all_features[3630]  & \all_features[3631]  & (\all_features[3628]  ? new_n7687_ : (new_n7686_ | ~new_n7687_));
  assign new_n7913_ = new_n7914_ & new_n7935_;
  assign new_n7914_ = ~new_n7915_ & (\all_features[5059]  | \all_features[5060]  | \all_features[5061]  | \all_features[5062]  | \all_features[5063] );
  assign new_n7915_ = ~new_n7929_ & (new_n7931_ | (~new_n7932_ & (new_n7933_ | (~new_n7916_ & ~new_n7934_))));
  assign new_n7916_ = ~new_n7917_ & (new_n7926_ | (new_n7928_ & (~new_n7919_ | (~new_n7924_ & new_n7922_))));
  assign new_n7917_ = ~new_n7918_ & ~\all_features[5063] ;
  assign new_n7918_ = \all_features[5061]  & \all_features[5062]  & (\all_features[5060]  | (\all_features[5058]  & \all_features[5059]  & \all_features[5057] ));
  assign new_n7919_ = \all_features[5063]  & (\all_features[5062]  | (\all_features[5061]  & (\all_features[5060]  | ~new_n7921_ | ~new_n7920_)));
  assign new_n7920_ = ~\all_features[5056]  & ~\all_features[5057] ;
  assign new_n7921_ = ~\all_features[5058]  & ~\all_features[5059] ;
  assign new_n7922_ = \all_features[5063]  & (\all_features[5062]  | (new_n7923_ & (\all_features[5058]  | \all_features[5059]  | \all_features[5057] )));
  assign new_n7923_ = \all_features[5060]  & \all_features[5061] ;
  assign new_n7924_ = ~\all_features[5061]  & \all_features[5062]  & \all_features[5063]  & (\all_features[5060]  ? new_n7921_ : (new_n7925_ | ~new_n7921_));
  assign new_n7925_ = \all_features[5056]  & \all_features[5057] ;
  assign new_n7926_ = ~\all_features[5063]  & (~\all_features[5062]  | ~new_n7925_ | ~new_n7923_ | ~new_n7927_);
  assign new_n7927_ = \all_features[5058]  & \all_features[5059] ;
  assign new_n7928_ = \all_features[5063]  & (\all_features[5061]  | \all_features[5062]  | \all_features[5060] );
  assign new_n7929_ = ~\all_features[5061]  & new_n7930_ & ((~\all_features[5058]  & new_n7920_) | ~\all_features[5060]  | ~\all_features[5059] );
  assign new_n7930_ = ~\all_features[5062]  & ~\all_features[5063] ;
  assign new_n7931_ = new_n7930_ & (~\all_features[5061]  | (~\all_features[5060]  & (~\all_features[5059]  | (~\all_features[5058]  & ~\all_features[5057] ))));
  assign new_n7932_ = new_n7930_ & (~\all_features[5059]  | ~new_n7923_ | (~\all_features[5058]  & ~new_n7925_));
  assign new_n7933_ = ~\all_features[5063]  & (~\all_features[5062]  | (~\all_features[5060]  & ~\all_features[5061]  & ~new_n7927_));
  assign new_n7934_ = ~\all_features[5063]  & (~\all_features[5062]  | (~\all_features[5061]  & (new_n7920_ | ~new_n7927_ | ~\all_features[5060] )));
  assign new_n7935_ = new_n7941_ & (~new_n7940_ | (~new_n7936_ & ~new_n7933_ & ~new_n7934_));
  assign new_n7936_ = ~new_n7926_ & ~new_n7917_ & (~new_n7928_ | ~new_n7919_ | new_n7937_);
  assign new_n7937_ = new_n7922_ & new_n7938_ & (new_n7939_ | ~\all_features[5061]  | ~\all_features[5062]  | ~\all_features[5063] );
  assign new_n7938_ = \all_features[5062]  & \all_features[5063]  & (\all_features[5060]  | \all_features[5061]  | new_n7925_ | ~new_n7921_);
  assign new_n7939_ = ~\all_features[5059]  & ~\all_features[5060]  & (~\all_features[5058]  | new_n7920_);
  assign new_n7940_ = ~new_n7931_ & ~new_n7932_;
  assign new_n7941_ = ~new_n7929_ & (\all_features[5059]  | \all_features[5060]  | \all_features[5061]  | \all_features[5062]  | \all_features[5063] );
  assign new_n7942_ = ~new_n7943_ & ~new_n7946_;
  assign new_n7943_ = new_n7940_ & new_n7941_ & (new_n7944_ | new_n7934_ | new_n7926_ | ~new_n7945_);
  assign new_n7944_ = new_n7928_ & new_n7938_ & new_n7919_ & new_n7922_;
  assign new_n7945_ = ~new_n7933_ & ~new_n7917_;
  assign new_n7946_ = new_n7941_ & new_n7940_ & new_n7945_ & ~new_n7934_ & ~new_n7926_;
  assign new_n7947_ = new_n7948_ & (~new_n7600_ | ((new_n7737_ | ~new_n7699_ | ~new_n7635_) & (~new_n7867_ | new_n7635_)));
  assign new_n7948_ = new_n7600_ | ((new_n7670_ | ~new_n7698_) & (new_n7803_ | ~new_n7949_ | new_n7698_));
  assign new_n7949_ = ~new_n7950_ & new_n6883_;
  assign new_n7950_ = ~new_n6869_ & ~new_n6880_;
  assign new_n7951_ = ~new_n7952_ & new_n8348_;
  assign new_n7952_ = new_n7953_ & (new_n8266_ | ~new_n8265_);
  assign new_n7953_ = new_n7954_ & (~new_n8163_ | ~new_n8200_ | ~new_n8231_) & (~new_n8162_ | ~new_n8164_);
  assign new_n7954_ = (new_n8133_ | ~new_n7955_ | ~new_n7992_) & (~new_n8029_ | (~new_n8098_ & new_n8060_));
  assign new_n7955_ = ~new_n7956_ & new_n7957_;
  assign new_n7956_ = ~new_n6378_ & new_n6384_;
  assign new_n7957_ = new_n7958_ & new_n7987_;
  assign new_n7958_ = new_n7959_ & new_n7980_;
  assign new_n7959_ = ~new_n7960_ & (\all_features[2155]  | \all_features[2156]  | \all_features[2157]  | \all_features[2158]  | \all_features[2159] );
  assign new_n7960_ = ~new_n7974_ & (new_n7979_ | (~new_n7976_ & (new_n7977_ | (~new_n7978_ & ~new_n7961_))));
  assign new_n7961_ = ~new_n7962_ & (new_n7964_ | (new_n7973_ & (~new_n7968_ | (~new_n7972_ & new_n7971_))));
  assign new_n7962_ = ~new_n7963_ & ~\all_features[2159] ;
  assign new_n7963_ = \all_features[2157]  & \all_features[2158]  & (\all_features[2156]  | (\all_features[2154]  & \all_features[2155]  & \all_features[2153] ));
  assign new_n7964_ = ~\all_features[2159]  & (~\all_features[2158]  | ~new_n7965_ | ~new_n7966_ | ~new_n7967_);
  assign new_n7965_ = \all_features[2152]  & \all_features[2153] ;
  assign new_n7966_ = \all_features[2156]  & \all_features[2157] ;
  assign new_n7967_ = \all_features[2154]  & \all_features[2155] ;
  assign new_n7968_ = \all_features[2159]  & (\all_features[2158]  | (\all_features[2157]  & (\all_features[2156]  | ~new_n7970_ | ~new_n7969_)));
  assign new_n7969_ = ~\all_features[2152]  & ~\all_features[2153] ;
  assign new_n7970_ = ~\all_features[2154]  & ~\all_features[2155] ;
  assign new_n7971_ = \all_features[2159]  & (\all_features[2158]  | (new_n7966_ & (\all_features[2154]  | \all_features[2155]  | \all_features[2153] )));
  assign new_n7972_ = ~\all_features[2157]  & \all_features[2158]  & \all_features[2159]  & (\all_features[2156]  ? new_n7970_ : (new_n7965_ | ~new_n7970_));
  assign new_n7973_ = \all_features[2159]  & (\all_features[2157]  | \all_features[2158]  | \all_features[2156] );
  assign new_n7974_ = ~\all_features[2157]  & new_n7975_ & ((~\all_features[2154]  & new_n7969_) | ~\all_features[2156]  | ~\all_features[2155] );
  assign new_n7975_ = ~\all_features[2158]  & ~\all_features[2159] ;
  assign new_n7976_ = new_n7975_ & (~\all_features[2155]  | ~new_n7966_ | (~\all_features[2154]  & ~new_n7965_));
  assign new_n7977_ = ~\all_features[2159]  & (~\all_features[2158]  | (~\all_features[2156]  & ~\all_features[2157]  & ~new_n7967_));
  assign new_n7978_ = ~\all_features[2159]  & (~\all_features[2158]  | (~\all_features[2157]  & (new_n7969_ | ~new_n7967_ | ~\all_features[2156] )));
  assign new_n7979_ = new_n7975_ & (~\all_features[2157]  | (~\all_features[2156]  & (~\all_features[2155]  | (~\all_features[2154]  & ~\all_features[2153] ))));
  assign new_n7980_ = new_n7986_ & (~new_n7985_ | (~new_n7981_ & ~new_n7977_ & ~new_n7978_));
  assign new_n7981_ = ~new_n7962_ & ~new_n7964_ & (~new_n7973_ | ~new_n7968_ | new_n7982_);
  assign new_n7982_ = new_n7971_ & new_n7983_ & (new_n7984_ | ~\all_features[2157]  | ~\all_features[2158]  | ~\all_features[2159] );
  assign new_n7983_ = \all_features[2158]  & \all_features[2159]  & (\all_features[2156]  | \all_features[2157]  | new_n7965_ | ~new_n7970_);
  assign new_n7984_ = ~\all_features[2155]  & ~\all_features[2156]  & (~\all_features[2154]  | new_n7969_);
  assign new_n7985_ = ~new_n7976_ & ~new_n7979_;
  assign new_n7986_ = ~new_n7974_ & (\all_features[2155]  | \all_features[2156]  | \all_features[2157]  | \all_features[2158]  | \all_features[2159] );
  assign new_n7987_ = new_n7988_ & new_n7991_;
  assign new_n7988_ = new_n7989_ & (~new_n7990_ | (new_n7983_ & new_n7973_ & new_n7968_ & new_n7971_));
  assign new_n7989_ = new_n7985_ & new_n7986_;
  assign new_n7990_ = ~new_n7964_ & ~new_n7962_ & ~new_n7977_ & ~new_n7978_;
  assign new_n7991_ = new_n7989_ & new_n7990_;
  assign new_n7992_ = new_n7993_ & new_n8028_;
  assign new_n7993_ = new_n7994_ & new_n8026_;
  assign new_n7994_ = new_n7995_ & new_n8022_;
  assign new_n7995_ = new_n8019_ & (~new_n8015_ | (~new_n7996_ & new_n8012_));
  assign new_n7996_ = new_n7997_ & ((~new_n8004_ & new_n8008_ & new_n8007_) | ~new_n8011_ | ~new_n8010_);
  assign new_n7997_ = ~new_n7998_ & ~new_n8000_;
  assign new_n7998_ = ~new_n7999_ & ~\all_features[2399] ;
  assign new_n7999_ = \all_features[2397]  & \all_features[2398]  & (\all_features[2396]  | (\all_features[2394]  & \all_features[2395]  & \all_features[2393] ));
  assign new_n8000_ = ~\all_features[2399]  & (~\all_features[2398]  | ~new_n8001_ | ~new_n8002_ | ~new_n8003_);
  assign new_n8001_ = \all_features[2394]  & \all_features[2395] ;
  assign new_n8002_ = \all_features[2392]  & \all_features[2393] ;
  assign new_n8003_ = \all_features[2396]  & \all_features[2397] ;
  assign new_n8004_ = \all_features[2399]  & \all_features[2398]  & ~new_n8005_ & \all_features[2397] ;
  assign new_n8005_ = ~\all_features[2395]  & ~\all_features[2396]  & (~\all_features[2394]  | new_n8006_);
  assign new_n8006_ = ~\all_features[2392]  & ~\all_features[2393] ;
  assign new_n8007_ = \all_features[2399]  & (\all_features[2398]  | (new_n8003_ & (\all_features[2394]  | \all_features[2395]  | \all_features[2393] )));
  assign new_n8008_ = \all_features[2398]  & \all_features[2399]  & (\all_features[2396]  | \all_features[2397]  | new_n8002_ | ~new_n8009_);
  assign new_n8009_ = ~\all_features[2394]  & ~\all_features[2395] ;
  assign new_n8010_ = \all_features[2399]  & (\all_features[2398]  | (\all_features[2397]  & (\all_features[2396]  | ~new_n8009_ | ~new_n8006_)));
  assign new_n8011_ = \all_features[2399]  & (\all_features[2397]  | \all_features[2398]  | \all_features[2396] );
  assign new_n8012_ = ~new_n8013_ & ~new_n8014_;
  assign new_n8013_ = ~\all_features[2399]  & (~\all_features[2398]  | (~\all_features[2396]  & ~\all_features[2397]  & ~new_n8001_));
  assign new_n8014_ = ~\all_features[2399]  & (~\all_features[2398]  | (~\all_features[2397]  & (new_n8006_ | ~\all_features[2396]  | ~new_n8001_)));
  assign new_n8015_ = ~new_n8016_ & ~new_n8018_;
  assign new_n8016_ = new_n8017_ & (~\all_features[2397]  | (~\all_features[2396]  & (~\all_features[2395]  | (~\all_features[2394]  & ~\all_features[2393] ))));
  assign new_n8017_ = ~\all_features[2398]  & ~\all_features[2399] ;
  assign new_n8018_ = new_n8017_ & (~\all_features[2395]  | ~new_n8003_ | (~\all_features[2394]  & ~new_n8002_));
  assign new_n8019_ = ~new_n8020_ & ~new_n8021_;
  assign new_n8020_ = ~\all_features[2397]  & new_n8017_ & ((~\all_features[2394]  & new_n8006_) | ~\all_features[2396]  | ~\all_features[2395] );
  assign new_n8021_ = ~\all_features[2399]  & ~\all_features[2398]  & ~\all_features[2397]  & ~\all_features[2395]  & ~\all_features[2396] ;
  assign new_n8022_ = ~new_n8021_ & (new_n8020_ | new_n8023_);
  assign new_n8023_ = ~new_n8016_ & (new_n8018_ | (~new_n8013_ & (new_n8014_ | (~new_n8024_ & ~new_n7998_))));
  assign new_n8024_ = ~new_n8000_ & (~new_n8011_ | (new_n8010_ & (~new_n8007_ | (~new_n8025_ & new_n8008_))));
  assign new_n8025_ = \all_features[2398]  & \all_features[2399]  & (\all_features[2397]  | (~new_n8009_ & \all_features[2396] ));
  assign new_n8026_ = new_n8015_ & new_n8019_ & (~new_n7997_ | ~new_n8012_ | (new_n8027_ & new_n8010_));
  assign new_n8027_ = new_n8011_ & new_n8007_ & new_n8008_;
  assign new_n8028_ = new_n8019_ & new_n7997_ & new_n8012_ & new_n8015_;
  assign new_n8029_ = new_n7956_ & new_n8030_;
  assign new_n8030_ = ~new_n8031_ & new_n8055_;
  assign new_n8031_ = new_n8052_ & (~new_n8046_ | (~new_n8032_ & ~new_n8050_ & ~new_n8054_));
  assign new_n8032_ = ~new_n8043_ & ~new_n8042_ & (~new_n8045_ | ~new_n8041_ | new_n8033_);
  assign new_n8033_ = new_n8034_ & new_n8036_ & (new_n8039_ | ~\all_features[3925]  | ~\all_features[3926]  | ~\all_features[3927] );
  assign new_n8034_ = \all_features[3927]  & (\all_features[3926]  | (new_n8035_ & (\all_features[3922]  | \all_features[3923]  | \all_features[3921] )));
  assign new_n8035_ = \all_features[3924]  & \all_features[3925] ;
  assign new_n8036_ = \all_features[3926]  & \all_features[3927]  & (\all_features[3924]  | \all_features[3925]  | new_n8037_ | ~new_n8038_);
  assign new_n8037_ = \all_features[3920]  & \all_features[3921] ;
  assign new_n8038_ = ~\all_features[3922]  & ~\all_features[3923] ;
  assign new_n8039_ = ~\all_features[3923]  & ~\all_features[3924]  & (~\all_features[3922]  | new_n8040_);
  assign new_n8040_ = ~\all_features[3920]  & ~\all_features[3921] ;
  assign new_n8041_ = \all_features[3927]  & (\all_features[3926]  | (\all_features[3925]  & (\all_features[3924]  | ~new_n8040_ | ~new_n8038_)));
  assign new_n8042_ = ~\all_features[3927]  & (~new_n8035_ | ~\all_features[3922]  | ~\all_features[3923]  | ~\all_features[3926]  | ~new_n8037_);
  assign new_n8043_ = ~new_n8044_ & ~\all_features[3927] ;
  assign new_n8044_ = \all_features[3925]  & \all_features[3926]  & (\all_features[3924]  | (\all_features[3922]  & \all_features[3923]  & \all_features[3921] ));
  assign new_n8045_ = \all_features[3927]  & (\all_features[3925]  | \all_features[3926]  | \all_features[3924] );
  assign new_n8046_ = ~new_n8047_ & ~new_n8049_;
  assign new_n8047_ = new_n8048_ & (~\all_features[3923]  | ~new_n8035_ | (~\all_features[3922]  & ~new_n8037_));
  assign new_n8048_ = ~\all_features[3926]  & ~\all_features[3927] ;
  assign new_n8049_ = new_n8048_ & (~\all_features[3925]  | (~\all_features[3924]  & (~\all_features[3923]  | (~\all_features[3922]  & ~\all_features[3921] ))));
  assign new_n8050_ = ~\all_features[3927]  & (~\all_features[3926]  | new_n8051_);
  assign new_n8051_ = ~\all_features[3925]  & (new_n8040_ | ~\all_features[3923]  | ~\all_features[3924]  | ~\all_features[3922] );
  assign new_n8052_ = ~new_n8053_ & (\all_features[3923]  | \all_features[3924]  | \all_features[3925]  | \all_features[3926]  | \all_features[3927] );
  assign new_n8053_ = ~\all_features[3925]  & new_n8048_ & ((~\all_features[3922]  & new_n8040_) | ~\all_features[3924]  | ~\all_features[3923] );
  assign new_n8054_ = ~\all_features[3927]  & (~\all_features[3926]  | (~\all_features[3925]  & ~\all_features[3924]  & (~\all_features[3923]  | ~\all_features[3922] )));
  assign new_n8055_ = ~new_n8056_ & ~new_n8059_;
  assign new_n8056_ = new_n8046_ & new_n8052_ & (new_n8050_ | new_n8057_ | new_n8042_ | ~new_n8058_);
  assign new_n8057_ = new_n8045_ & new_n8041_ & new_n8034_ & new_n8036_;
  assign new_n8058_ = ~new_n8043_ & ~new_n8054_;
  assign new_n8059_ = new_n8046_ & new_n8058_ & new_n8052_ & ~new_n8050_ & ~new_n8042_;
  assign new_n8060_ = ~new_n8061_ & new_n8093_;
  assign new_n8061_ = new_n8062_ & new_n8083_;
  assign new_n8062_ = ~new_n8063_ & (\all_features[1915]  | \all_features[1916]  | \all_features[1917]  | \all_features[1918]  | \all_features[1919] );
  assign new_n8063_ = ~new_n8077_ & (new_n8079_ | (~new_n8080_ & (new_n8081_ | (~new_n8064_ & ~new_n8082_))));
  assign new_n8064_ = ~new_n8072_ & (new_n8074_ | (~new_n8065_ & new_n8076_));
  assign new_n8065_ = \all_features[1919]  & ((~new_n8070_ & ~\all_features[1917]  & \all_features[1918] ) | (~new_n8068_ & (\all_features[1918]  | (~new_n8066_ & \all_features[1917] ))));
  assign new_n8066_ = new_n8067_ & ~\all_features[1916]  & ~\all_features[1914]  & ~\all_features[1915] ;
  assign new_n8067_ = ~\all_features[1912]  & ~\all_features[1913] ;
  assign new_n8068_ = \all_features[1919]  & (\all_features[1918]  | (new_n8069_ & (\all_features[1914]  | \all_features[1915]  | \all_features[1913] )));
  assign new_n8069_ = \all_features[1916]  & \all_features[1917] ;
  assign new_n8070_ = (\all_features[1916]  & (\all_features[1914]  | \all_features[1915] )) | (~new_n8071_ & ~\all_features[1914]  & ~\all_features[1915]  & ~\all_features[1916] );
  assign new_n8071_ = \all_features[1912]  & \all_features[1913] ;
  assign new_n8072_ = ~new_n8073_ & ~\all_features[1919] ;
  assign new_n8073_ = \all_features[1917]  & \all_features[1918]  & (\all_features[1916]  | (\all_features[1914]  & \all_features[1915]  & \all_features[1913] ));
  assign new_n8074_ = ~\all_features[1919]  & (~\all_features[1918]  | ~new_n8071_ | ~new_n8069_ | ~new_n8075_);
  assign new_n8075_ = \all_features[1914]  & \all_features[1915] ;
  assign new_n8076_ = \all_features[1919]  & (\all_features[1917]  | \all_features[1918]  | \all_features[1916] );
  assign new_n8077_ = ~\all_features[1917]  & new_n8078_ & ((~\all_features[1914]  & new_n8067_) | ~\all_features[1916]  | ~\all_features[1915] );
  assign new_n8078_ = ~\all_features[1918]  & ~\all_features[1919] ;
  assign new_n8079_ = new_n8078_ & (~\all_features[1917]  | (~\all_features[1916]  & (~\all_features[1915]  | (~\all_features[1914]  & ~\all_features[1913] ))));
  assign new_n8080_ = new_n8078_ & (~\all_features[1915]  | ~new_n8069_ | (~\all_features[1914]  & ~new_n8071_));
  assign new_n8081_ = ~\all_features[1919]  & (~\all_features[1918]  | (~\all_features[1916]  & ~\all_features[1917]  & ~new_n8075_));
  assign new_n8082_ = ~\all_features[1919]  & (~\all_features[1918]  | (~\all_features[1917]  & (new_n8067_ | ~new_n8075_ | ~\all_features[1916] )));
  assign new_n8083_ = new_n8089_ & (~new_n8090_ | (new_n8091_ & (~new_n8092_ | new_n8084_)));
  assign new_n8084_ = new_n8085_ & (~new_n8086_ | (~new_n8088_ & \all_features[1917]  & \all_features[1918]  & \all_features[1919] ));
  assign new_n8085_ = \all_features[1919]  & (\all_features[1918]  | (~new_n8066_ & \all_features[1917] ));
  assign new_n8086_ = \all_features[1919]  & \all_features[1918]  & ~new_n8087_ & new_n8068_;
  assign new_n8087_ = ~\all_features[1917]  & ~\all_features[1916]  & ~\all_features[1915]  & ~new_n8071_ & ~\all_features[1914] ;
  assign new_n8088_ = ~\all_features[1915]  & ~\all_features[1916]  & (~\all_features[1914]  | new_n8067_);
  assign new_n8089_ = ~new_n8077_ & (\all_features[1915]  | \all_features[1916]  | \all_features[1917]  | \all_features[1918]  | \all_features[1919] );
  assign new_n8090_ = ~new_n8079_ & ~new_n8080_;
  assign new_n8091_ = ~new_n8081_ & ~new_n8082_;
  assign new_n8092_ = ~new_n8072_ & ~new_n8074_;
  assign new_n8093_ = ~new_n8094_ & ~new_n8097_;
  assign new_n8094_ = new_n8095_ & (new_n8082_ | new_n8072_ | ~new_n8096_ | (new_n8086_ & new_n8085_));
  assign new_n8095_ = new_n8089_ & new_n8090_;
  assign new_n8096_ = ~new_n8081_ & ~new_n8074_;
  assign new_n8097_ = new_n8092_ & new_n8095_ & new_n8091_;
  assign new_n8098_ = ~new_n8099_ & new_n8128_;
  assign new_n8099_ = new_n8100_ & new_n8121_;
  assign new_n8100_ = ~new_n8101_ & (\all_features[2587]  | \all_features[2588]  | \all_features[2589]  | \all_features[2590]  | \all_features[2591] );
  assign new_n8101_ = ~new_n8115_ & (new_n8117_ | (~new_n8118_ & (new_n8119_ | (~new_n8102_ & ~new_n8120_))));
  assign new_n8102_ = ~new_n8103_ & (new_n8112_ | (new_n8114_ & (~new_n8105_ | (~new_n8110_ & new_n8108_))));
  assign new_n8103_ = ~new_n8104_ & ~\all_features[2591] ;
  assign new_n8104_ = \all_features[2589]  & \all_features[2590]  & (\all_features[2588]  | (\all_features[2586]  & \all_features[2587]  & \all_features[2585] ));
  assign new_n8105_ = \all_features[2591]  & (\all_features[2590]  | (\all_features[2589]  & (\all_features[2588]  | ~new_n8107_ | ~new_n8106_)));
  assign new_n8106_ = ~\all_features[2584]  & ~\all_features[2585] ;
  assign new_n8107_ = ~\all_features[2586]  & ~\all_features[2587] ;
  assign new_n8108_ = \all_features[2591]  & (\all_features[2590]  | (new_n8109_ & (\all_features[2586]  | \all_features[2587]  | \all_features[2585] )));
  assign new_n8109_ = \all_features[2588]  & \all_features[2589] ;
  assign new_n8110_ = ~\all_features[2589]  & \all_features[2590]  & \all_features[2591]  & (\all_features[2588]  ? new_n8107_ : (new_n8111_ | ~new_n8107_));
  assign new_n8111_ = \all_features[2584]  & \all_features[2585] ;
  assign new_n8112_ = ~\all_features[2591]  & (~\all_features[2590]  | ~new_n8111_ | ~new_n8109_ | ~new_n8113_);
  assign new_n8113_ = \all_features[2586]  & \all_features[2587] ;
  assign new_n8114_ = \all_features[2591]  & (\all_features[2589]  | \all_features[2590]  | \all_features[2588] );
  assign new_n8115_ = ~\all_features[2589]  & new_n8116_ & ((~\all_features[2586]  & new_n8106_) | ~\all_features[2588]  | ~\all_features[2587] );
  assign new_n8116_ = ~\all_features[2590]  & ~\all_features[2591] ;
  assign new_n8117_ = new_n8116_ & (~\all_features[2589]  | (~\all_features[2588]  & (~\all_features[2587]  | (~\all_features[2586]  & ~\all_features[2585] ))));
  assign new_n8118_ = new_n8116_ & (~\all_features[2587]  | ~new_n8109_ | (~\all_features[2586]  & ~new_n8111_));
  assign new_n8119_ = ~\all_features[2591]  & (~\all_features[2590]  | (~\all_features[2588]  & ~\all_features[2589]  & ~new_n8113_));
  assign new_n8120_ = ~\all_features[2591]  & (~\all_features[2590]  | (~\all_features[2589]  & (new_n8106_ | ~new_n8113_ | ~\all_features[2588] )));
  assign new_n8121_ = new_n8127_ & (~new_n8126_ | (~new_n8122_ & ~new_n8119_ & ~new_n8120_));
  assign new_n8122_ = ~new_n8112_ & ~new_n8103_ & (~new_n8114_ | ~new_n8105_ | new_n8123_);
  assign new_n8123_ = new_n8108_ & new_n8124_ & (new_n8125_ | ~\all_features[2589]  | ~\all_features[2590]  | ~\all_features[2591] );
  assign new_n8124_ = \all_features[2590]  & \all_features[2591]  & (\all_features[2588]  | \all_features[2589]  | new_n8111_ | ~new_n8107_);
  assign new_n8125_ = ~\all_features[2587]  & ~\all_features[2588]  & (~\all_features[2586]  | new_n8106_);
  assign new_n8126_ = ~new_n8117_ & ~new_n8118_;
  assign new_n8127_ = ~new_n8115_ & (\all_features[2587]  | \all_features[2588]  | \all_features[2589]  | \all_features[2590]  | \all_features[2591] );
  assign new_n8128_ = ~new_n8129_ & ~new_n8132_;
  assign new_n8129_ = new_n8126_ & new_n8127_ & (new_n8130_ | new_n8120_ | new_n8112_ | ~new_n8131_);
  assign new_n8130_ = new_n8114_ & new_n8124_ & new_n8105_ & new_n8108_;
  assign new_n8131_ = ~new_n8119_ & ~new_n8103_;
  assign new_n8132_ = new_n8127_ & new_n8126_ & new_n8131_ & ~new_n8120_ & ~new_n8112_;
  assign new_n8133_ = new_n8161_ & new_n8134_ & new_n8159_;
  assign new_n8134_ = new_n8135_ & (~new_n8149_ | (new_n8152_ & (new_n8141_ | new_n8156_ | new_n8157_)));
  assign new_n8135_ = ~new_n8136_ & ~new_n8139_;
  assign new_n8136_ = new_n8137_ & ~\all_features[4555]  & ~\all_features[4556] ;
  assign new_n8137_ = ~\all_features[4557]  & new_n8138_;
  assign new_n8138_ = ~\all_features[4558]  & ~\all_features[4559] ;
  assign new_n8139_ = new_n8137_ & ((~\all_features[4554]  & new_n8140_) | ~\all_features[4556]  | ~\all_features[4555] );
  assign new_n8140_ = ~\all_features[4552]  & ~\all_features[4553] ;
  assign new_n8141_ = new_n8142_ & (~new_n8144_ | (~new_n8148_ & \all_features[4557]  & \all_features[4558]  & \all_features[4559] ));
  assign new_n8142_ = \all_features[4559]  & (\all_features[4558]  | (~new_n8143_ & \all_features[4557] ));
  assign new_n8143_ = new_n8140_ & ~\all_features[4556]  & ~\all_features[4554]  & ~\all_features[4555] ;
  assign new_n8144_ = \all_features[4559]  & \all_features[4558]  & ~new_n8147_ & new_n8145_;
  assign new_n8145_ = \all_features[4559]  & (\all_features[4558]  | (new_n8146_ & (\all_features[4554]  | \all_features[4555]  | \all_features[4553] )));
  assign new_n8146_ = \all_features[4556]  & \all_features[4557] ;
  assign new_n8147_ = ~\all_features[4554]  & ~\all_features[4555]  & ~\all_features[4556]  & ~\all_features[4557]  & (~\all_features[4553]  | ~\all_features[4552] );
  assign new_n8148_ = ~\all_features[4555]  & ~\all_features[4556]  & (~\all_features[4554]  | new_n8140_);
  assign new_n8149_ = ~new_n8150_ & ~new_n8151_;
  assign new_n8150_ = new_n8138_ & (~new_n8146_ | ~\all_features[4555]  | (~\all_features[4554]  & (~\all_features[4552]  | ~\all_features[4553] )));
  assign new_n8151_ = new_n8138_ & (~\all_features[4557]  | (~\all_features[4556]  & (~\all_features[4555]  | (~\all_features[4554]  & ~\all_features[4553] ))));
  assign new_n8152_ = ~new_n8153_ & ~new_n8155_;
  assign new_n8153_ = ~\all_features[4559]  & (~\all_features[4558]  | (~\all_features[4556]  & ~\all_features[4557]  & ~new_n8154_));
  assign new_n8154_ = \all_features[4554]  & \all_features[4555] ;
  assign new_n8155_ = ~\all_features[4559]  & (~\all_features[4558]  | (~\all_features[4557]  & (new_n8140_ | ~new_n8154_ | ~\all_features[4556] )));
  assign new_n8156_ = ~\all_features[4559]  & (~new_n8154_ | ~\all_features[4552]  | ~\all_features[4553]  | ~\all_features[4558]  | ~new_n8146_);
  assign new_n8157_ = ~new_n8158_ & ~\all_features[4559] ;
  assign new_n8158_ = \all_features[4557]  & \all_features[4558]  & (\all_features[4556]  | (\all_features[4554]  & \all_features[4555]  & \all_features[4553] ));
  assign new_n8159_ = new_n8149_ & ~new_n8160_ & new_n8135_;
  assign new_n8160_ = ~new_n8153_ & ~new_n8155_ & ~new_n8156_ & ~new_n8157_ & (~new_n8144_ | ~new_n8142_);
  assign new_n8161_ = new_n8152_ & new_n8149_ & ~new_n8157_ & ~new_n8156_ & ~new_n8136_ & ~new_n8139_;
  assign new_n8162_ = ~new_n7992_ & new_n7955_;
  assign new_n8163_ = ~new_n7956_ & ~new_n7957_;
  assign new_n8164_ = new_n8165_ & new_n8191_;
  assign new_n8165_ = new_n8166_ & new_n8188_;
  assign new_n8166_ = ~new_n8187_ & ~new_n8186_ & ~new_n8185_ & ~new_n8167_ & ~new_n8183_;
  assign new_n8167_ = new_n8168_ & (~new_n8181_ | ~new_n8182_ | ~new_n8178_ | ~new_n8180_);
  assign new_n8168_ = ~new_n8175_ & ~new_n8174_ & ~new_n8169_ & ~new_n8172_;
  assign new_n8169_ = ~\all_features[2127]  & (~\all_features[2126]  | (~\all_features[2125]  & (new_n8170_ | ~new_n8171_ | ~\all_features[2124] )));
  assign new_n8170_ = ~\all_features[2120]  & ~\all_features[2121] ;
  assign new_n8171_ = \all_features[2122]  & \all_features[2123] ;
  assign new_n8172_ = ~new_n8173_ & ~\all_features[2127] ;
  assign new_n8173_ = \all_features[2125]  & \all_features[2126]  & (\all_features[2124]  | (\all_features[2122]  & \all_features[2123]  & \all_features[2121] ));
  assign new_n8174_ = ~\all_features[2127]  & (~\all_features[2126]  | (~\all_features[2124]  & ~\all_features[2125]  & ~new_n8171_));
  assign new_n8175_ = ~\all_features[2127]  & (~\all_features[2126]  | ~new_n8176_ | ~new_n8177_ | ~new_n8171_);
  assign new_n8176_ = \all_features[2124]  & \all_features[2125] ;
  assign new_n8177_ = \all_features[2120]  & \all_features[2121] ;
  assign new_n8178_ = \all_features[2127]  & (\all_features[2126]  | (\all_features[2125]  & (\all_features[2124]  | ~new_n8170_ | ~new_n8179_)));
  assign new_n8179_ = ~\all_features[2122]  & ~\all_features[2123] ;
  assign new_n8180_ = \all_features[2127]  & (\all_features[2126]  | (new_n8176_ & (\all_features[2122]  | \all_features[2123]  | \all_features[2121] )));
  assign new_n8181_ = \all_features[2126]  & \all_features[2127]  & (\all_features[2124]  | \all_features[2125]  | new_n8177_ | ~new_n8179_);
  assign new_n8182_ = \all_features[2127]  & (\all_features[2125]  | \all_features[2126]  | \all_features[2124] );
  assign new_n8183_ = new_n8184_ & (~\all_features[2125]  | (~\all_features[2124]  & (~\all_features[2123]  | (~\all_features[2122]  & ~\all_features[2121] ))));
  assign new_n8184_ = ~\all_features[2126]  & ~\all_features[2127] ;
  assign new_n8185_ = ~\all_features[2125]  & new_n8184_ & ((~\all_features[2122]  & new_n8170_) | ~\all_features[2124]  | ~\all_features[2123] );
  assign new_n8186_ = new_n8184_ & (~\all_features[2123]  | ~new_n8176_ | (~\all_features[2122]  & ~new_n8177_));
  assign new_n8187_ = ~\all_features[2127]  & ~\all_features[2126]  & ~\all_features[2125]  & ~\all_features[2123]  & ~\all_features[2124] ;
  assign new_n8188_ = new_n8190_ & new_n8189_ & ~new_n8185_ & ~new_n8175_ & ~new_n8169_ & ~new_n8172_;
  assign new_n8189_ = ~new_n8174_ & ~new_n8187_;
  assign new_n8190_ = ~new_n8183_ & ~new_n8186_;
  assign new_n8191_ = new_n8192_ & new_n8196_;
  assign new_n8192_ = ~new_n8185_ & ~new_n8187_ & (~new_n8190_ | (~new_n8193_ & ~new_n8169_ & ~new_n8174_));
  assign new_n8193_ = ~new_n8175_ & ~new_n8172_ & (~new_n8182_ | ~new_n8178_ | new_n8194_);
  assign new_n8194_ = new_n8180_ & new_n8181_ & (new_n8195_ | ~\all_features[2125]  | ~\all_features[2126]  | ~\all_features[2127] );
  assign new_n8195_ = ~\all_features[2123]  & ~\all_features[2124]  & (~\all_features[2122]  | new_n8170_);
  assign new_n8196_ = ~new_n8197_ & ~new_n8187_;
  assign new_n8197_ = ~new_n8185_ & (new_n8183_ | (~new_n8186_ & (new_n8174_ | (~new_n8169_ & ~new_n8198_))));
  assign new_n8198_ = ~new_n8172_ & (new_n8175_ | (new_n8182_ & (~new_n8178_ | (~new_n8199_ & new_n8180_))));
  assign new_n8199_ = ~\all_features[2125]  & \all_features[2126]  & \all_features[2127]  & (\all_features[2124]  ? new_n8179_ : (new_n8177_ | ~new_n8179_));
  assign new_n8200_ = ~new_n8227_ & new_n8201_;
  assign new_n8201_ = ~new_n8202_ & ~new_n8225_;
  assign new_n8202_ = new_n8222_ & ~new_n8203_ & new_n8219_;
  assign new_n8203_ = ~new_n8218_ & ~new_n8217_ & ~new_n8215_ & ~new_n8204_ & ~new_n8207_;
  assign new_n8204_ = ~\all_features[3031]  & (~\all_features[3030]  | new_n8205_);
  assign new_n8205_ = ~\all_features[3029]  & (new_n8206_ | ~\all_features[3027]  | ~\all_features[3028]  | ~\all_features[3026] );
  assign new_n8206_ = ~\all_features[3024]  & ~\all_features[3025] ;
  assign new_n8207_ = new_n8214_ & new_n8213_ & new_n8208_ & new_n8210_;
  assign new_n8208_ = \all_features[3031]  & (\all_features[3030]  | (new_n8209_ & (\all_features[3026]  | \all_features[3027]  | \all_features[3025] )));
  assign new_n8209_ = \all_features[3028]  & \all_features[3029] ;
  assign new_n8210_ = \all_features[3030]  & \all_features[3031]  & (\all_features[3028]  | \all_features[3029]  | new_n8212_ | ~new_n8211_);
  assign new_n8211_ = ~\all_features[3026]  & ~\all_features[3027] ;
  assign new_n8212_ = \all_features[3024]  & \all_features[3025] ;
  assign new_n8213_ = \all_features[3031]  & (\all_features[3030]  | (\all_features[3029]  & (\all_features[3028]  | ~new_n8211_ | ~new_n8206_)));
  assign new_n8214_ = \all_features[3031]  & (\all_features[3029]  | \all_features[3030]  | \all_features[3028] );
  assign new_n8215_ = ~new_n8216_ & ~\all_features[3031] ;
  assign new_n8216_ = \all_features[3029]  & \all_features[3030]  & (\all_features[3028]  | (\all_features[3026]  & \all_features[3027]  & \all_features[3025] ));
  assign new_n8217_ = ~\all_features[3031]  & (~new_n8212_ | ~\all_features[3026]  | ~\all_features[3027]  | ~\all_features[3030]  | ~new_n8209_);
  assign new_n8218_ = ~\all_features[3031]  & (~\all_features[3030]  | (~\all_features[3029]  & ~\all_features[3028]  & (~\all_features[3027]  | ~\all_features[3026] )));
  assign new_n8219_ = ~new_n8220_ & (\all_features[3027]  | \all_features[3028]  | \all_features[3029]  | \all_features[3030]  | \all_features[3031] );
  assign new_n8220_ = ~\all_features[3029]  & new_n8221_ & ((~\all_features[3026]  & new_n8206_) | ~\all_features[3028]  | ~\all_features[3027] );
  assign new_n8221_ = ~\all_features[3030]  & ~\all_features[3031] ;
  assign new_n8222_ = ~new_n8223_ & ~new_n8224_;
  assign new_n8223_ = new_n8221_ & (~\all_features[3029]  | (~\all_features[3028]  & (~\all_features[3027]  | (~\all_features[3026]  & ~\all_features[3025] ))));
  assign new_n8224_ = new_n8221_ & (~\all_features[3027]  | ~new_n8209_ | (~new_n8212_ & ~\all_features[3026] ));
  assign new_n8225_ = new_n8219_ & new_n8226_ & ~new_n8215_ & ~new_n8223_;
  assign new_n8226_ = ~new_n8218_ & ~new_n8224_ & ~new_n8204_ & ~new_n8217_;
  assign new_n8227_ = new_n8219_ & (~new_n8222_ | (~new_n8204_ & ~new_n8228_ & ~new_n8218_));
  assign new_n8228_ = ~new_n8217_ & ~new_n8215_ & (~new_n8214_ | ~new_n8213_ | new_n8229_);
  assign new_n8229_ = new_n8208_ & new_n8210_ & (new_n8230_ | ~\all_features[3029]  | ~\all_features[3030]  | ~\all_features[3031] );
  assign new_n8230_ = ~\all_features[3027]  & ~\all_features[3028]  & (~\all_features[3026]  | new_n8206_);
  assign new_n8231_ = new_n8264_ & (new_n8232_ | (new_n8255_ & new_n8260_));
  assign new_n8232_ = ~new_n8254_ & ~new_n8253_ & ~new_n8252_ & ~new_n8233_ & ~new_n8250_;
  assign new_n8233_ = ~new_n8234_ & ~new_n8248_ & new_n8237_ & (~new_n8249_ | ~new_n8241_);
  assign new_n8234_ = ~\all_features[5023]  & (~\all_features[5022]  | new_n8235_);
  assign new_n8235_ = ~\all_features[5021]  & (new_n8236_ | ~\all_features[5019]  | ~\all_features[5020]  | ~\all_features[5018] );
  assign new_n8236_ = ~\all_features[5016]  & ~\all_features[5017] ;
  assign new_n8237_ = ~new_n8238_ & ~new_n8240_;
  assign new_n8238_ = ~new_n8239_ & ~\all_features[5023] ;
  assign new_n8239_ = \all_features[5021]  & \all_features[5022]  & (\all_features[5020]  | (\all_features[5018]  & \all_features[5019]  & \all_features[5017] ));
  assign new_n8240_ = ~\all_features[5023]  & (~\all_features[5022]  | (~\all_features[5021]  & ~\all_features[5020]  & (~\all_features[5019]  | ~\all_features[5018] )));
  assign new_n8241_ = new_n8247_ & new_n8242_ & new_n8244_;
  assign new_n8242_ = \all_features[5023]  & (\all_features[5022]  | (new_n8243_ & (\all_features[5018]  | \all_features[5019]  | \all_features[5017] )));
  assign new_n8243_ = \all_features[5020]  & \all_features[5021] ;
  assign new_n8244_ = \all_features[5022]  & \all_features[5023]  & (\all_features[5020]  | \all_features[5021]  | new_n8245_ | ~new_n8246_);
  assign new_n8245_ = \all_features[5016]  & \all_features[5017] ;
  assign new_n8246_ = ~\all_features[5018]  & ~\all_features[5019] ;
  assign new_n8247_ = \all_features[5023]  & (\all_features[5021]  | \all_features[5022]  | \all_features[5020] );
  assign new_n8248_ = ~\all_features[5023]  & (~new_n8243_ | ~\all_features[5018]  | ~\all_features[5019]  | ~\all_features[5022]  | ~new_n8245_);
  assign new_n8249_ = \all_features[5023]  & (\all_features[5022]  | (\all_features[5021]  & (\all_features[5020]  | ~new_n8246_ | ~new_n8236_)));
  assign new_n8250_ = new_n8251_ & (~\all_features[5019]  | ~new_n8243_ | (~\all_features[5018]  & ~new_n8245_));
  assign new_n8251_ = ~\all_features[5022]  & ~\all_features[5023] ;
  assign new_n8252_ = new_n8251_ & (~\all_features[5021]  | (~\all_features[5020]  & (~\all_features[5019]  | (~\all_features[5018]  & ~\all_features[5017] ))));
  assign new_n8253_ = ~\all_features[5021]  & new_n8251_ & ((~\all_features[5018]  & new_n8236_) | ~\all_features[5020]  | ~\all_features[5019] );
  assign new_n8254_ = ~\all_features[5023]  & ~\all_features[5022]  & ~\all_features[5021]  & ~\all_features[5019]  & ~\all_features[5020] ;
  assign new_n8255_ = ~new_n8254_ & ~new_n8253_ & (~new_n8259_ | (~new_n8256_ & ~new_n8234_ & ~new_n8240_));
  assign new_n8256_ = ~new_n8248_ & ~new_n8238_ & (~new_n8247_ | ~new_n8249_ | new_n8257_);
  assign new_n8257_ = new_n8242_ & new_n8244_ & (new_n8258_ | ~\all_features[5021]  | ~\all_features[5022]  | ~\all_features[5023] );
  assign new_n8258_ = ~\all_features[5019]  & ~\all_features[5020]  & (~\all_features[5018]  | new_n8236_);
  assign new_n8259_ = ~new_n8250_ & ~new_n8252_;
  assign new_n8260_ = ~new_n8261_ & ~new_n8254_;
  assign new_n8261_ = ~new_n8253_ & (new_n8252_ | (~new_n8250_ & (new_n8240_ | (~new_n8234_ & ~new_n8262_))));
  assign new_n8262_ = ~new_n8238_ & (new_n8248_ | (new_n8247_ & (~new_n8249_ | (~new_n8263_ & new_n8242_))));
  assign new_n8263_ = ~\all_features[5021]  & \all_features[5022]  & \all_features[5023]  & (\all_features[5020]  ? new_n8246_ : (new_n8245_ | ~new_n8246_));
  assign new_n8264_ = new_n8259_ & new_n8237_ & ~new_n8254_ & ~new_n8248_ & ~new_n8234_ & ~new_n8253_;
  assign new_n8265_ = ~new_n8030_ & new_n7956_;
  assign new_n8266_ = (~new_n8344_ & (new_n8298_ | ~new_n8346_)) ? ~new_n8327_ : new_n8267_;
  assign new_n8267_ = ~new_n8295_ & new_n8268_;
  assign new_n8268_ = ~new_n8269_ & ~new_n8292_;
  assign new_n8269_ = new_n8270_ & (new_n8289_ | new_n8290_ | ~new_n8285_ | (new_n8282_ & new_n8280_));
  assign new_n8270_ = new_n8271_ & new_n8277_;
  assign new_n8271_ = ~new_n8272_ & ~new_n8275_;
  assign new_n8272_ = ~\all_features[3206]  & ~\all_features[3207]  & (~\all_features[3203]  | ~new_n8274_ | (~\all_features[3202]  & ~new_n8273_));
  assign new_n8273_ = \all_features[3200]  & \all_features[3201] ;
  assign new_n8274_ = \all_features[3204]  & \all_features[3205] ;
  assign new_n8275_ = ~\all_features[3207]  & ~new_n8276_ & ~\all_features[3206] ;
  assign new_n8276_ = \all_features[3205]  & (\all_features[3204]  | (\all_features[3203]  & (\all_features[3202]  | \all_features[3201] )));
  assign new_n8277_ = ~new_n8279_ | (\all_features[3203]  & \all_features[3204]  & (\all_features[3202]  | ~new_n8278_));
  assign new_n8278_ = ~\all_features[3200]  & ~\all_features[3201] ;
  assign new_n8279_ = ~\all_features[3207]  & ~\all_features[3205]  & ~\all_features[3206] ;
  assign new_n8280_ = \all_features[3207]  & (\all_features[3206]  | (~new_n8281_ & \all_features[3205] ));
  assign new_n8281_ = new_n8278_ & ~\all_features[3204]  & ~\all_features[3202]  & ~\all_features[3203] ;
  assign new_n8282_ = \all_features[3207]  & \all_features[3206]  & ~new_n8284_ & new_n8283_;
  assign new_n8283_ = \all_features[3207]  & (\all_features[3206]  | (new_n8274_ & (\all_features[3202]  | \all_features[3203]  | \all_features[3201] )));
  assign new_n8284_ = ~\all_features[3205]  & ~\all_features[3204]  & ~\all_features[3203]  & ~new_n8273_ & ~\all_features[3202] ;
  assign new_n8285_ = ~new_n8286_ & ~new_n8288_;
  assign new_n8286_ = ~\all_features[3207]  & (~\all_features[3206]  | (~\all_features[3204]  & ~\all_features[3205]  & ~new_n8287_));
  assign new_n8287_ = \all_features[3202]  & \all_features[3203] ;
  assign new_n8288_ = ~\all_features[3207]  & (~\all_features[3206]  | ~new_n8273_ | ~new_n8274_ | ~new_n8287_);
  assign new_n8289_ = ~\all_features[3207]  & (~\all_features[3206]  | (~\all_features[3205]  & (new_n8278_ | ~new_n8287_ | ~\all_features[3204] )));
  assign new_n8290_ = ~new_n8291_ & ~\all_features[3207] ;
  assign new_n8291_ = \all_features[3205]  & \all_features[3206]  & (\all_features[3204]  | (\all_features[3202]  & \all_features[3203]  & \all_features[3201] ));
  assign new_n8292_ = new_n8294_ & new_n8270_ & new_n8293_;
  assign new_n8293_ = ~new_n8286_ & ~new_n8289_;
  assign new_n8294_ = ~new_n8288_ & ~new_n8290_;
  assign new_n8295_ = new_n8277_ & (~new_n8271_ | (new_n8293_ & (~new_n8294_ | new_n8296_)));
  assign new_n8296_ = new_n8280_ & (~new_n8282_ | (~new_n8297_ & \all_features[3205]  & \all_features[3206]  & \all_features[3207] ));
  assign new_n8297_ = ~\all_features[3203]  & ~\all_features[3204]  & (~\all_features[3202]  | new_n8278_);
  assign new_n8298_ = ~new_n8299_ & ~new_n8320_;
  assign new_n8299_ = ~new_n8300_ & (\all_features[2355]  | \all_features[2356]  | \all_features[2357]  | \all_features[2358]  | \all_features[2359] );
  assign new_n8300_ = ~new_n8316_ & (new_n8314_ | (~new_n8318_ & (new_n8319_ | (~new_n8317_ & ~new_n8301_))));
  assign new_n8301_ = ~new_n8302_ & (new_n8304_ | (new_n8313_ & (~new_n8308_ | (~new_n8312_ & new_n8311_))));
  assign new_n8302_ = ~new_n8303_ & ~\all_features[2359] ;
  assign new_n8303_ = \all_features[2357]  & \all_features[2358]  & (\all_features[2356]  | (\all_features[2354]  & \all_features[2355]  & \all_features[2353] ));
  assign new_n8304_ = ~\all_features[2359]  & (~\all_features[2358]  | ~new_n8305_ | ~new_n8306_ | ~new_n8307_);
  assign new_n8305_ = \all_features[2354]  & \all_features[2355] ;
  assign new_n8306_ = \all_features[2352]  & \all_features[2353] ;
  assign new_n8307_ = \all_features[2356]  & \all_features[2357] ;
  assign new_n8308_ = \all_features[2359]  & (\all_features[2358]  | (\all_features[2357]  & (\all_features[2356]  | ~new_n8310_ | ~new_n8309_)));
  assign new_n8309_ = ~\all_features[2352]  & ~\all_features[2353] ;
  assign new_n8310_ = ~\all_features[2354]  & ~\all_features[2355] ;
  assign new_n8311_ = \all_features[2359]  & (\all_features[2358]  | (new_n8307_ & (\all_features[2354]  | \all_features[2355]  | \all_features[2353] )));
  assign new_n8312_ = ~\all_features[2357]  & \all_features[2358]  & \all_features[2359]  & (\all_features[2356]  ? new_n8310_ : (new_n8306_ | ~new_n8310_));
  assign new_n8313_ = \all_features[2359]  & (\all_features[2357]  | \all_features[2358]  | \all_features[2356] );
  assign new_n8314_ = new_n8315_ & (~\all_features[2357]  | (~\all_features[2356]  & (~\all_features[2355]  | (~\all_features[2354]  & ~\all_features[2353] ))));
  assign new_n8315_ = ~\all_features[2358]  & ~\all_features[2359] ;
  assign new_n8316_ = ~\all_features[2357]  & new_n8315_ & ((~\all_features[2354]  & new_n8309_) | ~\all_features[2356]  | ~\all_features[2355] );
  assign new_n8317_ = ~\all_features[2359]  & (~\all_features[2358]  | (~\all_features[2357]  & (new_n8309_ | ~new_n8305_ | ~\all_features[2356] )));
  assign new_n8318_ = new_n8315_ & (~\all_features[2355]  | ~new_n8307_ | (~\all_features[2354]  & ~new_n8306_));
  assign new_n8319_ = ~\all_features[2359]  & (~\all_features[2358]  | (~\all_features[2356]  & ~\all_features[2357]  & ~new_n8305_));
  assign new_n8320_ = new_n8325_ & (~new_n8326_ | (~new_n8321_ & ~new_n8317_ & ~new_n8319_));
  assign new_n8321_ = ~new_n8302_ & ~new_n8304_ & (~new_n8313_ | ~new_n8308_ | new_n8322_);
  assign new_n8322_ = new_n8311_ & new_n8323_ & (new_n8324_ | ~\all_features[2357]  | ~\all_features[2358]  | ~\all_features[2359] );
  assign new_n8323_ = \all_features[2358]  & \all_features[2359]  & (\all_features[2356]  | \all_features[2357]  | new_n8306_ | ~new_n8310_);
  assign new_n8324_ = ~\all_features[2355]  & ~\all_features[2356]  & (~\all_features[2354]  | new_n8309_);
  assign new_n8325_ = ~new_n8316_ & (\all_features[2355]  | \all_features[2356]  | \all_features[2357]  | \all_features[2358]  | \all_features[2359] );
  assign new_n8326_ = ~new_n8314_ & ~new_n8318_;
  assign new_n8327_ = new_n8334_ & new_n8328_ & ~new_n8343_ & ~new_n8341_ & ~new_n8338_ & ~new_n8340_;
  assign new_n8328_ = ~new_n8329_ & ~new_n8333_;
  assign new_n8329_ = ~\all_features[3335]  & (~\all_features[3334]  | ~new_n8330_ | ~new_n8331_ | ~new_n8332_);
  assign new_n8330_ = \all_features[3328]  & \all_features[3329] ;
  assign new_n8331_ = \all_features[3332]  & \all_features[3333] ;
  assign new_n8332_ = \all_features[3330]  & \all_features[3331] ;
  assign new_n8333_ = ~\all_features[3335]  & ~\all_features[3334]  & ~\all_features[3333]  & ~\all_features[3331]  & ~\all_features[3332] ;
  assign new_n8334_ = ~new_n8335_ & ~new_n8337_;
  assign new_n8335_ = new_n8336_ & (~\all_features[3331]  | ~new_n8331_ | (~\all_features[3330]  & ~new_n8330_));
  assign new_n8336_ = ~\all_features[3334]  & ~\all_features[3335] ;
  assign new_n8337_ = new_n8336_ & (~\all_features[3333]  | (~\all_features[3332]  & (~\all_features[3331]  | (~\all_features[3330]  & ~\all_features[3329] ))));
  assign new_n8338_ = ~new_n8339_ & ~\all_features[3335] ;
  assign new_n8339_ = \all_features[3333]  & \all_features[3334]  & (\all_features[3332]  | (\all_features[3330]  & \all_features[3331]  & \all_features[3329] ));
  assign new_n8340_ = ~\all_features[3335]  & (~\all_features[3334]  | (~\all_features[3332]  & ~\all_features[3333]  & ~new_n8332_));
  assign new_n8341_ = ~\all_features[3333]  & new_n8336_ & ((~\all_features[3330]  & new_n8342_) | ~\all_features[3332]  | ~\all_features[3331] );
  assign new_n8342_ = ~\all_features[3328]  & ~\all_features[3329] ;
  assign new_n8343_ = ~\all_features[3335]  & (~\all_features[3334]  | (~\all_features[3333]  & (new_n8342_ | ~\all_features[3332]  | ~new_n8332_)));
  assign new_n8344_ = new_n8345_ & new_n8325_ & ~new_n8318_ & ~new_n8317_ & ~new_n8302_ & ~new_n8314_;
  assign new_n8345_ = ~new_n8304_ & ~new_n8319_;
  assign new_n8346_ = new_n8325_ & new_n8326_ & (new_n8347_ | new_n8302_ | new_n8317_ | ~new_n8345_);
  assign new_n8347_ = new_n8313_ & new_n8323_ & new_n8308_ & new_n8311_;
  assign new_n8348_ = new_n8349_ & (~new_n8266_ | ~new_n8265_) & (~new_n8162_ | new_n8164_);
  assign new_n8349_ = (new_n8098_ | ~new_n8029_ | ~new_n8060_) & (~new_n8163_ | (new_n8231_ & new_n8200_));
  assign new_n8350_ = ~new_n8351_ & new_n8536_;
  assign new_n8351_ = ~new_n8480_ & new_n8352_ & (~new_n8506_ | ~new_n8479_);
  assign new_n8352_ = new_n8353_ & (~new_n8476_ | (new_n8477_ & new_n7866_) | (~new_n6638_ & ~new_n7866_));
  assign new_n8353_ = (new_n8446_ | ~new_n8407_) & (~new_n8354_ | ~new_n8410_);
  assign new_n8354_ = new_n8355_ & ~new_n8391_ & new_n8390_;
  assign new_n8355_ = ~new_n8388_ & (~new_n8385_ | ~new_n8356_);
  assign new_n8356_ = new_n8357_ & new_n8381_;
  assign new_n8357_ = ~new_n8379_ & ~new_n8378_ & (~new_n8372_ | (~new_n8358_ & ~new_n8376_ & ~new_n8380_));
  assign new_n8358_ = ~new_n8367_ & ~new_n8369_ & (~new_n8371_ | ~new_n8370_ | new_n8359_);
  assign new_n8359_ = new_n8360_ & new_n8362_ & (new_n8365_ | ~\all_features[4325]  | ~\all_features[4326]  | ~\all_features[4327] );
  assign new_n8360_ = \all_features[4327]  & (\all_features[4326]  | (new_n8361_ & (\all_features[4322]  | \all_features[4323]  | \all_features[4321] )));
  assign new_n8361_ = \all_features[4324]  & \all_features[4325] ;
  assign new_n8362_ = \all_features[4326]  & \all_features[4327]  & (\all_features[4324]  | \all_features[4325]  | new_n8363_ | ~new_n8364_);
  assign new_n8363_ = \all_features[4320]  & \all_features[4321] ;
  assign new_n8364_ = ~\all_features[4322]  & ~\all_features[4323] ;
  assign new_n8365_ = ~\all_features[4323]  & ~\all_features[4324]  & (~\all_features[4322]  | new_n8366_);
  assign new_n8366_ = ~\all_features[4320]  & ~\all_features[4321] ;
  assign new_n8367_ = ~new_n8368_ & ~\all_features[4327] ;
  assign new_n8368_ = \all_features[4325]  & \all_features[4326]  & (\all_features[4324]  | (\all_features[4322]  & \all_features[4323]  & \all_features[4321] ));
  assign new_n8369_ = ~\all_features[4327]  & (~new_n8361_ | ~\all_features[4322]  | ~\all_features[4323]  | ~\all_features[4326]  | ~new_n8363_);
  assign new_n8370_ = \all_features[4327]  & (\all_features[4326]  | (\all_features[4325]  & (\all_features[4324]  | ~new_n8364_ | ~new_n8366_)));
  assign new_n8371_ = \all_features[4327]  & (\all_features[4325]  | \all_features[4326]  | \all_features[4324] );
  assign new_n8372_ = ~new_n8373_ & ~new_n8375_;
  assign new_n8373_ = new_n8374_ & (~\all_features[4323]  | ~new_n8361_ | (~\all_features[4322]  & ~new_n8363_));
  assign new_n8374_ = ~\all_features[4326]  & ~\all_features[4327] ;
  assign new_n8375_ = new_n8374_ & (~\all_features[4325]  | (~\all_features[4324]  & (~\all_features[4323]  | (~\all_features[4322]  & ~\all_features[4321] ))));
  assign new_n8376_ = ~\all_features[4327]  & (~\all_features[4326]  | new_n8377_);
  assign new_n8377_ = ~\all_features[4325]  & (new_n8366_ | ~\all_features[4323]  | ~\all_features[4324]  | ~\all_features[4322] );
  assign new_n8378_ = ~\all_features[4325]  & new_n8374_ & ((~\all_features[4322]  & new_n8366_) | ~\all_features[4324]  | ~\all_features[4323] );
  assign new_n8379_ = ~\all_features[4327]  & ~\all_features[4326]  & ~\all_features[4325]  & ~\all_features[4323]  & ~\all_features[4324] ;
  assign new_n8380_ = ~\all_features[4327]  & (~\all_features[4326]  | (~\all_features[4325]  & ~\all_features[4324]  & (~\all_features[4323]  | ~\all_features[4322] )));
  assign new_n8381_ = ~new_n8382_ & ~new_n8379_;
  assign new_n8382_ = ~new_n8378_ & (new_n8375_ | (~new_n8373_ & (new_n8380_ | (~new_n8376_ & ~new_n8383_))));
  assign new_n8383_ = ~new_n8367_ & (new_n8369_ | (new_n8371_ & (~new_n8370_ | (~new_n8384_ & new_n8360_))));
  assign new_n8384_ = ~\all_features[4325]  & \all_features[4326]  & \all_features[4327]  & (\all_features[4324]  ? new_n8364_ : (new_n8363_ | ~new_n8364_));
  assign new_n8385_ = ~new_n8379_ & ~new_n8375_ & ~new_n8373_ & ~new_n8386_ & ~new_n8378_;
  assign new_n8386_ = ~new_n8380_ & ~new_n8369_ & ~new_n8367_ & ~new_n8376_ & ~new_n8387_;
  assign new_n8387_ = new_n8371_ & new_n8362_ & new_n8370_ & new_n8360_;
  assign new_n8388_ = new_n8372_ & new_n8389_ & ~new_n8380_ & ~new_n8378_ & ~new_n8376_ & ~new_n8367_;
  assign new_n8389_ = ~new_n8369_ & ~new_n8379_;
  assign new_n8390_ = new_n6424_ & new_n6411_ & new_n6421_;
  assign new_n8391_ = new_n8396_ & new_n8392_ & ~new_n8406_ & ~new_n8405_ & ~new_n8402_ & ~new_n8404_;
  assign new_n8392_ = ~new_n8393_ & (\all_features[1419]  | \all_features[1420]  | \all_features[1421]  | \all_features[1422]  | \all_features[1423] );
  assign new_n8393_ = ~\all_features[1421]  & new_n8394_ & ((~\all_features[1418]  & new_n8395_) | ~\all_features[1420]  | ~\all_features[1419] );
  assign new_n8394_ = ~\all_features[1422]  & ~\all_features[1423] ;
  assign new_n8395_ = ~\all_features[1416]  & ~\all_features[1417] ;
  assign new_n8396_ = ~new_n8397_ & ~new_n8401_;
  assign new_n8397_ = ~\all_features[1423]  & (~\all_features[1422]  | ~new_n8398_ | ~new_n8399_ | ~new_n8400_);
  assign new_n8398_ = \all_features[1418]  & \all_features[1419] ;
  assign new_n8399_ = \all_features[1416]  & \all_features[1417] ;
  assign new_n8400_ = \all_features[1420]  & \all_features[1421] ;
  assign new_n8401_ = ~\all_features[1423]  & (~\all_features[1422]  | (~\all_features[1420]  & ~\all_features[1421]  & ~new_n8398_));
  assign new_n8402_ = ~new_n8403_ & ~\all_features[1423] ;
  assign new_n8403_ = \all_features[1421]  & \all_features[1422]  & (\all_features[1420]  | (\all_features[1418]  & \all_features[1419]  & \all_features[1417] ));
  assign new_n8404_ = new_n8394_ & (~\all_features[1421]  | (~\all_features[1420]  & (~\all_features[1419]  | (~\all_features[1418]  & ~\all_features[1417] ))));
  assign new_n8405_ = ~\all_features[1423]  & (~\all_features[1422]  | (~\all_features[1421]  & (new_n8395_ | ~new_n8398_ | ~\all_features[1420] )));
  assign new_n8406_ = new_n8394_ & (~\all_features[1419]  | ~new_n8400_ | (~\all_features[1418]  & ~new_n8399_));
  assign new_n8407_ = ~new_n8408_ & new_n8391_;
  assign new_n8408_ = new_n7946_ & (new_n7943_ | ~new_n8409_);
  assign new_n8409_ = ~new_n7914_ & ~new_n7935_;
  assign new_n8410_ = new_n8411_ & new_n8437_;
  assign new_n8411_ = new_n8412_ & new_n8434_;
  assign new_n8412_ = ~new_n8433_ & ~new_n8432_ & ~new_n8431_ & ~new_n8413_ & ~new_n8429_;
  assign new_n8413_ = new_n8414_ & (~new_n8427_ | ~new_n8428_ | ~new_n8424_ | ~new_n8426_);
  assign new_n8414_ = ~new_n8421_ & ~new_n8420_ & ~new_n8415_ & ~new_n8418_;
  assign new_n8415_ = ~\all_features[4079]  & (~\all_features[4078]  | (~\all_features[4077]  & (new_n8416_ | ~new_n8417_ | ~\all_features[4076] )));
  assign new_n8416_ = ~\all_features[4072]  & ~\all_features[4073] ;
  assign new_n8417_ = \all_features[4074]  & \all_features[4075] ;
  assign new_n8418_ = ~new_n8419_ & ~\all_features[4079] ;
  assign new_n8419_ = \all_features[4077]  & \all_features[4078]  & (\all_features[4076]  | (\all_features[4074]  & \all_features[4075]  & \all_features[4073] ));
  assign new_n8420_ = ~\all_features[4079]  & (~\all_features[4078]  | (~\all_features[4076]  & ~\all_features[4077]  & ~new_n8417_));
  assign new_n8421_ = ~\all_features[4079]  & (~\all_features[4078]  | ~new_n8422_ | ~new_n8423_ | ~new_n8417_);
  assign new_n8422_ = \all_features[4076]  & \all_features[4077] ;
  assign new_n8423_ = \all_features[4072]  & \all_features[4073] ;
  assign new_n8424_ = \all_features[4079]  & (\all_features[4078]  | (\all_features[4077]  & (\all_features[4076]  | ~new_n8416_ | ~new_n8425_)));
  assign new_n8425_ = ~\all_features[4074]  & ~\all_features[4075] ;
  assign new_n8426_ = \all_features[4079]  & (\all_features[4078]  | (new_n8422_ & (\all_features[4074]  | \all_features[4075]  | \all_features[4073] )));
  assign new_n8427_ = \all_features[4078]  & \all_features[4079]  & (\all_features[4076]  | \all_features[4077]  | new_n8423_ | ~new_n8425_);
  assign new_n8428_ = \all_features[4079]  & (\all_features[4077]  | \all_features[4078]  | \all_features[4076] );
  assign new_n8429_ = new_n8430_ & (~\all_features[4077]  | (~\all_features[4076]  & (~\all_features[4075]  | (~\all_features[4074]  & ~\all_features[4073] ))));
  assign new_n8430_ = ~\all_features[4078]  & ~\all_features[4079] ;
  assign new_n8431_ = ~\all_features[4077]  & new_n8430_ & ((~\all_features[4074]  & new_n8416_) | ~\all_features[4076]  | ~\all_features[4075] );
  assign new_n8432_ = new_n8430_ & (~\all_features[4075]  | ~new_n8422_ | (~\all_features[4074]  & ~new_n8423_));
  assign new_n8433_ = ~\all_features[4079]  & ~\all_features[4078]  & ~\all_features[4077]  & ~\all_features[4075]  & ~\all_features[4076] ;
  assign new_n8434_ = new_n8436_ & new_n8435_ & ~new_n8431_ & ~new_n8421_ & ~new_n8415_ & ~new_n8418_;
  assign new_n8435_ = ~new_n8420_ & ~new_n8433_;
  assign new_n8436_ = ~new_n8429_ & ~new_n8432_;
  assign new_n8437_ = new_n8438_ & new_n8442_;
  assign new_n8438_ = ~new_n8431_ & ~new_n8433_ & (~new_n8436_ | (~new_n8439_ & ~new_n8415_ & ~new_n8420_));
  assign new_n8439_ = ~new_n8421_ & ~new_n8418_ & (~new_n8428_ | ~new_n8424_ | new_n8440_);
  assign new_n8440_ = new_n8426_ & new_n8427_ & (new_n8441_ | ~\all_features[4077]  | ~\all_features[4078]  | ~\all_features[4079] );
  assign new_n8441_ = ~\all_features[4075]  & ~\all_features[4076]  & (~\all_features[4074]  | new_n8416_);
  assign new_n8442_ = ~new_n8443_ & ~new_n8433_;
  assign new_n8443_ = ~new_n8431_ & (new_n8429_ | (~new_n8432_ & (new_n8420_ | (~new_n8415_ & ~new_n8444_))));
  assign new_n8444_ = ~new_n8418_ & (new_n8421_ | (new_n8428_ & (~new_n8424_ | (~new_n8445_ & new_n8426_))));
  assign new_n8445_ = ~\all_features[4077]  & \all_features[4078]  & \all_features[4079]  & (\all_features[4076]  ? new_n8425_ : (new_n8423_ | ~new_n8425_));
  assign new_n8446_ = ~new_n8475_ & (~new_n8471_ | ~new_n8447_);
  assign new_n8447_ = new_n8468_ & ~new_n8448_ & new_n8464_;
  assign new_n8448_ = ~new_n8458_ & ~new_n8460_ & ~new_n8461_ & ~new_n8463_ & (~new_n8453_ | ~new_n8449_);
  assign new_n8449_ = \all_features[2511]  & (\all_features[2510]  | (~new_n8450_ & \all_features[2509] ));
  assign new_n8450_ = new_n8451_ & ~\all_features[2508]  & new_n8452_;
  assign new_n8451_ = ~\all_features[2504]  & ~\all_features[2505] ;
  assign new_n8452_ = ~\all_features[2506]  & ~\all_features[2507] ;
  assign new_n8453_ = \all_features[2511]  & \all_features[2510]  & ~new_n8456_ & new_n8454_;
  assign new_n8454_ = \all_features[2511]  & (\all_features[2510]  | (new_n8455_ & (\all_features[2506]  | \all_features[2507]  | \all_features[2505] )));
  assign new_n8455_ = \all_features[2508]  & \all_features[2509] ;
  assign new_n8456_ = new_n8452_ & ~\all_features[2509]  & ~new_n8457_ & ~\all_features[2508] ;
  assign new_n8457_ = \all_features[2504]  & \all_features[2505] ;
  assign new_n8458_ = ~\all_features[2511]  & (~\all_features[2510]  | (~\all_features[2508]  & ~\all_features[2509]  & ~new_n8459_));
  assign new_n8459_ = \all_features[2506]  & \all_features[2507] ;
  assign new_n8460_ = ~\all_features[2511]  & (~\all_features[2510]  | (~\all_features[2509]  & (new_n8451_ | ~\all_features[2508]  | ~new_n8459_)));
  assign new_n8461_ = ~new_n8462_ & ~\all_features[2511] ;
  assign new_n8462_ = \all_features[2509]  & \all_features[2510]  & (\all_features[2508]  | (\all_features[2506]  & \all_features[2507]  & \all_features[2505] ));
  assign new_n8463_ = ~\all_features[2511]  & (~\all_features[2510]  | ~new_n8459_ | ~new_n8457_ | ~new_n8455_);
  assign new_n8464_ = ~new_n8465_ & ~new_n8467_;
  assign new_n8465_ = new_n8466_ & (~\all_features[2507]  | ~new_n8455_ | (~\all_features[2506]  & ~new_n8457_));
  assign new_n8466_ = ~\all_features[2510]  & ~\all_features[2511] ;
  assign new_n8467_ = new_n8466_ & (~\all_features[2509]  | (~\all_features[2508]  & (~\all_features[2507]  | (~\all_features[2506]  & ~\all_features[2505] ))));
  assign new_n8468_ = ~new_n8469_ & ~new_n8470_;
  assign new_n8469_ = ~\all_features[2509]  & new_n8466_ & ((~\all_features[2506]  & new_n8451_) | ~\all_features[2508]  | ~\all_features[2507] );
  assign new_n8470_ = ~\all_features[2511]  & ~\all_features[2510]  & ~\all_features[2509]  & ~\all_features[2507]  & ~\all_features[2508] ;
  assign new_n8471_ = new_n8468_ & (~new_n8464_ | (new_n8474_ & (new_n8472_ | new_n8461_ | new_n8463_)));
  assign new_n8472_ = new_n8449_ & (~new_n8453_ | (~new_n8473_ & \all_features[2509]  & \all_features[2510]  & \all_features[2511] ));
  assign new_n8473_ = ~\all_features[2507]  & ~\all_features[2508]  & (~\all_features[2506]  | new_n8451_);
  assign new_n8474_ = ~new_n8458_ & ~new_n8460_;
  assign new_n8475_ = new_n8464_ & new_n8474_ & new_n8468_ & ~new_n8461_ & ~new_n8463_;
  assign new_n8476_ = new_n8408_ & new_n8391_;
  assign new_n8477_ = ~new_n8478_ & new_n6734_;
  assign new_n8478_ = ~new_n6732_ & ~new_n6723_;
  assign new_n8479_ = new_n8407_ & new_n8446_;
  assign new_n8480_ = ~new_n8391_ & ((~new_n8355_ & ~new_n7509_ & new_n8390_) | (~new_n8481_ & ~new_n8390_));
  assign new_n8481_ = ~new_n7902_ & new_n8483_ & (~new_n7899_ | ~new_n8482_);
  assign new_n8482_ = new_n7870_ & new_n7895_;
  assign new_n8483_ = new_n8505_ & new_n8503_ & new_n8502_ & new_n8500_ & new_n8484_ & new_n8493_;
  assign new_n8484_ = new_n8485_ & ~new_n8489_ & ~new_n8490_;
  assign new_n8485_ = ~new_n8486_ & (\all_features[3323]  | \all_features[3324]  | \all_features[3325]  | \all_features[3326]  | \all_features[3327] );
  assign new_n8486_ = ~\all_features[3325]  & new_n8488_ & ((~\all_features[3322]  & new_n8487_) | ~\all_features[3324]  | ~\all_features[3323] );
  assign new_n8487_ = ~\all_features[3320]  & ~\all_features[3321] ;
  assign new_n8488_ = ~\all_features[3326]  & ~\all_features[3327] ;
  assign new_n8489_ = new_n8488_ & (~\all_features[3325]  | (~\all_features[3324]  & (~\all_features[3323]  | (~\all_features[3322]  & ~\all_features[3321] ))));
  assign new_n8490_ = new_n8488_ & (~\all_features[3323]  | ~new_n8492_ | (~\all_features[3322]  & ~new_n8491_));
  assign new_n8491_ = \all_features[3320]  & \all_features[3321] ;
  assign new_n8492_ = \all_features[3324]  & \all_features[3325] ;
  assign new_n8493_ = ~new_n8499_ & ~new_n8498_ & ~new_n8494_ & ~new_n8496_;
  assign new_n8494_ = ~\all_features[3327]  & (~\all_features[3326]  | (~\all_features[3325]  & (new_n8487_ | ~\all_features[3324]  | ~new_n8495_)));
  assign new_n8495_ = \all_features[3322]  & \all_features[3323] ;
  assign new_n8496_ = ~new_n8497_ & ~\all_features[3327] ;
  assign new_n8497_ = \all_features[3325]  & \all_features[3326]  & (\all_features[3324]  | (\all_features[3322]  & \all_features[3323]  & \all_features[3321] ));
  assign new_n8498_ = ~\all_features[3327]  & (~\all_features[3326]  | ~new_n8495_ | ~new_n8491_ | ~new_n8492_);
  assign new_n8499_ = ~\all_features[3327]  & (~\all_features[3326]  | (~\all_features[3324]  & ~\all_features[3325]  & ~new_n8495_));
  assign new_n8500_ = \all_features[3327]  & (\all_features[3326]  | (\all_features[3325]  & (\all_features[3324]  | ~new_n8501_ | ~new_n8487_)));
  assign new_n8501_ = ~\all_features[3322]  & ~\all_features[3323] ;
  assign new_n8502_ = \all_features[3327]  & (\all_features[3326]  | (new_n8492_ & (\all_features[3322]  | \all_features[3323]  | \all_features[3321] )));
  assign new_n8503_ = new_n8504_ & (new_n8491_ | \all_features[3324]  | \all_features[3325]  | ~new_n8501_);
  assign new_n8504_ = \all_features[3326]  & \all_features[3327] ;
  assign new_n8505_ = \all_features[3327]  & (\all_features[3325]  | \all_features[3326]  | \all_features[3324] );
  assign new_n8506_ = ~new_n8535_ & new_n8507_;
  assign new_n8507_ = ~new_n8508_ & ~new_n8533_;
  assign new_n8508_ = new_n8509_ & (~new_n8527_ | (new_n8523_ & (new_n8515_ | new_n8530_ | new_n8532_)));
  assign new_n8509_ = ~new_n8510_ & ~new_n8514_;
  assign new_n8510_ = new_n8511_ & ((~\all_features[3082]  & new_n8513_) | ~\all_features[3084]  | ~\all_features[3083] );
  assign new_n8511_ = ~\all_features[3085]  & new_n8512_;
  assign new_n8512_ = ~\all_features[3086]  & ~\all_features[3087] ;
  assign new_n8513_ = ~\all_features[3080]  & ~\all_features[3081] ;
  assign new_n8514_ = new_n8511_ & ~\all_features[3083]  & ~\all_features[3084] ;
  assign new_n8515_ = new_n8516_ & (~new_n8518_ | (~new_n8522_ & \all_features[3085]  & \all_features[3086]  & \all_features[3087] ));
  assign new_n8516_ = \all_features[3087]  & (\all_features[3086]  | (~new_n8517_ & \all_features[3085] ));
  assign new_n8517_ = new_n8513_ & ~\all_features[3084]  & ~\all_features[3082]  & ~\all_features[3083] ;
  assign new_n8518_ = \all_features[3087]  & \all_features[3086]  & ~new_n8521_ & new_n8519_;
  assign new_n8519_ = \all_features[3087]  & (\all_features[3086]  | (new_n8520_ & (\all_features[3082]  | \all_features[3083]  | \all_features[3081] )));
  assign new_n8520_ = \all_features[3084]  & \all_features[3085] ;
  assign new_n8521_ = ~\all_features[3082]  & ~\all_features[3083]  & ~\all_features[3084]  & ~\all_features[3085]  & (~\all_features[3081]  | ~\all_features[3080] );
  assign new_n8522_ = ~\all_features[3083]  & ~\all_features[3084]  & (~\all_features[3082]  | new_n8513_);
  assign new_n8523_ = ~new_n8524_ & ~new_n8526_;
  assign new_n8524_ = ~\all_features[3087]  & (~\all_features[3086]  | (~\all_features[3084]  & ~\all_features[3085]  & ~new_n8525_));
  assign new_n8525_ = \all_features[3082]  & \all_features[3083] ;
  assign new_n8526_ = ~\all_features[3087]  & (~\all_features[3086]  | (~\all_features[3085]  & (new_n8513_ | ~\all_features[3084]  | ~new_n8525_)));
  assign new_n8527_ = ~new_n8528_ & ~new_n8529_;
  assign new_n8528_ = new_n8512_ & (~new_n8520_ | ~\all_features[3083]  | (~\all_features[3082]  & (~\all_features[3080]  | ~\all_features[3081] )));
  assign new_n8529_ = new_n8512_ & (~\all_features[3085]  | (~\all_features[3084]  & (~\all_features[3083]  | (~\all_features[3082]  & ~\all_features[3081] ))));
  assign new_n8530_ = ~new_n8531_ & ~\all_features[3087] ;
  assign new_n8531_ = \all_features[3085]  & \all_features[3086]  & (\all_features[3084]  | (\all_features[3082]  & \all_features[3083]  & \all_features[3081] ));
  assign new_n8532_ = ~\all_features[3087]  & (~new_n8520_ | ~\all_features[3080]  | ~\all_features[3081]  | ~\all_features[3086]  | ~new_n8525_);
  assign new_n8533_ = new_n8527_ & ~new_n8534_ & new_n8509_;
  assign new_n8534_ = ~new_n8524_ & ~new_n8526_ & ~new_n8530_ & ~new_n8532_ & (~new_n8518_ | ~new_n8516_);
  assign new_n8535_ = new_n8527_ & new_n8523_ & ~new_n8532_ & ~new_n8530_ & ~new_n8510_ & ~new_n8514_;
  assign new_n8536_ = new_n8537_ & (new_n8506_ | ~new_n8479_);
  assign new_n8537_ = (~new_n8354_ | new_n8410_) & (new_n6638_ | new_n7866_ | ~new_n8476_);
  assign new_n8538_ = new_n8539_ & (new_n8541_ | ~new_n8543_ | (new_n8776_ ? new_n8740_ : new_n8703_));
  assign new_n8539_ = ~new_n8540_ & (~new_n8541_ | (new_n7270_ & new_n7293_ & ~new_n8667_) | (new_n8630_ & new_n8667_));
  assign new_n8540_ = ~new_n8543_ & ~new_n8541_ & (~new_n8595_ | ~new_n8621_) & (~new_n8558_ | ~new_n8590_);
  assign new_n8541_ = new_n6869_ & new_n6849_ & new_n8542_;
  assign new_n8542_ = new_n6880_ & new_n6883_;
  assign new_n8543_ = new_n8544_ & new_n6955_;
  assign new_n8544_ = new_n8545_ & new_n8554_;
  assign new_n8545_ = new_n8553_ & ~new_n8546_ & new_n6961_;
  assign new_n8546_ = new_n8547_ & (~new_n8551_ | ~new_n8552_ | ~new_n8548_ | ~new_n8550_);
  assign new_n8547_ = ~new_n6968_ & ~new_n6969_ & ~new_n6957_ & ~new_n6959_;
  assign new_n8548_ = \all_features[4151]  & (\all_features[4150]  | (\all_features[4149]  & (\all_features[4148]  | ~new_n8549_ | ~new_n6960_)));
  assign new_n8549_ = ~\all_features[4146]  & ~\all_features[4147] ;
  assign new_n8550_ = \all_features[4151]  & (\all_features[4150]  | (new_n6965_ & (\all_features[4146]  | \all_features[4147]  | \all_features[4145] )));
  assign new_n8551_ = \all_features[4150]  & \all_features[4151]  & (\all_features[4148]  | \all_features[4149]  | new_n6964_ | ~new_n8549_);
  assign new_n8552_ = \all_features[4151]  & (\all_features[4149]  | \all_features[4150]  | \all_features[4148] );
  assign new_n8553_ = ~new_n6971_ & (\all_features[4147]  | \all_features[4148]  | \all_features[4149]  | \all_features[4150]  | \all_features[4151] );
  assign new_n8554_ = new_n8553_ & (~new_n6961_ | (new_n6956_ & (new_n8555_ | new_n6969_ | new_n6968_)));
  assign new_n8555_ = new_n8548_ & new_n8552_ & (~new_n8551_ | ~new_n8550_ | new_n8556_);
  assign new_n8556_ = \all_features[4151]  & \all_features[4150]  & ~new_n8557_ & \all_features[4149] ;
  assign new_n8557_ = ~\all_features[4147]  & ~\all_features[4148]  & (~\all_features[4146]  | new_n6960_);
  assign new_n8558_ = new_n8559_ & new_n8580_;
  assign new_n8559_ = ~new_n8560_ & (\all_features[3979]  | \all_features[3980]  | \all_features[3981]  | \all_features[3982]  | \all_features[3983] );
  assign new_n8560_ = ~new_n8574_ & (new_n8576_ | (~new_n8577_ & (new_n8578_ | (~new_n8561_ & ~new_n8579_))));
  assign new_n8561_ = ~new_n8569_ & (new_n8571_ | (~new_n8562_ & new_n8573_));
  assign new_n8562_ = \all_features[3983]  & ((~new_n8567_ & ~\all_features[3981]  & \all_features[3982] ) | (~new_n8565_ & (\all_features[3982]  | (~new_n8563_ & \all_features[3981] ))));
  assign new_n8563_ = new_n8564_ & ~\all_features[3980]  & ~\all_features[3978]  & ~\all_features[3979] ;
  assign new_n8564_ = ~\all_features[3976]  & ~\all_features[3977] ;
  assign new_n8565_ = \all_features[3983]  & (\all_features[3982]  | (new_n8566_ & (\all_features[3978]  | \all_features[3979]  | \all_features[3977] )));
  assign new_n8566_ = \all_features[3980]  & \all_features[3981] ;
  assign new_n8567_ = (\all_features[3980]  & (\all_features[3978]  | \all_features[3979] )) | (~new_n8568_ & ~\all_features[3978]  & ~\all_features[3979]  & ~\all_features[3980] );
  assign new_n8568_ = \all_features[3976]  & \all_features[3977] ;
  assign new_n8569_ = ~new_n8570_ & ~\all_features[3983] ;
  assign new_n8570_ = \all_features[3981]  & \all_features[3982]  & (\all_features[3980]  | (\all_features[3978]  & \all_features[3979]  & \all_features[3977] ));
  assign new_n8571_ = ~\all_features[3983]  & (~\all_features[3982]  | ~new_n8568_ | ~new_n8566_ | ~new_n8572_);
  assign new_n8572_ = \all_features[3978]  & \all_features[3979] ;
  assign new_n8573_ = \all_features[3983]  & (\all_features[3981]  | \all_features[3982]  | \all_features[3980] );
  assign new_n8574_ = ~\all_features[3981]  & new_n8575_ & ((~\all_features[3978]  & new_n8564_) | ~\all_features[3980]  | ~\all_features[3979] );
  assign new_n8575_ = ~\all_features[3982]  & ~\all_features[3983] ;
  assign new_n8576_ = new_n8575_ & (~\all_features[3981]  | (~\all_features[3980]  & (~\all_features[3979]  | (~\all_features[3978]  & ~\all_features[3977] ))));
  assign new_n8577_ = new_n8575_ & (~\all_features[3979]  | ~new_n8566_ | (~\all_features[3978]  & ~new_n8568_));
  assign new_n8578_ = ~\all_features[3983]  & (~\all_features[3982]  | (~\all_features[3980]  & ~\all_features[3981]  & ~new_n8572_));
  assign new_n8579_ = ~\all_features[3983]  & (~\all_features[3982]  | (~\all_features[3981]  & (new_n8564_ | ~new_n8572_ | ~\all_features[3980] )));
  assign new_n8580_ = new_n8586_ & (~new_n8587_ | (new_n8588_ & (~new_n8589_ | new_n8581_)));
  assign new_n8581_ = new_n8582_ & (~new_n8583_ | (~new_n8585_ & \all_features[3981]  & \all_features[3982]  & \all_features[3983] ));
  assign new_n8582_ = \all_features[3983]  & (\all_features[3982]  | (~new_n8563_ & \all_features[3981] ));
  assign new_n8583_ = \all_features[3983]  & \all_features[3982]  & ~new_n8584_ & new_n8565_;
  assign new_n8584_ = ~\all_features[3981]  & ~\all_features[3980]  & ~\all_features[3979]  & ~new_n8568_ & ~\all_features[3978] ;
  assign new_n8585_ = ~\all_features[3979]  & ~\all_features[3980]  & (~\all_features[3978]  | new_n8564_);
  assign new_n8586_ = ~new_n8574_ & (\all_features[3979]  | \all_features[3980]  | \all_features[3981]  | \all_features[3982]  | \all_features[3983] );
  assign new_n8587_ = ~new_n8576_ & ~new_n8577_;
  assign new_n8588_ = ~new_n8578_ & ~new_n8579_;
  assign new_n8589_ = ~new_n8569_ & ~new_n8571_;
  assign new_n8590_ = new_n8591_ & new_n8594_;
  assign new_n8591_ = new_n8592_ & (new_n8579_ | new_n8569_ | ~new_n8593_ | (new_n8583_ & new_n8582_));
  assign new_n8592_ = new_n8586_ & new_n8587_;
  assign new_n8593_ = ~new_n8578_ & ~new_n8571_;
  assign new_n8594_ = new_n8589_ & new_n8592_ & new_n8588_;
  assign new_n8595_ = ~new_n8596_ & ~new_n8619_;
  assign new_n8596_ = new_n8614_ & ~new_n8618_ & ~new_n8597_ & ~new_n8617_;
  assign new_n8597_ = ~new_n8612_ & ~new_n8613_ & new_n8605_ & (~new_n8610_ | ~new_n8598_);
  assign new_n8598_ = new_n8604_ & new_n8599_ & new_n8601_;
  assign new_n8599_ = \all_features[983]  & (\all_features[982]  | (new_n8600_ & (\all_features[978]  | \all_features[979]  | \all_features[977] )));
  assign new_n8600_ = \all_features[980]  & \all_features[981] ;
  assign new_n8601_ = \all_features[982]  & \all_features[983]  & (\all_features[980]  | \all_features[981]  | new_n8603_ | ~new_n8602_);
  assign new_n8602_ = ~\all_features[978]  & ~\all_features[979] ;
  assign new_n8603_ = \all_features[976]  & \all_features[977] ;
  assign new_n8604_ = \all_features[983]  & (\all_features[981]  | \all_features[982]  | \all_features[980] );
  assign new_n8605_ = ~new_n8606_ & ~new_n8608_;
  assign new_n8606_ = ~new_n8607_ & ~\all_features[983] ;
  assign new_n8607_ = \all_features[981]  & \all_features[982]  & (\all_features[980]  | (\all_features[978]  & \all_features[979]  & \all_features[977] ));
  assign new_n8608_ = ~\all_features[983]  & (~\all_features[982]  | (~\all_features[980]  & ~\all_features[981]  & ~new_n8609_));
  assign new_n8609_ = \all_features[978]  & \all_features[979] ;
  assign new_n8610_ = \all_features[983]  & (\all_features[982]  | (\all_features[981]  & (\all_features[980]  | ~new_n8611_ | ~new_n8602_)));
  assign new_n8611_ = ~\all_features[976]  & ~\all_features[977] ;
  assign new_n8612_ = ~\all_features[983]  & (~\all_features[982]  | (~\all_features[981]  & (new_n8611_ | ~new_n8609_ | ~\all_features[980] )));
  assign new_n8613_ = ~\all_features[983]  & (~\all_features[982]  | ~new_n8600_ | ~new_n8603_ | ~new_n8609_);
  assign new_n8614_ = ~new_n8615_ & (\all_features[979]  | \all_features[980]  | \all_features[981]  | \all_features[982]  | \all_features[983] );
  assign new_n8615_ = ~\all_features[981]  & new_n8616_ & ((~\all_features[978]  & new_n8611_) | ~\all_features[980]  | ~\all_features[979] );
  assign new_n8616_ = ~\all_features[982]  & ~\all_features[983] ;
  assign new_n8617_ = new_n8616_ & (~\all_features[981]  | (~\all_features[980]  & (~\all_features[979]  | (~\all_features[978]  & ~\all_features[977] ))));
  assign new_n8618_ = new_n8616_ & (~\all_features[979]  | ~new_n8600_ | (~\all_features[978]  & ~new_n8603_));
  assign new_n8619_ = new_n8614_ & new_n8605_ & new_n8620_ & ~new_n8612_ & ~new_n8613_;
  assign new_n8620_ = ~new_n8617_ & ~new_n8618_;
  assign new_n8621_ = ~new_n8622_ & ~new_n8626_;
  assign new_n8622_ = new_n8614_ & (~new_n8620_ | (~new_n8623_ & ~new_n8608_ & ~new_n8612_));
  assign new_n8623_ = ~new_n8613_ & ~new_n8606_ & (~new_n8604_ | ~new_n8610_ | new_n8624_);
  assign new_n8624_ = new_n8599_ & new_n8601_ & (new_n8625_ | ~\all_features[981]  | ~\all_features[982]  | ~\all_features[983] );
  assign new_n8625_ = ~\all_features[979]  & ~\all_features[980]  & (~\all_features[978]  | new_n8611_);
  assign new_n8626_ = ~new_n8627_ & (\all_features[979]  | \all_features[980]  | \all_features[981]  | \all_features[982]  | \all_features[983] );
  assign new_n8627_ = ~new_n8615_ & (new_n8617_ | (~new_n8618_ & (new_n8608_ | (~new_n8612_ & ~new_n8628_))));
  assign new_n8628_ = ~new_n8606_ & (new_n8613_ | (new_n8604_ & (~new_n8610_ | (~new_n8629_ & new_n8599_))));
  assign new_n8629_ = ~\all_features[981]  & \all_features[982]  & \all_features[983]  & (\all_features[980]  ? new_n8602_ : (new_n8603_ | ~new_n8602_));
  assign new_n8630_ = new_n8631_ & new_n8662_;
  assign new_n8631_ = new_n8632_ & new_n8652_;
  assign new_n8632_ = (new_n8633_ | (new_n8651_ & (~\all_features[4579]  | ~\all_features[4580]  | (~\all_features[4578]  & new_n8637_)))) & (~new_n8651_ | \all_features[4579]  | \all_features[4580] );
  assign new_n8633_ = ~new_n8644_ & (new_n8646_ | (~new_n8647_ & (new_n8648_ | (~new_n8634_ & ~new_n8649_))));
  assign new_n8634_ = ~new_n8642_ & (~\all_features[4583]  | new_n8635_ | (~\all_features[4580]  & ~\all_features[4581]  & ~\all_features[4582] ));
  assign new_n8635_ = \all_features[4583]  & ((~new_n8638_ & ~\all_features[4581]  & \all_features[4582] ) | (~new_n8640_ & (\all_features[4582]  | (~new_n8636_ & \all_features[4581] ))));
  assign new_n8636_ = new_n8637_ & ~\all_features[4580]  & ~\all_features[4578]  & ~\all_features[4579] ;
  assign new_n8637_ = ~\all_features[4576]  & ~\all_features[4577] ;
  assign new_n8638_ = (\all_features[4580]  & (\all_features[4578]  | \all_features[4579] )) | (~new_n8639_ & ~\all_features[4578]  & ~\all_features[4579]  & ~\all_features[4580] );
  assign new_n8639_ = \all_features[4576]  & \all_features[4577] ;
  assign new_n8640_ = \all_features[4583]  & (\all_features[4582]  | (new_n8641_ & (\all_features[4578]  | \all_features[4579]  | \all_features[4577] )));
  assign new_n8641_ = \all_features[4580]  & \all_features[4581] ;
  assign new_n8642_ = ~\all_features[4583]  & (~\all_features[4582]  | ~new_n8639_ | ~new_n8641_ | ~new_n8643_);
  assign new_n8643_ = \all_features[4578]  & \all_features[4579] ;
  assign new_n8644_ = ~\all_features[4583]  & ~new_n8645_ & ~\all_features[4582] ;
  assign new_n8645_ = \all_features[4581]  & (\all_features[4580]  | (\all_features[4579]  & (\all_features[4578]  | \all_features[4577] )));
  assign new_n8646_ = ~\all_features[4582]  & ~\all_features[4583]  & (~\all_features[4579]  | ~new_n8641_ | (~\all_features[4578]  & ~new_n8639_));
  assign new_n8647_ = ~\all_features[4583]  & (~\all_features[4582]  | (~\all_features[4580]  & ~\all_features[4581]  & ~new_n8643_));
  assign new_n8648_ = ~\all_features[4583]  & (~\all_features[4582]  | (~\all_features[4581]  & (new_n8637_ | ~new_n8643_ | ~\all_features[4580] )));
  assign new_n8649_ = ~new_n8650_ & ~\all_features[4583] ;
  assign new_n8650_ = \all_features[4581]  & \all_features[4582]  & (\all_features[4580]  | (\all_features[4578]  & \all_features[4579]  & \all_features[4577] ));
  assign new_n8651_ = ~\all_features[4583]  & ~\all_features[4581]  & ~\all_features[4582] ;
  assign new_n8652_ = new_n8661_ & (~new_n8658_ | (new_n8659_ & (~new_n8660_ | new_n8653_)));
  assign new_n8653_ = new_n8654_ & (~new_n8655_ | (~new_n8657_ & \all_features[4581]  & \all_features[4582]  & \all_features[4583] ));
  assign new_n8654_ = \all_features[4583]  & (\all_features[4582]  | (~new_n8636_ & \all_features[4581] ));
  assign new_n8655_ = \all_features[4583]  & \all_features[4582]  & ~new_n8656_ & new_n8640_;
  assign new_n8656_ = ~\all_features[4581]  & ~\all_features[4580]  & ~\all_features[4579]  & ~new_n8639_ & ~\all_features[4578] ;
  assign new_n8657_ = ~\all_features[4579]  & ~\all_features[4580]  & (~\all_features[4578]  | new_n8637_);
  assign new_n8658_ = ~new_n8644_ & ~new_n8646_;
  assign new_n8659_ = ~new_n8647_ & ~new_n8648_;
  assign new_n8660_ = ~new_n8649_ & ~new_n8642_;
  assign new_n8661_ = ~new_n8651_ | (\all_features[4579]  & \all_features[4580]  & (\all_features[4578]  | ~new_n8637_));
  assign new_n8662_ = new_n8663_ & new_n8666_;
  assign new_n8663_ = new_n8664_ & (new_n8648_ | new_n8649_ | ~new_n8665_ | (new_n8655_ & new_n8654_));
  assign new_n8664_ = new_n8658_ & new_n8661_;
  assign new_n8665_ = ~new_n8647_ & ~new_n8642_;
  assign new_n8666_ = new_n8660_ & new_n8664_ & new_n8659_;
  assign new_n8667_ = ~new_n8668_ & new_n8697_;
  assign new_n8668_ = ~new_n8669_ & ~new_n8693_;
  assign new_n8669_ = new_n8684_ & (~new_n8689_ | (~new_n8687_ & ~new_n8670_ & ~new_n8692_));
  assign new_n8670_ = ~new_n8682_ & ~new_n8680_ & (~new_n8683_ | ~new_n8679_ | new_n8671_);
  assign new_n8671_ = new_n8672_ & new_n8676_ & (new_n8674_ | ~\all_features[3933]  | ~\all_features[3934]  | ~\all_features[3935] );
  assign new_n8672_ = \all_features[3935]  & (\all_features[3934]  | (new_n8673_ & (\all_features[3930]  | \all_features[3931]  | \all_features[3929] )));
  assign new_n8673_ = \all_features[3932]  & \all_features[3933] ;
  assign new_n8674_ = ~\all_features[3931]  & ~\all_features[3932]  & (~\all_features[3930]  | new_n8675_);
  assign new_n8675_ = ~\all_features[3928]  & ~\all_features[3929] ;
  assign new_n8676_ = \all_features[3934]  & \all_features[3935]  & (\all_features[3932]  | \all_features[3933]  | new_n8678_ | ~new_n8677_);
  assign new_n8677_ = ~\all_features[3930]  & ~\all_features[3931] ;
  assign new_n8678_ = \all_features[3928]  & \all_features[3929] ;
  assign new_n8679_ = \all_features[3935]  & (\all_features[3934]  | (\all_features[3933]  & (\all_features[3932]  | ~new_n8677_ | ~new_n8675_)));
  assign new_n8680_ = ~new_n8681_ & ~\all_features[3935] ;
  assign new_n8681_ = \all_features[3933]  & \all_features[3934]  & (\all_features[3932]  | (\all_features[3930]  & \all_features[3931]  & \all_features[3929] ));
  assign new_n8682_ = ~\all_features[3935]  & (~new_n8678_ | ~\all_features[3930]  | ~\all_features[3931]  | ~\all_features[3934]  | ~new_n8673_);
  assign new_n8683_ = \all_features[3935]  & (\all_features[3933]  | \all_features[3934]  | \all_features[3932] );
  assign new_n8684_ = ~new_n8685_ & (\all_features[3931]  | \all_features[3932]  | \all_features[3933]  | \all_features[3934]  | \all_features[3935] );
  assign new_n8685_ = ~\all_features[3933]  & new_n8686_ & ((~\all_features[3930]  & new_n8675_) | ~\all_features[3932]  | ~\all_features[3931] );
  assign new_n8686_ = ~\all_features[3934]  & ~\all_features[3935] ;
  assign new_n8687_ = ~\all_features[3935]  & (~\all_features[3934]  | new_n8688_);
  assign new_n8688_ = ~\all_features[3933]  & (new_n8675_ | ~\all_features[3931]  | ~\all_features[3932]  | ~\all_features[3930] );
  assign new_n8689_ = ~new_n8690_ & ~new_n8691_;
  assign new_n8690_ = new_n8686_ & (~\all_features[3933]  | (~\all_features[3932]  & (~\all_features[3931]  | (~\all_features[3930]  & ~\all_features[3929] ))));
  assign new_n8691_ = new_n8686_ & (~\all_features[3931]  | ~new_n8673_ | (~new_n8678_ & ~\all_features[3930] ));
  assign new_n8692_ = ~\all_features[3935]  & (~\all_features[3934]  | (~\all_features[3933]  & ~\all_features[3932]  & (~\all_features[3931]  | ~\all_features[3930] )));
  assign new_n8693_ = ~new_n8694_ & (\all_features[3931]  | \all_features[3932]  | \all_features[3933]  | \all_features[3934]  | \all_features[3935] );
  assign new_n8694_ = ~new_n8685_ & (new_n8690_ | (~new_n8691_ & (new_n8692_ | (~new_n8687_ & ~new_n8695_))));
  assign new_n8695_ = ~new_n8680_ & (new_n8682_ | (new_n8683_ & (~new_n8679_ | (~new_n8696_ & new_n8672_))));
  assign new_n8696_ = ~\all_features[3933]  & \all_features[3934]  & \all_features[3935]  & (\all_features[3932]  ? new_n8677_ : (new_n8678_ | ~new_n8677_));
  assign new_n8697_ = new_n8698_ & new_n8701_;
  assign new_n8698_ = new_n8689_ & ~new_n8699_ & new_n8684_;
  assign new_n8699_ = ~new_n8692_ & ~new_n8682_ & ~new_n8680_ & ~new_n8687_ & ~new_n8700_;
  assign new_n8700_ = new_n8683_ & new_n8679_ & new_n8672_ & new_n8676_;
  assign new_n8701_ = new_n8684_ & new_n8702_ & ~new_n8680_ & ~new_n8690_;
  assign new_n8702_ = ~new_n8692_ & ~new_n8691_ & ~new_n8687_ & ~new_n8682_;
  assign new_n8703_ = new_n8704_ & new_n8735_;
  assign new_n8704_ = new_n8705_ & new_n8725_;
  assign new_n8705_ = (new_n8706_ | (new_n8724_ & (~\all_features[2827]  | ~\all_features[2828]  | (~\all_features[2826]  & new_n8710_)))) & (~new_n8724_ | \all_features[2827]  | \all_features[2828] );
  assign new_n8706_ = ~new_n8717_ & (new_n8719_ | (~new_n8720_ & (new_n8721_ | (~new_n8707_ & ~new_n8722_))));
  assign new_n8707_ = ~new_n8715_ & (~\all_features[2831]  | new_n8708_ | (~\all_features[2828]  & ~\all_features[2829]  & ~\all_features[2830] ));
  assign new_n8708_ = \all_features[2831]  & ((~new_n8711_ & ~\all_features[2829]  & \all_features[2830] ) | (~new_n8713_ & (\all_features[2830]  | (~new_n8709_ & \all_features[2829] ))));
  assign new_n8709_ = new_n8710_ & ~\all_features[2828]  & ~\all_features[2826]  & ~\all_features[2827] ;
  assign new_n8710_ = ~\all_features[2824]  & ~\all_features[2825] ;
  assign new_n8711_ = (\all_features[2828]  & (\all_features[2826]  | \all_features[2827] )) | (~new_n8712_ & ~\all_features[2826]  & ~\all_features[2827]  & ~\all_features[2828] );
  assign new_n8712_ = \all_features[2824]  & \all_features[2825] ;
  assign new_n8713_ = \all_features[2831]  & (\all_features[2830]  | (new_n8714_ & (\all_features[2826]  | \all_features[2827]  | \all_features[2825] )));
  assign new_n8714_ = \all_features[2828]  & \all_features[2829] ;
  assign new_n8715_ = ~\all_features[2831]  & (~\all_features[2830]  | ~new_n8712_ | ~new_n8714_ | ~new_n8716_);
  assign new_n8716_ = \all_features[2826]  & \all_features[2827] ;
  assign new_n8717_ = ~\all_features[2831]  & ~new_n8718_ & ~\all_features[2830] ;
  assign new_n8718_ = \all_features[2829]  & (\all_features[2828]  | (\all_features[2827]  & (\all_features[2826]  | \all_features[2825] )));
  assign new_n8719_ = ~\all_features[2830]  & ~\all_features[2831]  & (~\all_features[2827]  | ~new_n8714_ | (~\all_features[2826]  & ~new_n8712_));
  assign new_n8720_ = ~\all_features[2831]  & (~\all_features[2830]  | (~\all_features[2828]  & ~\all_features[2829]  & ~new_n8716_));
  assign new_n8721_ = ~\all_features[2831]  & (~\all_features[2830]  | (~\all_features[2829]  & (new_n8710_ | ~new_n8716_ | ~\all_features[2828] )));
  assign new_n8722_ = ~new_n8723_ & ~\all_features[2831] ;
  assign new_n8723_ = \all_features[2829]  & \all_features[2830]  & (\all_features[2828]  | (\all_features[2826]  & \all_features[2827]  & \all_features[2825] ));
  assign new_n8724_ = ~\all_features[2831]  & ~\all_features[2829]  & ~\all_features[2830] ;
  assign new_n8725_ = new_n8734_ & (~new_n8731_ | (new_n8732_ & (~new_n8733_ | new_n8726_)));
  assign new_n8726_ = new_n8727_ & (~new_n8728_ | (~new_n8730_ & \all_features[2829]  & \all_features[2830]  & \all_features[2831] ));
  assign new_n8727_ = \all_features[2831]  & (\all_features[2830]  | (~new_n8709_ & \all_features[2829] ));
  assign new_n8728_ = \all_features[2831]  & \all_features[2830]  & ~new_n8729_ & new_n8713_;
  assign new_n8729_ = ~\all_features[2829]  & ~\all_features[2828]  & ~\all_features[2827]  & ~new_n8712_ & ~\all_features[2826] ;
  assign new_n8730_ = ~\all_features[2827]  & ~\all_features[2828]  & (~\all_features[2826]  | new_n8710_);
  assign new_n8731_ = ~new_n8717_ & ~new_n8719_;
  assign new_n8732_ = ~new_n8720_ & ~new_n8721_;
  assign new_n8733_ = ~new_n8722_ & ~new_n8715_;
  assign new_n8734_ = ~new_n8724_ | (\all_features[2827]  & \all_features[2828]  & (\all_features[2826]  | ~new_n8710_));
  assign new_n8735_ = new_n8736_ & new_n8739_;
  assign new_n8736_ = new_n8737_ & (new_n8721_ | new_n8722_ | ~new_n8738_ | (new_n8728_ & new_n8727_));
  assign new_n8737_ = new_n8731_ & new_n8734_;
  assign new_n8738_ = ~new_n8720_ & ~new_n8715_;
  assign new_n8739_ = new_n8733_ & new_n8737_ & new_n8732_;
  assign new_n8740_ = ~new_n8772_ & new_n8741_;
  assign new_n8741_ = ~new_n8768_ & new_n8742_;
  assign new_n8742_ = ~new_n8743_ & ~new_n8765_;
  assign new_n8743_ = new_n8760_ & ~new_n8764_ & ~new_n8744_ & ~new_n8763_;
  assign new_n8744_ = new_n8745_ & ~new_n8753_ & (~new_n8758_ | ~new_n8759_ | ~new_n8755_ | ~new_n8757_);
  assign new_n8745_ = ~new_n8750_ & ~new_n8746_ & ~new_n8748_;
  assign new_n8746_ = ~\all_features[5079]  & (~\all_features[5078]  | (~\all_features[5076]  & ~\all_features[5077]  & ~new_n8747_));
  assign new_n8747_ = \all_features[5074]  & \all_features[5075] ;
  assign new_n8748_ = ~new_n8749_ & ~\all_features[5079] ;
  assign new_n8749_ = \all_features[5077]  & \all_features[5078]  & (\all_features[5076]  | (\all_features[5074]  & \all_features[5075]  & \all_features[5073] ));
  assign new_n8750_ = ~\all_features[5079]  & (~\all_features[5078]  | ~new_n8751_ | ~new_n8752_ | ~new_n8747_);
  assign new_n8751_ = \all_features[5072]  & \all_features[5073] ;
  assign new_n8752_ = \all_features[5076]  & \all_features[5077] ;
  assign new_n8753_ = ~\all_features[5079]  & (~\all_features[5078]  | (~\all_features[5077]  & (new_n8754_ | ~new_n8747_ | ~\all_features[5076] )));
  assign new_n8754_ = ~\all_features[5072]  & ~\all_features[5073] ;
  assign new_n8755_ = \all_features[5079]  & (\all_features[5078]  | (\all_features[5077]  & (\all_features[5076]  | ~new_n8756_ | ~new_n8754_)));
  assign new_n8756_ = ~\all_features[5074]  & ~\all_features[5075] ;
  assign new_n8757_ = \all_features[5079]  & (\all_features[5078]  | (new_n8752_ & (\all_features[5074]  | \all_features[5075]  | \all_features[5073] )));
  assign new_n8758_ = \all_features[5078]  & \all_features[5079]  & (\all_features[5076]  | \all_features[5077]  | new_n8751_ | ~new_n8756_);
  assign new_n8759_ = \all_features[5079]  & (\all_features[5077]  | \all_features[5078]  | \all_features[5076] );
  assign new_n8760_ = ~new_n8761_ & (\all_features[5075]  | \all_features[5076]  | \all_features[5077]  | \all_features[5078]  | \all_features[5079] );
  assign new_n8761_ = new_n8762_ & (~\all_features[5075]  | ~new_n8752_ | (~\all_features[5074]  & ~new_n8751_));
  assign new_n8762_ = ~\all_features[5078]  & ~\all_features[5079] ;
  assign new_n8763_ = ~\all_features[5077]  & new_n8762_ & ((~\all_features[5074]  & new_n8754_) | ~\all_features[5076]  | ~\all_features[5075] );
  assign new_n8764_ = new_n8762_ & (~\all_features[5077]  | (~\all_features[5076]  & (~\all_features[5075]  | (~\all_features[5074]  & ~\all_features[5073] ))));
  assign new_n8765_ = new_n8745_ & new_n8767_ & ~new_n8753_ & new_n8766_;
  assign new_n8766_ = ~new_n8763_ & (\all_features[5075]  | \all_features[5076]  | \all_features[5077]  | \all_features[5078]  | \all_features[5079] );
  assign new_n8767_ = ~new_n8764_ & ~new_n8761_;
  assign new_n8768_ = new_n8766_ & (~new_n8767_ | (~new_n8769_ & ~new_n8746_ & ~new_n8753_));
  assign new_n8769_ = ~new_n8748_ & ~new_n8750_ & (~new_n8759_ | ~new_n8755_ | new_n8770_);
  assign new_n8770_ = new_n8757_ & new_n8758_ & (new_n8771_ | ~\all_features[5077]  | ~\all_features[5078]  | ~\all_features[5079] );
  assign new_n8771_ = ~\all_features[5075]  & ~\all_features[5076]  & (~\all_features[5074]  | new_n8754_);
  assign new_n8772_ = ~new_n8773_ & (\all_features[5075]  | \all_features[5076]  | \all_features[5077]  | \all_features[5078]  | \all_features[5079] );
  assign new_n8773_ = ~new_n8763_ & (new_n8764_ | (~new_n8761_ & (new_n8746_ | (~new_n8774_ & ~new_n8753_))));
  assign new_n8774_ = ~new_n8748_ & (new_n8750_ | (new_n8759_ & (~new_n8755_ | (~new_n8775_ & new_n8757_))));
  assign new_n8775_ = ~\all_features[5077]  & \all_features[5078]  & \all_features[5079]  & (\all_features[5076]  ? new_n8756_ : (new_n8751_ | ~new_n8756_));
  assign new_n8776_ = new_n8777_ & new_n8806_;
  assign new_n8777_ = ~new_n8778_ & ~new_n8802_;
  assign new_n8778_ = new_n8793_ & (~new_n8798_ | (~new_n8796_ & ~new_n8779_ & ~new_n8801_));
  assign new_n8779_ = ~new_n8791_ & ~new_n8789_ & (~new_n8792_ | ~new_n8788_ | new_n8780_);
  assign new_n8780_ = new_n8781_ & new_n8783_ & (new_n8786_ | ~\all_features[5269]  | ~\all_features[5270]  | ~\all_features[5271] );
  assign new_n8781_ = \all_features[5271]  & (\all_features[5270]  | (new_n8782_ & (\all_features[5266]  | \all_features[5267]  | \all_features[5265] )));
  assign new_n8782_ = \all_features[5268]  & \all_features[5269] ;
  assign new_n8783_ = \all_features[5270]  & \all_features[5271]  & (\all_features[5268]  | \all_features[5269]  | new_n8785_ | ~new_n8784_);
  assign new_n8784_ = ~\all_features[5266]  & ~\all_features[5267] ;
  assign new_n8785_ = \all_features[5264]  & \all_features[5265] ;
  assign new_n8786_ = ~\all_features[5267]  & ~\all_features[5268]  & (~\all_features[5266]  | new_n8787_);
  assign new_n8787_ = ~\all_features[5264]  & ~\all_features[5265] ;
  assign new_n8788_ = \all_features[5271]  & (\all_features[5270]  | (\all_features[5269]  & (\all_features[5268]  | ~new_n8784_ | ~new_n8787_)));
  assign new_n8789_ = ~new_n8790_ & ~\all_features[5271] ;
  assign new_n8790_ = \all_features[5269]  & \all_features[5270]  & (\all_features[5268]  | (\all_features[5266]  & \all_features[5267]  & \all_features[5265] ));
  assign new_n8791_ = ~\all_features[5271]  & (~new_n8785_ | ~\all_features[5266]  | ~\all_features[5267]  | ~\all_features[5270]  | ~new_n8782_);
  assign new_n8792_ = \all_features[5271]  & (\all_features[5269]  | \all_features[5270]  | \all_features[5268] );
  assign new_n8793_ = ~new_n8794_ & (\all_features[5267]  | \all_features[5268]  | \all_features[5269]  | \all_features[5270]  | \all_features[5271] );
  assign new_n8794_ = ~\all_features[5269]  & new_n8795_ & ((~\all_features[5266]  & new_n8787_) | ~\all_features[5268]  | ~\all_features[5267] );
  assign new_n8795_ = ~\all_features[5270]  & ~\all_features[5271] ;
  assign new_n8796_ = ~\all_features[5271]  & (~\all_features[5270]  | new_n8797_);
  assign new_n8797_ = ~\all_features[5269]  & (new_n8787_ | ~\all_features[5267]  | ~\all_features[5268]  | ~\all_features[5266] );
  assign new_n8798_ = ~new_n8799_ & ~new_n8800_;
  assign new_n8799_ = new_n8795_ & (~\all_features[5269]  | (~\all_features[5268]  & (~\all_features[5267]  | (~\all_features[5266]  & ~\all_features[5265] ))));
  assign new_n8800_ = new_n8795_ & (~\all_features[5267]  | ~new_n8782_ | (~new_n8785_ & ~\all_features[5266] ));
  assign new_n8801_ = ~\all_features[5271]  & (~\all_features[5270]  | (~\all_features[5269]  & ~\all_features[5268]  & (~\all_features[5267]  | ~\all_features[5266] )));
  assign new_n8802_ = ~new_n8803_ & (\all_features[5267]  | \all_features[5268]  | \all_features[5269]  | \all_features[5270]  | \all_features[5271] );
  assign new_n8803_ = ~new_n8794_ & (new_n8799_ | (~new_n8800_ & (new_n8801_ | (~new_n8796_ & ~new_n8804_))));
  assign new_n8804_ = ~new_n8789_ & (new_n8791_ | (new_n8792_ & (~new_n8788_ | (~new_n8805_ & new_n8781_))));
  assign new_n8805_ = ~\all_features[5269]  & \all_features[5270]  & \all_features[5271]  & (\all_features[5268]  ? new_n8784_ : (new_n8785_ | ~new_n8784_));
  assign new_n8806_ = ~new_n8807_ & ~new_n8810_;
  assign new_n8807_ = new_n8798_ & ~new_n8808_ & new_n8793_;
  assign new_n8808_ = ~new_n8801_ & ~new_n8791_ & ~new_n8789_ & ~new_n8796_ & ~new_n8809_;
  assign new_n8809_ = new_n8792_ & new_n8788_ & new_n8781_ & new_n8783_;
  assign new_n8810_ = new_n8793_ & new_n8811_ & ~new_n8789_ & ~new_n8799_;
  assign new_n8811_ = ~new_n8801_ & ~new_n8800_ & ~new_n8796_ & ~new_n8791_;
  assign new_n8812_ = new_n8813_ ? (~new_n9608_ ^ new_n9895_) : (new_n9608_ ^ new_n9895_);
  assign new_n8813_ = new_n8814_ ? (new_n9061_ ^ new_n9383_) : (~new_n9061_ ^ new_n9383_);
  assign new_n8814_ = ~new_n8815_ & new_n9059_;
  assign new_n8815_ = ~new_n8990_ & new_n8816_;
  assign new_n8816_ = (~new_n8928_ & ~new_n8889_ & (new_n8892_ ? ~new_n8891_ : ~new_n8961_)) | (~new_n8817_ & new_n8889_);
  assign new_n8817_ = new_n7407_ & ~new_n8855_ & new_n8818_;
  assign new_n8818_ = new_n8819_ & ~new_n8851_ & ~new_n8854_;
  assign new_n8819_ = ~new_n8820_ & ~new_n8841_;
  assign new_n8820_ = ~new_n8821_ & (\all_features[3275]  | \all_features[3276]  | \all_features[3277]  | \all_features[3278]  | \all_features[3279] );
  assign new_n8821_ = ~new_n8835_ & (new_n8837_ | (~new_n8838_ & (new_n8839_ | (~new_n8822_ & ~new_n8840_))));
  assign new_n8822_ = ~new_n8830_ & (new_n8832_ | (~new_n8823_ & new_n8834_));
  assign new_n8823_ = \all_features[3279]  & ((~new_n8828_ & ~\all_features[3277]  & \all_features[3278] ) | (~new_n8826_ & (\all_features[3278]  | (~new_n8824_ & \all_features[3277] ))));
  assign new_n8824_ = new_n8825_ & ~\all_features[3276]  & ~\all_features[3274]  & ~\all_features[3275] ;
  assign new_n8825_ = ~\all_features[3272]  & ~\all_features[3273] ;
  assign new_n8826_ = \all_features[3279]  & (\all_features[3278]  | (new_n8827_ & (\all_features[3274]  | \all_features[3275]  | \all_features[3273] )));
  assign new_n8827_ = \all_features[3276]  & \all_features[3277] ;
  assign new_n8828_ = (\all_features[3276]  & (\all_features[3274]  | \all_features[3275] )) | (~new_n8829_ & ~\all_features[3274]  & ~\all_features[3275]  & ~\all_features[3276] );
  assign new_n8829_ = \all_features[3272]  & \all_features[3273] ;
  assign new_n8830_ = ~new_n8831_ & ~\all_features[3279] ;
  assign new_n8831_ = \all_features[3277]  & \all_features[3278]  & (\all_features[3276]  | (\all_features[3274]  & \all_features[3275]  & \all_features[3273] ));
  assign new_n8832_ = ~\all_features[3279]  & (~\all_features[3278]  | ~new_n8829_ | ~new_n8827_ | ~new_n8833_);
  assign new_n8833_ = \all_features[3274]  & \all_features[3275] ;
  assign new_n8834_ = \all_features[3279]  & (\all_features[3277]  | \all_features[3278]  | \all_features[3276] );
  assign new_n8835_ = ~\all_features[3277]  & new_n8836_ & ((~\all_features[3274]  & new_n8825_) | ~\all_features[3276]  | ~\all_features[3275] );
  assign new_n8836_ = ~\all_features[3278]  & ~\all_features[3279] ;
  assign new_n8837_ = new_n8836_ & (~\all_features[3277]  | (~\all_features[3276]  & (~\all_features[3275]  | (~\all_features[3274]  & ~\all_features[3273] ))));
  assign new_n8838_ = new_n8836_ & (~\all_features[3275]  | ~new_n8827_ | (~\all_features[3274]  & ~new_n8829_));
  assign new_n8839_ = ~\all_features[3279]  & (~\all_features[3278]  | (~\all_features[3276]  & ~\all_features[3277]  & ~new_n8833_));
  assign new_n8840_ = ~\all_features[3279]  & (~\all_features[3278]  | (~\all_features[3277]  & (new_n8825_ | ~new_n8833_ | ~\all_features[3276] )));
  assign new_n8841_ = new_n8847_ & (~new_n8848_ | (new_n8849_ & (~new_n8850_ | new_n8842_)));
  assign new_n8842_ = new_n8843_ & (~new_n8844_ | (~new_n8846_ & \all_features[3277]  & \all_features[3278]  & \all_features[3279] ));
  assign new_n8843_ = \all_features[3279]  & (\all_features[3278]  | (~new_n8824_ & \all_features[3277] ));
  assign new_n8844_ = \all_features[3279]  & \all_features[3278]  & ~new_n8845_ & new_n8826_;
  assign new_n8845_ = ~\all_features[3277]  & ~\all_features[3276]  & ~\all_features[3275]  & ~new_n8829_ & ~\all_features[3274] ;
  assign new_n8846_ = ~\all_features[3275]  & ~\all_features[3276]  & (~\all_features[3274]  | new_n8825_);
  assign new_n8847_ = ~new_n8835_ & (\all_features[3275]  | \all_features[3276]  | \all_features[3277]  | \all_features[3278]  | \all_features[3279] );
  assign new_n8848_ = ~new_n8837_ & ~new_n8838_;
  assign new_n8849_ = ~new_n8839_ & ~new_n8840_;
  assign new_n8850_ = ~new_n8830_ & ~new_n8832_;
  assign new_n8851_ = new_n8852_ & (new_n8840_ | new_n8830_ | ~new_n8853_ | (new_n8844_ & new_n8843_));
  assign new_n8852_ = new_n8847_ & new_n8848_;
  assign new_n8853_ = ~new_n8839_ & ~new_n8832_;
  assign new_n8854_ = new_n8850_ & new_n8852_ & new_n8849_;
  assign new_n8855_ = new_n8856_ & ~new_n8881_ & ~new_n8885_;
  assign new_n8856_ = ~new_n8857_ & ~new_n8879_;
  assign new_n8857_ = new_n8874_ & ~new_n8878_ & ~new_n8858_ & ~new_n8877_;
  assign new_n8858_ = new_n8859_ & (~new_n8872_ | ~new_n8873_ | ~new_n8869_ | ~new_n8871_);
  assign new_n8859_ = ~new_n8866_ & ~new_n8864_ & ~new_n8860_ & ~new_n8862_;
  assign new_n8860_ = ~\all_features[4095]  & (~\all_features[4094]  | (~\all_features[4092]  & ~\all_features[4093]  & ~new_n8861_));
  assign new_n8861_ = \all_features[4090]  & \all_features[4091] ;
  assign new_n8862_ = ~\all_features[4095]  & (~\all_features[4094]  | (~\all_features[4093]  & (new_n8863_ | ~new_n8861_ | ~\all_features[4092] )));
  assign new_n8863_ = ~\all_features[4088]  & ~\all_features[4089] ;
  assign new_n8864_ = ~new_n8865_ & ~\all_features[4095] ;
  assign new_n8865_ = \all_features[4093]  & \all_features[4094]  & (\all_features[4092]  | (\all_features[4090]  & \all_features[4091]  & \all_features[4089] ));
  assign new_n8866_ = ~\all_features[4095]  & (~\all_features[4094]  | ~new_n8867_ | ~new_n8868_ | ~new_n8861_);
  assign new_n8867_ = \all_features[4088]  & \all_features[4089] ;
  assign new_n8868_ = \all_features[4092]  & \all_features[4093] ;
  assign new_n8869_ = \all_features[4095]  & (\all_features[4094]  | (\all_features[4093]  & (\all_features[4092]  | ~new_n8870_ | ~new_n8863_)));
  assign new_n8870_ = ~\all_features[4090]  & ~\all_features[4091] ;
  assign new_n8871_ = \all_features[4095]  & (\all_features[4094]  | (new_n8868_ & (\all_features[4090]  | \all_features[4091]  | \all_features[4089] )));
  assign new_n8872_ = \all_features[4094]  & \all_features[4095]  & (\all_features[4092]  | \all_features[4093]  | new_n8867_ | ~new_n8870_);
  assign new_n8873_ = \all_features[4095]  & (\all_features[4093]  | \all_features[4094]  | \all_features[4092] );
  assign new_n8874_ = ~new_n8875_ & (\all_features[4091]  | \all_features[4092]  | \all_features[4093]  | \all_features[4094]  | \all_features[4095] );
  assign new_n8875_ = ~\all_features[4093]  & new_n8876_ & ((~\all_features[4090]  & new_n8863_) | ~\all_features[4092]  | ~\all_features[4091] );
  assign new_n8876_ = ~\all_features[4094]  & ~\all_features[4095] ;
  assign new_n8877_ = new_n8876_ & (~\all_features[4093]  | (~\all_features[4092]  & (~\all_features[4091]  | (~\all_features[4090]  & ~\all_features[4089] ))));
  assign new_n8878_ = new_n8876_ & (~\all_features[4091]  | ~new_n8868_ | (~\all_features[4090]  & ~new_n8867_));
  assign new_n8879_ = new_n8880_ & new_n8874_ & ~new_n8877_ & ~new_n8864_;
  assign new_n8880_ = ~new_n8866_ & ~new_n8862_ & ~new_n8878_ & ~new_n8860_;
  assign new_n8881_ = ~new_n8882_ & (\all_features[4091]  | \all_features[4092]  | \all_features[4093]  | \all_features[4094]  | \all_features[4095] );
  assign new_n8882_ = ~new_n8875_ & (new_n8877_ | (~new_n8878_ & (new_n8860_ | (~new_n8883_ & ~new_n8862_))));
  assign new_n8883_ = ~new_n8864_ & (new_n8866_ | (new_n8873_ & (~new_n8869_ | (~new_n8884_ & new_n8871_))));
  assign new_n8884_ = ~\all_features[4093]  & \all_features[4094]  & \all_features[4095]  & (\all_features[4092]  ? new_n8870_ : (new_n8867_ | ~new_n8870_));
  assign new_n8885_ = new_n8874_ & (new_n8878_ | new_n8877_ | (~new_n8886_ & ~new_n8860_ & ~new_n8862_));
  assign new_n8886_ = ~new_n8864_ & ~new_n8866_ & (~new_n8873_ | ~new_n8869_ | new_n8887_);
  assign new_n8887_ = new_n8871_ & new_n8872_ & (new_n8888_ | ~\all_features[4093]  | ~\all_features[4094]  | ~\all_features[4095] );
  assign new_n8888_ = ~\all_features[4091]  & ~\all_features[4092]  & (~\all_features[4090]  | new_n8863_);
  assign new_n8889_ = new_n7327_ & (new_n7305_ | new_n8890_);
  assign new_n8890_ = new_n7330_ & new_n7334_;
  assign new_n8891_ = new_n7946_ & (new_n7943_ | new_n7913_);
  assign new_n8892_ = new_n8893_ & new_n8923_;
  assign new_n8893_ = ~new_n8894_ & ~new_n8915_;
  assign new_n8894_ = ~new_n8895_ & (\all_features[2563]  | \all_features[2564]  | \all_features[2565]  | \all_features[2566]  | \all_features[2567] );
  assign new_n8895_ = ~new_n8909_ & (new_n8914_ | (~new_n8911_ & (new_n8912_ | (~new_n8913_ & ~new_n8896_))));
  assign new_n8896_ = ~new_n8897_ & (new_n8906_ | (new_n8908_ & (~new_n8899_ | (~new_n8904_ & new_n8902_))));
  assign new_n8897_ = ~new_n8898_ & ~\all_features[2567] ;
  assign new_n8898_ = \all_features[2565]  & \all_features[2566]  & (\all_features[2564]  | (\all_features[2562]  & \all_features[2563]  & \all_features[2561] ));
  assign new_n8899_ = \all_features[2567]  & (\all_features[2566]  | (\all_features[2565]  & (\all_features[2564]  | ~new_n8901_ | ~new_n8900_)));
  assign new_n8900_ = ~\all_features[2560]  & ~\all_features[2561] ;
  assign new_n8901_ = ~\all_features[2562]  & ~\all_features[2563] ;
  assign new_n8902_ = \all_features[2567]  & (\all_features[2566]  | (new_n8903_ & (\all_features[2562]  | \all_features[2563]  | \all_features[2561] )));
  assign new_n8903_ = \all_features[2564]  & \all_features[2565] ;
  assign new_n8904_ = ~\all_features[2565]  & \all_features[2566]  & \all_features[2567]  & (\all_features[2564]  ? new_n8901_ : (new_n8905_ | ~new_n8901_));
  assign new_n8905_ = \all_features[2560]  & \all_features[2561] ;
  assign new_n8906_ = ~\all_features[2567]  & (~\all_features[2566]  | ~new_n8905_ | ~new_n8903_ | ~new_n8907_);
  assign new_n8907_ = \all_features[2562]  & \all_features[2563] ;
  assign new_n8908_ = \all_features[2567]  & (\all_features[2565]  | \all_features[2566]  | \all_features[2564] );
  assign new_n8909_ = ~\all_features[2565]  & new_n8910_ & ((~\all_features[2562]  & new_n8900_) | ~\all_features[2564]  | ~\all_features[2563] );
  assign new_n8910_ = ~\all_features[2566]  & ~\all_features[2567] ;
  assign new_n8911_ = new_n8910_ & (~\all_features[2563]  | ~new_n8903_ | (~\all_features[2562]  & ~new_n8905_));
  assign new_n8912_ = ~\all_features[2567]  & (~\all_features[2566]  | (~\all_features[2564]  & ~\all_features[2565]  & ~new_n8907_));
  assign new_n8913_ = ~\all_features[2567]  & (~\all_features[2566]  | (~\all_features[2565]  & (new_n8900_ | ~new_n8907_ | ~\all_features[2564] )));
  assign new_n8914_ = new_n8910_ & (~\all_features[2565]  | (~\all_features[2564]  & (~\all_features[2563]  | (~\all_features[2562]  & ~\all_features[2561] ))));
  assign new_n8915_ = new_n8921_ & (~new_n8922_ | (~new_n8916_ & ~new_n8912_ & ~new_n8913_));
  assign new_n8916_ = new_n8919_ & ((~new_n8917_ & new_n8902_ & new_n8920_) | ~new_n8908_ | ~new_n8899_);
  assign new_n8917_ = \all_features[2567]  & \all_features[2566]  & ~new_n8918_ & \all_features[2565] ;
  assign new_n8918_ = ~\all_features[2563]  & ~\all_features[2564]  & (~\all_features[2562]  | new_n8900_);
  assign new_n8919_ = ~new_n8897_ & ~new_n8906_;
  assign new_n8920_ = \all_features[2566]  & \all_features[2567]  & (\all_features[2564]  | \all_features[2565]  | new_n8905_ | ~new_n8901_);
  assign new_n8921_ = ~new_n8909_ & (\all_features[2563]  | \all_features[2564]  | \all_features[2565]  | \all_features[2566]  | \all_features[2567] );
  assign new_n8922_ = ~new_n8911_ & ~new_n8914_;
  assign new_n8923_ = ~new_n8924_ & ~new_n8927_;
  assign new_n8924_ = new_n8922_ & ~new_n8925_ & new_n8921_;
  assign new_n8925_ = new_n8926_ & (~new_n8920_ | ~new_n8908_ | ~new_n8899_ | ~new_n8902_);
  assign new_n8926_ = ~new_n8906_ & ~new_n8897_ & ~new_n8912_ & ~new_n8913_;
  assign new_n8927_ = new_n8919_ & new_n8921_ & ~new_n8914_ & ~new_n8913_ & ~new_n8911_ & ~new_n8912_;
  assign new_n8928_ = ~new_n8957_ & new_n8929_;
  assign new_n8929_ = ~new_n8930_ & ~new_n8956_;
  assign new_n8930_ = new_n8943_ & (~new_n8931_ | (new_n8954_ & new_n8955_ & new_n8951_ & new_n8952_));
  assign new_n8931_ = new_n8932_ & new_n8939_;
  assign new_n8932_ = ~new_n8933_ & ~new_n8935_;
  assign new_n8933_ = ~new_n8934_ & ~\all_features[1199] ;
  assign new_n8934_ = \all_features[1197]  & \all_features[1198]  & (\all_features[1196]  | (\all_features[1194]  & \all_features[1195]  & \all_features[1193] ));
  assign new_n8935_ = ~\all_features[1199]  & (~\all_features[1198]  | ~new_n8936_ | ~new_n8937_ | ~new_n8938_);
  assign new_n8936_ = \all_features[1196]  & \all_features[1197] ;
  assign new_n8937_ = \all_features[1192]  & \all_features[1193] ;
  assign new_n8938_ = \all_features[1194]  & \all_features[1195] ;
  assign new_n8939_ = ~new_n8940_ & ~new_n8941_;
  assign new_n8940_ = ~\all_features[1199]  & (~\all_features[1198]  | (~\all_features[1196]  & ~\all_features[1197]  & ~new_n8938_));
  assign new_n8941_ = ~\all_features[1199]  & (~\all_features[1198]  | (~\all_features[1197]  & (new_n8942_ | ~new_n8938_ | ~\all_features[1196] )));
  assign new_n8942_ = ~\all_features[1192]  & ~\all_features[1193] ;
  assign new_n8943_ = new_n8944_ & new_n8948_;
  assign new_n8944_ = ~new_n8945_ & ~new_n8947_;
  assign new_n8945_ = new_n8946_ & (~\all_features[1197]  | (~\all_features[1196]  & (~\all_features[1195]  | (~\all_features[1194]  & ~\all_features[1193] ))));
  assign new_n8946_ = ~\all_features[1198]  & ~\all_features[1199] ;
  assign new_n8947_ = new_n8946_ & (~\all_features[1195]  | ~new_n8936_ | (~\all_features[1194]  & ~new_n8937_));
  assign new_n8948_ = ~new_n8949_ & ~new_n8950_;
  assign new_n8949_ = ~\all_features[1197]  & new_n8946_ & ((~\all_features[1194]  & new_n8942_) | ~\all_features[1196]  | ~\all_features[1195] );
  assign new_n8950_ = ~\all_features[1199]  & ~\all_features[1198]  & ~\all_features[1197]  & ~\all_features[1195]  & ~\all_features[1196] ;
  assign new_n8951_ = \all_features[1199]  & (\all_features[1198]  | (new_n8936_ & (\all_features[1194]  | \all_features[1195]  | \all_features[1193] )));
  assign new_n8952_ = \all_features[1198]  & \all_features[1199]  & (\all_features[1196]  | \all_features[1197]  | new_n8937_ | ~new_n8953_);
  assign new_n8953_ = ~\all_features[1194]  & ~\all_features[1195] ;
  assign new_n8954_ = \all_features[1199]  & (\all_features[1198]  | (\all_features[1197]  & (\all_features[1196]  | ~new_n8953_ | ~new_n8942_)));
  assign new_n8955_ = \all_features[1199]  & (\all_features[1197]  | \all_features[1198]  | \all_features[1196] );
  assign new_n8956_ = new_n8931_ & new_n8943_;
  assign new_n8957_ = new_n8948_ & (~new_n8944_ | (~new_n8958_ & new_n8939_));
  assign new_n8958_ = new_n8932_ & ((~new_n8959_ & new_n8952_ & new_n8951_) | ~new_n8955_ | ~new_n8954_);
  assign new_n8959_ = \all_features[1199]  & \all_features[1198]  & ~new_n8960_ & \all_features[1197] ;
  assign new_n8960_ = ~\all_features[1195]  & ~\all_features[1196]  & (~\all_features[1194]  | new_n8942_);
  assign new_n8961_ = new_n8962_ & new_n8987_;
  assign new_n8962_ = new_n8963_ & new_n8985_;
  assign new_n8963_ = new_n8982_ & ~new_n8964_ & new_n8978_;
  assign new_n8964_ = ~new_n8972_ & ~new_n8974_ & ~new_n8976_ & ~new_n8977_ & (~new_n8968_ | ~new_n8965_);
  assign new_n8965_ = \all_features[1687]  & (\all_features[1686]  | (~new_n8966_ & \all_features[1685] ));
  assign new_n8966_ = new_n8967_ & ~\all_features[1684]  & ~\all_features[1682]  & ~\all_features[1683] ;
  assign new_n8967_ = ~\all_features[1680]  & ~\all_features[1681] ;
  assign new_n8968_ = \all_features[1687]  & \all_features[1686]  & ~new_n8971_ & new_n8969_;
  assign new_n8969_ = \all_features[1687]  & (\all_features[1686]  | (new_n8970_ & (\all_features[1682]  | \all_features[1683]  | \all_features[1681] )));
  assign new_n8970_ = \all_features[1684]  & \all_features[1685] ;
  assign new_n8971_ = ~\all_features[1682]  & ~\all_features[1683]  & ~\all_features[1684]  & ~\all_features[1685]  & (~\all_features[1681]  | ~\all_features[1680] );
  assign new_n8972_ = ~\all_features[1687]  & (~\all_features[1686]  | (~\all_features[1685]  & (new_n8967_ | ~new_n8973_ | ~\all_features[1684] )));
  assign new_n8973_ = \all_features[1682]  & \all_features[1683] ;
  assign new_n8974_ = ~new_n8975_ & ~\all_features[1687] ;
  assign new_n8975_ = \all_features[1685]  & \all_features[1686]  & (\all_features[1684]  | (\all_features[1682]  & \all_features[1683]  & \all_features[1681] ));
  assign new_n8976_ = ~\all_features[1687]  & (~new_n8973_ | ~\all_features[1680]  | ~\all_features[1681]  | ~\all_features[1686]  | ~new_n8970_);
  assign new_n8977_ = ~\all_features[1687]  & (~\all_features[1686]  | (~\all_features[1684]  & ~\all_features[1685]  & ~new_n8973_));
  assign new_n8978_ = ~new_n8979_ & ~new_n8981_;
  assign new_n8979_ = ~\all_features[1685]  & new_n8980_ & ((~\all_features[1682]  & new_n8967_) | ~\all_features[1684]  | ~\all_features[1683] );
  assign new_n8980_ = ~\all_features[1686]  & ~\all_features[1687] ;
  assign new_n8981_ = ~\all_features[1687]  & ~\all_features[1686]  & ~\all_features[1685]  & ~\all_features[1683]  & ~\all_features[1684] ;
  assign new_n8982_ = ~new_n8983_ & ~new_n8984_;
  assign new_n8983_ = new_n8980_ & (~new_n8970_ | ~\all_features[1683]  | (~\all_features[1682]  & (~\all_features[1680]  | ~\all_features[1681] )));
  assign new_n8984_ = new_n8980_ & (~\all_features[1685]  | (~\all_features[1684]  & (~\all_features[1683]  | (~\all_features[1682]  & ~\all_features[1681] ))));
  assign new_n8985_ = new_n8982_ & new_n8978_ & new_n8986_ & ~new_n8974_ & ~new_n8976_;
  assign new_n8986_ = ~new_n8972_ & ~new_n8977_;
  assign new_n8987_ = new_n8978_ & (~new_n8982_ | (new_n8986_ & (new_n8988_ | new_n8974_ | new_n8976_)));
  assign new_n8988_ = new_n8965_ & (~new_n8968_ | (~new_n8989_ & \all_features[1685]  & \all_features[1686]  & \all_features[1687] ));
  assign new_n8989_ = ~\all_features[1683]  & ~\all_features[1684]  & (~\all_features[1682]  | new_n8967_);
  assign new_n8990_ = new_n8889_ & (new_n7407_ ? (new_n8855_ ? ~new_n8991_ : ~new_n8818_) : new_n9027_);
  assign new_n8991_ = ~new_n9023_ & new_n8992_ & (new_n9014_ | (~new_n9020_ & ~new_n9012_));
  assign new_n8992_ = ~new_n8993_ & ~new_n9018_;
  assign new_n8993_ = new_n9015_ & ~new_n8994_ & new_n9011_;
  assign new_n8994_ = new_n9001_ & (~new_n9009_ | ~new_n9010_ | ~new_n8998_ | ~new_n8995_);
  assign new_n8995_ = \all_features[1895]  & (\all_features[1894]  | new_n8996_);
  assign new_n8996_ = \all_features[1893]  & (\all_features[1890]  | \all_features[1891]  | \all_features[1892]  | ~new_n8997_);
  assign new_n8997_ = ~\all_features[1888]  & ~\all_features[1889] ;
  assign new_n8998_ = \all_features[1895]  & ~new_n8999_ & \all_features[1894] ;
  assign new_n8999_ = ~\all_features[1893]  & ~\all_features[1892]  & ~\all_features[1891]  & ~new_n9000_ & ~\all_features[1890] ;
  assign new_n9000_ = \all_features[1888]  & \all_features[1889] ;
  assign new_n9001_ = ~new_n9007_ & ~new_n9005_ & ~new_n9002_ & ~new_n9004_;
  assign new_n9002_ = ~\all_features[1895]  & (~\all_features[1894]  | (~\all_features[1892]  & ~\all_features[1893]  & ~new_n9003_));
  assign new_n9003_ = \all_features[1890]  & \all_features[1891] ;
  assign new_n9004_ = ~\all_features[1895]  & (~\all_features[1894]  | (~\all_features[1893]  & (new_n8997_ | ~new_n9003_ | ~\all_features[1892] )));
  assign new_n9005_ = ~new_n9006_ & ~\all_features[1895] ;
  assign new_n9006_ = \all_features[1893]  & \all_features[1894]  & (\all_features[1892]  | (\all_features[1890]  & \all_features[1891]  & \all_features[1889] ));
  assign new_n9007_ = ~\all_features[1895]  & (~\all_features[1894]  | ~new_n9000_ | ~new_n9008_ | ~new_n9003_);
  assign new_n9008_ = \all_features[1892]  & \all_features[1893] ;
  assign new_n9009_ = \all_features[1895]  & (\all_features[1894]  | (new_n9008_ & (\all_features[1890]  | \all_features[1891]  | \all_features[1889] )));
  assign new_n9010_ = \all_features[1895]  & (\all_features[1893]  | \all_features[1894]  | \all_features[1892] );
  assign new_n9011_ = ~new_n9012_ & ~new_n9014_;
  assign new_n9012_ = ~\all_features[1893]  & new_n9013_ & ((~\all_features[1890]  & new_n8997_) | ~\all_features[1892]  | ~\all_features[1891] );
  assign new_n9013_ = ~\all_features[1894]  & ~\all_features[1895] ;
  assign new_n9014_ = ~\all_features[1895]  & ~\all_features[1894]  & ~\all_features[1893]  & ~\all_features[1891]  & ~\all_features[1892] ;
  assign new_n9015_ = ~new_n9016_ & ~new_n9017_;
  assign new_n9016_ = new_n9013_ & (~\all_features[1893]  | (~\all_features[1892]  & (~\all_features[1891]  | (~\all_features[1890]  & ~\all_features[1889] ))));
  assign new_n9017_ = new_n9013_ & (~\all_features[1891]  | ~new_n9008_ | (~\all_features[1890]  & ~new_n9000_));
  assign new_n9018_ = new_n9019_ & new_n9011_ & ~new_n9016_ & ~new_n9005_;
  assign new_n9019_ = ~new_n9007_ & ~new_n9004_ & ~new_n9017_ & ~new_n9002_;
  assign new_n9020_ = ~new_n9016_ & (new_n9017_ | (~new_n9002_ & (new_n9004_ | (~new_n9021_ & ~new_n9005_))));
  assign new_n9021_ = ~new_n9007_ & (~new_n9010_ | (new_n8995_ & (~new_n9009_ | (~new_n9022_ & new_n8998_))));
  assign new_n9022_ = \all_features[1894]  & \all_features[1895]  & (\all_features[1893]  | (\all_features[1892]  & (\all_features[1891]  | \all_features[1890] )));
  assign new_n9023_ = new_n9011_ & (~new_n9015_ | (~new_n9024_ & ~new_n9002_ & ~new_n9004_));
  assign new_n9024_ = ~new_n9007_ & ~new_n9005_ & (~new_n9010_ | new_n9025_ | ~new_n8995_);
  assign new_n9025_ = ~new_n8999_ & new_n9009_ & \all_features[1894]  & \all_features[1895]  & (~\all_features[1893]  | new_n9026_);
  assign new_n9026_ = ~\all_features[1891]  & ~\all_features[1892]  & (~\all_features[1890]  | new_n8997_);
  assign new_n9027_ = new_n9055_ & new_n9057_ & new_n9045_ & (new_n9052_ | new_n9028_);
  assign new_n9028_ = ~new_n9038_ & (new_n9040_ | (~new_n9041_ & (new_n9042_ | (~new_n9029_ & ~new_n9043_))));
  assign new_n9029_ = ~new_n9036_ & (~\all_features[1023]  | new_n9030_ | (~\all_features[1020]  & ~\all_features[1021]  & ~\all_features[1022] ));
  assign new_n9030_ = \all_features[1023]  & ((~new_n9035_ & ~\all_features[1021]  & \all_features[1022] ) | (~new_n9033_ & (\all_features[1022]  | (~new_n9031_ & \all_features[1021] ))));
  assign new_n9031_ = new_n9032_ & ~\all_features[1020]  & ~\all_features[1018]  & ~\all_features[1019] ;
  assign new_n9032_ = ~\all_features[1016]  & ~\all_features[1017] ;
  assign new_n9033_ = \all_features[1023]  & (\all_features[1022]  | (new_n9034_ & (\all_features[1018]  | \all_features[1019]  | \all_features[1017] )));
  assign new_n9034_ = \all_features[1020]  & \all_features[1021] ;
  assign new_n9035_ = (~\all_features[1018]  & ~\all_features[1019]  & ~\all_features[1020]  & (~\all_features[1017]  | ~\all_features[1016] )) | (\all_features[1020]  & (\all_features[1018]  | \all_features[1019] ));
  assign new_n9036_ = ~\all_features[1023]  & (~new_n9037_ | ~\all_features[1016]  | ~\all_features[1017]  | ~\all_features[1022]  | ~new_n9034_);
  assign new_n9037_ = \all_features[1018]  & \all_features[1019] ;
  assign new_n9038_ = new_n9039_ & (~\all_features[1021]  | (~\all_features[1020]  & (~\all_features[1019]  | (~\all_features[1018]  & ~\all_features[1017] ))));
  assign new_n9039_ = ~\all_features[1022]  & ~\all_features[1023] ;
  assign new_n9040_ = new_n9039_ & (~new_n9034_ | ~\all_features[1019]  | (~\all_features[1018]  & (~\all_features[1016]  | ~\all_features[1017] )));
  assign new_n9041_ = ~\all_features[1023]  & (~\all_features[1022]  | (~\all_features[1020]  & ~\all_features[1021]  & ~new_n9037_));
  assign new_n9042_ = ~\all_features[1023]  & (~\all_features[1022]  | (~\all_features[1021]  & (new_n9032_ | ~new_n9037_ | ~\all_features[1020] )));
  assign new_n9043_ = ~new_n9044_ & ~\all_features[1023] ;
  assign new_n9044_ = \all_features[1021]  & \all_features[1022]  & (\all_features[1020]  | (\all_features[1018]  & \all_features[1019]  & \all_features[1017] ));
  assign new_n9045_ = new_n9051_ & (~new_n9053_ | (new_n9054_ & (new_n9046_ | new_n9043_ | new_n9036_)));
  assign new_n9046_ = new_n9047_ & (~new_n9048_ | (~new_n9050_ & \all_features[1021]  & \all_features[1022]  & \all_features[1023] ));
  assign new_n9047_ = \all_features[1023]  & (\all_features[1022]  | (~new_n9031_ & \all_features[1021] ));
  assign new_n9048_ = \all_features[1023]  & \all_features[1022]  & ~new_n9049_ & new_n9033_;
  assign new_n9049_ = ~\all_features[1018]  & ~\all_features[1019]  & ~\all_features[1020]  & ~\all_features[1021]  & (~\all_features[1017]  | ~\all_features[1016] );
  assign new_n9050_ = ~\all_features[1019]  & ~\all_features[1020]  & (~\all_features[1018]  | new_n9032_);
  assign new_n9051_ = ~new_n9052_ & (\all_features[1019]  | \all_features[1020]  | \all_features[1021]  | \all_features[1022]  | \all_features[1023] );
  assign new_n9052_ = ~\all_features[1021]  & new_n9039_ & ((~\all_features[1018]  & new_n9032_) | ~\all_features[1020]  | ~\all_features[1019] );
  assign new_n9053_ = ~new_n9038_ & ~new_n9040_;
  assign new_n9054_ = ~new_n9041_ & ~new_n9042_;
  assign new_n9055_ = new_n9053_ & ~new_n9056_ & new_n9051_;
  assign new_n9056_ = ~new_n9041_ & ~new_n9042_ & ~new_n9043_ & ~new_n9036_ & (~new_n9048_ | ~new_n9047_);
  assign new_n9057_ = new_n9058_ & (\all_features[1019]  | \all_features[1020]  | \all_features[1021]  | \all_features[1022]  | \all_features[1023] );
  assign new_n9058_ = new_n9053_ & new_n9051_ & new_n9054_ & ~new_n9043_ & ~new_n9036_;
  assign new_n9059_ = (new_n8928_ | new_n8889_ | (new_n8892_ ? new_n8891_ : new_n8961_)) & (~new_n9060_ | ~new_n8889_);
  assign new_n9060_ = ~new_n9027_ & ~new_n7407_;
  assign new_n9061_ = ~new_n9062_ & new_n9381_;
  assign new_n9062_ = ~new_n9169_ & ~new_n9063_ & (~new_n9277_ | new_n9278_) & (~new_n9276_ | ~new_n9345_);
  assign new_n9063_ = ~new_n9167_ & (new_n9099_ ? (new_n9133_ | ~new_n9098_) : new_n9064_);
  assign new_n9064_ = new_n9097_ & (new_n9093_ | new_n9065_);
  assign new_n9065_ = ~new_n9066_ & (\all_features[1763]  | \all_features[1764]  | \all_features[1765]  | \all_features[1766]  | \all_features[1767] );
  assign new_n9066_ = new_n9067_ & (new_n9090_ | (~new_n9088_ & (new_n9081_ | (~new_n9091_ & ~new_n9083_))));
  assign new_n9067_ = ~new_n9085_ & ~new_n9089_ & ~new_n9087_ & (new_n9090_ | new_n9088_ | new_n9068_);
  assign new_n9068_ = ~new_n9081_ & ~new_n9083_ & (~new_n9075_ | (~new_n9079_ & new_n9069_));
  assign new_n9069_ = \all_features[1767]  & \all_features[1766]  & ~new_n9070_ & new_n9073_;
  assign new_n9070_ = new_n9072_ & ~\all_features[1765]  & ~new_n9071_ & ~\all_features[1764] ;
  assign new_n9071_ = \all_features[1760]  & \all_features[1761] ;
  assign new_n9072_ = ~\all_features[1762]  & ~\all_features[1763] ;
  assign new_n9073_ = \all_features[1767]  & (\all_features[1766]  | (new_n9074_ & (\all_features[1762]  | \all_features[1763]  | \all_features[1761] )));
  assign new_n9074_ = \all_features[1764]  & \all_features[1765] ;
  assign new_n9075_ = new_n9076_ & new_n9078_;
  assign new_n9076_ = \all_features[1767]  & (\all_features[1766]  | (\all_features[1765]  & (\all_features[1764]  | ~new_n9072_ | ~new_n9077_)));
  assign new_n9077_ = ~\all_features[1760]  & ~\all_features[1761] ;
  assign new_n9078_ = \all_features[1767]  & (\all_features[1765]  | \all_features[1766]  | \all_features[1764] );
  assign new_n9079_ = \all_features[1767]  & \all_features[1766]  & ~new_n9080_ & \all_features[1765] ;
  assign new_n9080_ = ~\all_features[1763]  & ~\all_features[1764]  & (~\all_features[1762]  | new_n9077_);
  assign new_n9081_ = ~new_n9082_ & ~\all_features[1767] ;
  assign new_n9082_ = \all_features[1765]  & \all_features[1766]  & (\all_features[1764]  | (\all_features[1762]  & \all_features[1763]  & \all_features[1761] ));
  assign new_n9083_ = ~\all_features[1767]  & (~\all_features[1766]  | ~new_n9084_ | ~new_n9071_ | ~new_n9074_);
  assign new_n9084_ = \all_features[1762]  & \all_features[1763] ;
  assign new_n9085_ = new_n9086_ & (~\all_features[1765]  | (~\all_features[1764]  & (~\all_features[1763]  | (~\all_features[1762]  & ~\all_features[1761] ))));
  assign new_n9086_ = ~\all_features[1766]  & ~\all_features[1767] ;
  assign new_n9087_ = ~\all_features[1765]  & new_n9086_ & ((~\all_features[1762]  & new_n9077_) | ~\all_features[1764]  | ~\all_features[1763] );
  assign new_n9088_ = ~\all_features[1767]  & (~\all_features[1766]  | (~\all_features[1765]  & (new_n9077_ | ~new_n9084_ | ~\all_features[1764] )));
  assign new_n9089_ = new_n9086_ & (~\all_features[1763]  | ~new_n9074_ | (~\all_features[1762]  & ~new_n9071_));
  assign new_n9090_ = ~\all_features[1767]  & (~\all_features[1766]  | (~\all_features[1764]  & ~\all_features[1765]  & ~new_n9084_));
  assign new_n9091_ = new_n9078_ & (~new_n9076_ | (~new_n9092_ & new_n9073_));
  assign new_n9092_ = ~\all_features[1765]  & \all_features[1766]  & \all_features[1767]  & (\all_features[1764]  ? new_n9072_ : (new_n9071_ | ~new_n9072_));
  assign new_n9093_ = new_n9096_ & ~new_n9089_ & ~new_n9094_ & ~new_n9085_;
  assign new_n9094_ = ~new_n9081_ & ~new_n9088_ & new_n9095_ & (~new_n9075_ | ~new_n9069_);
  assign new_n9095_ = ~new_n9083_ & ~new_n9090_;
  assign new_n9096_ = ~new_n9087_ & (\all_features[1763]  | \all_features[1764]  | \all_features[1765]  | \all_features[1766]  | \all_features[1767] );
  assign new_n9097_ = new_n9095_ & new_n9096_ & ~new_n9089_ & ~new_n9088_ & ~new_n9081_ & ~new_n9085_;
  assign new_n9098_ = ~new_n6734_ & (~new_n6732_ | new_n6702_);
  assign new_n9099_ = ~new_n9129_ & (~new_n9131_ | ~new_n9100_);
  assign new_n9100_ = new_n9101_ & new_n9122_;
  assign new_n9101_ = ~new_n9102_ & (\all_features[3267]  | \all_features[3268]  | \all_features[3269]  | \all_features[3270]  | \all_features[3271] );
  assign new_n9102_ = ~new_n9118_ & (new_n9116_ | (~new_n9120_ & (new_n9121_ | (~new_n9119_ & ~new_n9103_))));
  assign new_n9103_ = ~new_n9104_ & (new_n9106_ | (new_n9115_ & (~new_n9110_ | (~new_n9114_ & new_n9113_))));
  assign new_n9104_ = ~new_n9105_ & ~\all_features[3271] ;
  assign new_n9105_ = \all_features[3269]  & \all_features[3270]  & (\all_features[3268]  | (\all_features[3266]  & \all_features[3267]  & \all_features[3265] ));
  assign new_n9106_ = ~\all_features[3271]  & (~\all_features[3270]  | ~new_n9107_ | ~new_n9108_ | ~new_n9109_);
  assign new_n9107_ = \all_features[3266]  & \all_features[3267] ;
  assign new_n9108_ = \all_features[3264]  & \all_features[3265] ;
  assign new_n9109_ = \all_features[3268]  & \all_features[3269] ;
  assign new_n9110_ = \all_features[3271]  & (\all_features[3270]  | (\all_features[3269]  & (\all_features[3268]  | ~new_n9112_ | ~new_n9111_)));
  assign new_n9111_ = ~\all_features[3264]  & ~\all_features[3265] ;
  assign new_n9112_ = ~\all_features[3266]  & ~\all_features[3267] ;
  assign new_n9113_ = \all_features[3271]  & (\all_features[3270]  | (new_n9109_ & (\all_features[3266]  | \all_features[3267]  | \all_features[3265] )));
  assign new_n9114_ = ~\all_features[3269]  & \all_features[3270]  & \all_features[3271]  & (\all_features[3268]  ? new_n9112_ : (new_n9108_ | ~new_n9112_));
  assign new_n9115_ = \all_features[3271]  & (\all_features[3269]  | \all_features[3270]  | \all_features[3268] );
  assign new_n9116_ = new_n9117_ & (~\all_features[3269]  | (~\all_features[3268]  & (~\all_features[3267]  | (~\all_features[3266]  & ~\all_features[3265] ))));
  assign new_n9117_ = ~\all_features[3270]  & ~\all_features[3271] ;
  assign new_n9118_ = ~\all_features[3269]  & new_n9117_ & ((~\all_features[3266]  & new_n9111_) | ~\all_features[3268]  | ~\all_features[3267] );
  assign new_n9119_ = ~\all_features[3271]  & (~\all_features[3270]  | (~\all_features[3269]  & (new_n9111_ | ~new_n9107_ | ~\all_features[3268] )));
  assign new_n9120_ = new_n9117_ & (~\all_features[3267]  | ~new_n9109_ | (~\all_features[3266]  & ~new_n9108_));
  assign new_n9121_ = ~\all_features[3271]  & (~\all_features[3270]  | (~\all_features[3268]  & ~\all_features[3269]  & ~new_n9107_));
  assign new_n9122_ = new_n9127_ & (~new_n9128_ | (~new_n9123_ & ~new_n9119_ & ~new_n9121_));
  assign new_n9123_ = ~new_n9104_ & ~new_n9106_ & (~new_n9115_ | ~new_n9110_ | new_n9124_);
  assign new_n9124_ = new_n9113_ & new_n9125_ & (new_n9126_ | ~\all_features[3269]  | ~\all_features[3270]  | ~\all_features[3271] );
  assign new_n9125_ = \all_features[3270]  & \all_features[3271]  & (\all_features[3268]  | \all_features[3269]  | new_n9108_ | ~new_n9112_);
  assign new_n9126_ = ~\all_features[3267]  & ~\all_features[3268]  & (~\all_features[3266]  | new_n9111_);
  assign new_n9127_ = ~new_n9118_ & (\all_features[3267]  | \all_features[3268]  | \all_features[3269]  | \all_features[3270]  | \all_features[3271] );
  assign new_n9128_ = ~new_n9116_ & ~new_n9120_;
  assign new_n9129_ = new_n9130_ & new_n9127_ & ~new_n9120_ & ~new_n9119_ & ~new_n9104_ & ~new_n9116_;
  assign new_n9130_ = ~new_n9106_ & ~new_n9121_;
  assign new_n9131_ = new_n9127_ & new_n9128_ & (new_n9132_ | new_n9104_ | new_n9119_ | ~new_n9130_);
  assign new_n9132_ = new_n9115_ & new_n9125_ & new_n9110_ & new_n9113_;
  assign new_n9133_ = ~new_n9163_ & (~new_n9165_ | new_n9134_);
  assign new_n9134_ = ~new_n9135_ & ~new_n9159_;
  assign new_n9135_ = new_n9151_ & (~new_n9154_ | (~new_n9136_ & ~new_n9157_ & ~new_n9158_));
  assign new_n9136_ = ~new_n9145_ & ~new_n9147_ & (~new_n9150_ | ~new_n9149_ | new_n9137_);
  assign new_n9137_ = new_n9138_ & new_n9140_ & (new_n9143_ | ~\all_features[1989]  | ~\all_features[1990]  | ~\all_features[1991] );
  assign new_n9138_ = \all_features[1991]  & (\all_features[1990]  | (new_n9139_ & (\all_features[1986]  | \all_features[1987]  | \all_features[1985] )));
  assign new_n9139_ = \all_features[1988]  & \all_features[1989] ;
  assign new_n9140_ = \all_features[1990]  & \all_features[1991]  & (\all_features[1988]  | \all_features[1989]  | new_n9141_ | ~new_n9142_);
  assign new_n9141_ = \all_features[1984]  & \all_features[1985] ;
  assign new_n9142_ = ~\all_features[1986]  & ~\all_features[1987] ;
  assign new_n9143_ = ~\all_features[1987]  & ~\all_features[1988]  & (~\all_features[1986]  | new_n9144_);
  assign new_n9144_ = ~\all_features[1984]  & ~\all_features[1985] ;
  assign new_n9145_ = ~new_n9146_ & ~\all_features[1991] ;
  assign new_n9146_ = \all_features[1989]  & \all_features[1990]  & (\all_features[1988]  | (\all_features[1986]  & \all_features[1987]  & \all_features[1985] ));
  assign new_n9147_ = ~\all_features[1991]  & (~\all_features[1990]  | ~new_n9148_ | ~new_n9141_ | ~new_n9139_);
  assign new_n9148_ = \all_features[1986]  & \all_features[1987] ;
  assign new_n9149_ = \all_features[1991]  & (\all_features[1990]  | (\all_features[1989]  & (\all_features[1988]  | ~new_n9142_ | ~new_n9144_)));
  assign new_n9150_ = \all_features[1991]  & (\all_features[1989]  | \all_features[1990]  | \all_features[1988] );
  assign new_n9151_ = ~new_n9152_ & (\all_features[1987]  | \all_features[1988]  | \all_features[1989]  | \all_features[1990]  | \all_features[1991] );
  assign new_n9152_ = ~\all_features[1989]  & new_n9153_ & ((~\all_features[1986]  & new_n9144_) | ~\all_features[1988]  | ~\all_features[1987] );
  assign new_n9153_ = ~\all_features[1990]  & ~\all_features[1991] ;
  assign new_n9154_ = ~new_n9155_ & ~new_n9156_;
  assign new_n9155_ = new_n9153_ & (~\all_features[1989]  | (~\all_features[1988]  & (~\all_features[1987]  | (~\all_features[1986]  & ~\all_features[1985] ))));
  assign new_n9156_ = new_n9153_ & (~\all_features[1987]  | ~new_n9139_ | (~\all_features[1986]  & ~new_n9141_));
  assign new_n9157_ = ~\all_features[1991]  & (~\all_features[1990]  | (~\all_features[1989]  & (new_n9144_ | ~new_n9148_ | ~\all_features[1988] )));
  assign new_n9158_ = ~\all_features[1991]  & (~\all_features[1990]  | (~\all_features[1988]  & ~\all_features[1989]  & ~new_n9148_));
  assign new_n9159_ = ~new_n9160_ & (\all_features[1987]  | \all_features[1988]  | \all_features[1989]  | \all_features[1990]  | \all_features[1991] );
  assign new_n9160_ = ~new_n9152_ & (new_n9155_ | (~new_n9156_ & (new_n9158_ | (~new_n9157_ & ~new_n9161_))));
  assign new_n9161_ = ~new_n9145_ & (new_n9147_ | (new_n9150_ & (~new_n9149_ | (~new_n9162_ & new_n9138_))));
  assign new_n9162_ = ~\all_features[1989]  & \all_features[1990]  & \all_features[1991]  & (\all_features[1988]  ? new_n9142_ : (new_n9141_ | ~new_n9142_));
  assign new_n9163_ = new_n9164_ & new_n9151_ & ~new_n9156_ & ~new_n9157_ & ~new_n9145_ & ~new_n9155_;
  assign new_n9164_ = ~new_n9147_ & ~new_n9158_;
  assign new_n9165_ = new_n9151_ & new_n9154_ & (new_n9166_ | new_n9145_ | new_n9157_ | ~new_n9164_);
  assign new_n9166_ = new_n9150_ & new_n9140_ & new_n9149_ & new_n9138_;
  assign new_n9167_ = new_n9168_ & new_n7902_;
  assign new_n9168_ = new_n7899_ & new_n7870_;
  assign new_n9169_ = new_n9208_ & (new_n9170_ ? ~new_n9247_ : new_n9245_);
  assign new_n9170_ = ~new_n9171_ & new_n9203_;
  assign new_n9171_ = ~new_n9172_ & ~new_n9193_;
  assign new_n9172_ = ~new_n9173_ & (\all_features[3547]  | \all_features[3548]  | \all_features[3549]  | \all_features[3550]  | \all_features[3551] );
  assign new_n9173_ = ~new_n9187_ & (new_n9189_ | (~new_n9190_ & (new_n9191_ | (~new_n9174_ & ~new_n9192_))));
  assign new_n9174_ = ~new_n9182_ & (new_n9184_ | (~new_n9175_ & new_n9186_));
  assign new_n9175_ = \all_features[3551]  & ((~new_n9180_ & ~\all_features[3549]  & \all_features[3550] ) | (~new_n9178_ & (\all_features[3550]  | (~new_n9176_ & \all_features[3549] ))));
  assign new_n9176_ = new_n9177_ & ~\all_features[3548]  & ~\all_features[3546]  & ~\all_features[3547] ;
  assign new_n9177_ = ~\all_features[3544]  & ~\all_features[3545] ;
  assign new_n9178_ = \all_features[3551]  & (\all_features[3550]  | (new_n9179_ & (\all_features[3546]  | \all_features[3547]  | \all_features[3545] )));
  assign new_n9179_ = \all_features[3548]  & \all_features[3549] ;
  assign new_n9180_ = (\all_features[3548]  & (\all_features[3546]  | \all_features[3547] )) | (~new_n9181_ & ~\all_features[3546]  & ~\all_features[3547]  & ~\all_features[3548] );
  assign new_n9181_ = \all_features[3544]  & \all_features[3545] ;
  assign new_n9182_ = ~new_n9183_ & ~\all_features[3551] ;
  assign new_n9183_ = \all_features[3549]  & \all_features[3550]  & (\all_features[3548]  | (\all_features[3546]  & \all_features[3547]  & \all_features[3545] ));
  assign new_n9184_ = ~\all_features[3551]  & (~\all_features[3550]  | ~new_n9181_ | ~new_n9179_ | ~new_n9185_);
  assign new_n9185_ = \all_features[3546]  & \all_features[3547] ;
  assign new_n9186_ = \all_features[3551]  & (\all_features[3549]  | \all_features[3550]  | \all_features[3548] );
  assign new_n9187_ = ~\all_features[3549]  & new_n9188_ & ((~\all_features[3546]  & new_n9177_) | ~\all_features[3548]  | ~\all_features[3547] );
  assign new_n9188_ = ~\all_features[3550]  & ~\all_features[3551] ;
  assign new_n9189_ = new_n9188_ & (~\all_features[3549]  | (~\all_features[3548]  & (~\all_features[3547]  | (~\all_features[3546]  & ~\all_features[3545] ))));
  assign new_n9190_ = new_n9188_ & (~\all_features[3547]  | ~new_n9179_ | (~\all_features[3546]  & ~new_n9181_));
  assign new_n9191_ = ~\all_features[3551]  & (~\all_features[3550]  | (~\all_features[3548]  & ~\all_features[3549]  & ~new_n9185_));
  assign new_n9192_ = ~\all_features[3551]  & (~\all_features[3550]  | (~\all_features[3549]  & (new_n9177_ | ~new_n9185_ | ~\all_features[3548] )));
  assign new_n9193_ = new_n9199_ & (~new_n9200_ | (new_n9201_ & (~new_n9202_ | new_n9194_)));
  assign new_n9194_ = new_n9195_ & (~new_n9196_ | (~new_n9198_ & \all_features[3549]  & \all_features[3550]  & \all_features[3551] ));
  assign new_n9195_ = \all_features[3551]  & (\all_features[3550]  | (~new_n9176_ & \all_features[3549] ));
  assign new_n9196_ = \all_features[3551]  & \all_features[3550]  & ~new_n9197_ & new_n9178_;
  assign new_n9197_ = ~\all_features[3549]  & ~\all_features[3548]  & ~\all_features[3547]  & ~new_n9181_ & ~\all_features[3546] ;
  assign new_n9198_ = ~\all_features[3547]  & ~\all_features[3548]  & (~\all_features[3546]  | new_n9177_);
  assign new_n9199_ = ~new_n9187_ & (\all_features[3547]  | \all_features[3548]  | \all_features[3549]  | \all_features[3550]  | \all_features[3551] );
  assign new_n9200_ = ~new_n9189_ & ~new_n9190_;
  assign new_n9201_ = ~new_n9191_ & ~new_n9192_;
  assign new_n9202_ = ~new_n9182_ & ~new_n9184_;
  assign new_n9203_ = new_n9204_ & new_n9207_;
  assign new_n9204_ = new_n9205_ & (new_n9192_ | new_n9182_ | ~new_n9206_ | (new_n9196_ & new_n9195_));
  assign new_n9205_ = new_n9199_ & new_n9200_;
  assign new_n9206_ = ~new_n9191_ & ~new_n9184_;
  assign new_n9207_ = new_n9202_ & new_n9205_ & new_n9201_;
  assign new_n9208_ = ~new_n9209_ & new_n9167_;
  assign new_n9209_ = new_n9210_ & new_n9236_;
  assign new_n9210_ = ~new_n9211_ & ~new_n9234_;
  assign new_n9211_ = new_n9229_ & ~new_n9233_ & ~new_n9212_ & ~new_n9232_;
  assign new_n9212_ = ~new_n9227_ & ~new_n9228_ & new_n9220_ & (~new_n9225_ | ~new_n9213_);
  assign new_n9213_ = new_n9219_ & new_n9214_ & new_n9216_;
  assign new_n9214_ = \all_features[1871]  & (\all_features[1870]  | (new_n9215_ & (\all_features[1866]  | \all_features[1867]  | \all_features[1865] )));
  assign new_n9215_ = \all_features[1868]  & \all_features[1869] ;
  assign new_n9216_ = \all_features[1870]  & \all_features[1871]  & (\all_features[1868]  | \all_features[1869]  | new_n9218_ | ~new_n9217_);
  assign new_n9217_ = ~\all_features[1866]  & ~\all_features[1867] ;
  assign new_n9218_ = \all_features[1864]  & \all_features[1865] ;
  assign new_n9219_ = \all_features[1871]  & (\all_features[1869]  | \all_features[1870]  | \all_features[1868] );
  assign new_n9220_ = ~new_n9221_ & ~new_n9223_;
  assign new_n9221_ = ~new_n9222_ & ~\all_features[1871] ;
  assign new_n9222_ = \all_features[1869]  & \all_features[1870]  & (\all_features[1868]  | (\all_features[1866]  & \all_features[1867]  & \all_features[1865] ));
  assign new_n9223_ = ~\all_features[1871]  & (~\all_features[1870]  | (~\all_features[1868]  & ~\all_features[1869]  & ~new_n9224_));
  assign new_n9224_ = \all_features[1866]  & \all_features[1867] ;
  assign new_n9225_ = \all_features[1871]  & (\all_features[1870]  | (\all_features[1869]  & (\all_features[1868]  | ~new_n9226_ | ~new_n9217_)));
  assign new_n9226_ = ~\all_features[1864]  & ~\all_features[1865] ;
  assign new_n9227_ = ~\all_features[1871]  & (~\all_features[1870]  | (~\all_features[1869]  & (new_n9226_ | ~new_n9224_ | ~\all_features[1868] )));
  assign new_n9228_ = ~\all_features[1871]  & (~\all_features[1870]  | ~new_n9215_ | ~new_n9218_ | ~new_n9224_);
  assign new_n9229_ = ~new_n9230_ & (\all_features[1867]  | \all_features[1868]  | \all_features[1869]  | \all_features[1870]  | \all_features[1871] );
  assign new_n9230_ = ~\all_features[1869]  & new_n9231_ & ((~\all_features[1866]  & new_n9226_) | ~\all_features[1868]  | ~\all_features[1867] );
  assign new_n9231_ = ~\all_features[1870]  & ~\all_features[1871] ;
  assign new_n9232_ = new_n9231_ & (~\all_features[1869]  | (~\all_features[1868]  & (~\all_features[1867]  | (~\all_features[1866]  & ~\all_features[1865] ))));
  assign new_n9233_ = new_n9231_ & (~\all_features[1867]  | ~new_n9215_ | (~\all_features[1866]  & ~new_n9218_));
  assign new_n9234_ = new_n9229_ & new_n9220_ & new_n9235_ & ~new_n9227_ & ~new_n9228_;
  assign new_n9235_ = ~new_n9232_ & ~new_n9233_;
  assign new_n9236_ = ~new_n9237_ & ~new_n9241_;
  assign new_n9237_ = ~new_n9238_ & (\all_features[1867]  | \all_features[1868]  | \all_features[1869]  | \all_features[1870]  | \all_features[1871] );
  assign new_n9238_ = ~new_n9230_ & (new_n9232_ | (~new_n9233_ & (new_n9223_ | (~new_n9227_ & ~new_n9239_))));
  assign new_n9239_ = ~new_n9221_ & (new_n9228_ | (new_n9219_ & (~new_n9225_ | (~new_n9240_ & new_n9214_))));
  assign new_n9240_ = ~\all_features[1869]  & \all_features[1870]  & \all_features[1871]  & (\all_features[1868]  ? new_n9217_ : (new_n9218_ | ~new_n9217_));
  assign new_n9241_ = new_n9229_ & (~new_n9235_ | (~new_n9242_ & ~new_n9223_ & ~new_n9227_));
  assign new_n9242_ = ~new_n9228_ & ~new_n9221_ & (~new_n9219_ | ~new_n9225_ | new_n9243_);
  assign new_n9243_ = new_n9214_ & new_n9216_ & (new_n9244_ | ~\all_features[1869]  | ~\all_features[1870]  | ~\all_features[1871] );
  assign new_n9244_ = ~\all_features[1867]  & ~\all_features[1868]  & (~\all_features[1866]  | new_n9226_);
  assign new_n9245_ = ~new_n8777_ & new_n9246_;
  assign new_n9246_ = new_n8807_ & new_n8810_;
  assign new_n9247_ = ~new_n9248_ & new_n9275_;
  assign new_n9248_ = ~new_n9249_ & ~new_n9271_;
  assign new_n9249_ = new_n9250_ & (~new_n9259_ | (new_n9269_ & new_n9270_ & new_n9266_ & new_n9268_));
  assign new_n9250_ = new_n9251_ & ~new_n9255_ & ~new_n9256_;
  assign new_n9251_ = ~new_n9252_ & (\all_features[3003]  | \all_features[3004]  | \all_features[3005]  | \all_features[3006]  | \all_features[3007] );
  assign new_n9252_ = ~\all_features[3005]  & new_n9254_ & ((~\all_features[3002]  & new_n9253_) | ~\all_features[3004]  | ~\all_features[3003] );
  assign new_n9253_ = ~\all_features[3000]  & ~\all_features[3001] ;
  assign new_n9254_ = ~\all_features[3006]  & ~\all_features[3007] ;
  assign new_n9255_ = new_n9254_ & (~\all_features[3005]  | (~\all_features[3004]  & (~\all_features[3003]  | (~\all_features[3002]  & ~\all_features[3001] ))));
  assign new_n9256_ = new_n9254_ & (~\all_features[3003]  | ~new_n9257_ | (~\all_features[3002]  & ~new_n9258_));
  assign new_n9257_ = \all_features[3004]  & \all_features[3005] ;
  assign new_n9258_ = \all_features[3000]  & \all_features[3001] ;
  assign new_n9259_ = ~new_n9265_ & ~new_n9264_ & ~new_n9260_ & ~new_n9262_;
  assign new_n9260_ = ~\all_features[3007]  & (~\all_features[3006]  | (~\all_features[3005]  & (new_n9253_ | ~new_n9261_ | ~\all_features[3004] )));
  assign new_n9261_ = \all_features[3002]  & \all_features[3003] ;
  assign new_n9262_ = ~new_n9263_ & ~\all_features[3007] ;
  assign new_n9263_ = \all_features[3005]  & \all_features[3006]  & (\all_features[3004]  | (\all_features[3002]  & \all_features[3003]  & \all_features[3001] ));
  assign new_n9264_ = ~\all_features[3007]  & (~\all_features[3006]  | ~new_n9257_ | ~new_n9258_ | ~new_n9261_);
  assign new_n9265_ = ~\all_features[3007]  & (~\all_features[3006]  | (~\all_features[3004]  & ~\all_features[3005]  & ~new_n9261_));
  assign new_n9266_ = \all_features[3007]  & (\all_features[3006]  | (\all_features[3005]  & (\all_features[3004]  | ~new_n9253_ | ~new_n9267_)));
  assign new_n9267_ = ~\all_features[3002]  & ~\all_features[3003] ;
  assign new_n9268_ = \all_features[3007]  & (\all_features[3006]  | (new_n9257_ & (\all_features[3002]  | \all_features[3003]  | \all_features[3001] )));
  assign new_n9269_ = \all_features[3006]  & \all_features[3007]  & (\all_features[3004]  | \all_features[3005]  | new_n9258_ | ~new_n9267_);
  assign new_n9270_ = \all_features[3007]  & (\all_features[3005]  | \all_features[3006]  | \all_features[3004] );
  assign new_n9271_ = new_n9251_ & (new_n9256_ | new_n9255_ | (~new_n9260_ & ~new_n9265_ & ~new_n9272_));
  assign new_n9272_ = ~new_n9264_ & ~new_n9262_ & (~new_n9270_ | ~new_n9266_ | new_n9273_);
  assign new_n9273_ = new_n9268_ & new_n9269_ & (new_n9274_ | ~\all_features[3005]  | ~\all_features[3006]  | ~\all_features[3007] );
  assign new_n9274_ = ~\all_features[3003]  & ~\all_features[3004]  & (~\all_features[3002]  | new_n9253_);
  assign new_n9275_ = new_n9250_ & new_n9259_;
  assign new_n9276_ = ~new_n9167_ & ~new_n9064_ & ~new_n9099_;
  assign new_n9277_ = new_n9167_ & new_n9209_;
  assign new_n9278_ = ~new_n9279_ & new_n9312_;
  assign new_n9279_ = ~new_n9280_ & new_n9308_;
  assign new_n9280_ = ~new_n9307_ & (new_n9300_ | new_n9303_ | new_n9305_ | new_n9306_ | new_n9281_);
  assign new_n9281_ = ~new_n9294_ & ~new_n9299_ & ((~new_n9282_ & new_n9291_) | new_n9298_ | new_n9296_);
  assign new_n9282_ = new_n9283_ & (new_n9289_ | ~\all_features[813]  | ~\all_features[814]  | ~\all_features[815] );
  assign new_n9283_ = \all_features[815]  & \all_features[814]  & ~new_n9284_ & new_n9287_;
  assign new_n9284_ = new_n9285_ & ~\all_features[813]  & ~new_n9286_ & ~\all_features[812] ;
  assign new_n9285_ = ~\all_features[810]  & ~\all_features[811] ;
  assign new_n9286_ = \all_features[808]  & \all_features[809] ;
  assign new_n9287_ = \all_features[815]  & (\all_features[814]  | (new_n9288_ & (\all_features[810]  | \all_features[811]  | \all_features[809] )));
  assign new_n9288_ = \all_features[812]  & \all_features[813] ;
  assign new_n9289_ = ~\all_features[811]  & ~\all_features[812]  & (~\all_features[810]  | new_n9290_);
  assign new_n9290_ = ~\all_features[808]  & ~\all_features[809] ;
  assign new_n9291_ = new_n9292_ & new_n9293_;
  assign new_n9292_ = \all_features[815]  & (\all_features[814]  | (\all_features[813]  & (\all_features[812]  | ~new_n9290_ | ~new_n9285_)));
  assign new_n9293_ = \all_features[815]  & (\all_features[813]  | \all_features[814]  | \all_features[812] );
  assign new_n9294_ = ~\all_features[815]  & (~\all_features[814]  | (~\all_features[813]  & (new_n9290_ | ~new_n9295_ | ~\all_features[812] )));
  assign new_n9295_ = \all_features[810]  & \all_features[811] ;
  assign new_n9296_ = ~new_n9297_ & ~\all_features[815] ;
  assign new_n9297_ = \all_features[813]  & \all_features[814]  & (\all_features[812]  | (\all_features[810]  & \all_features[811]  & \all_features[809] ));
  assign new_n9298_ = ~\all_features[815]  & (~\all_features[814]  | ~new_n9286_ | ~new_n9288_ | ~new_n9295_);
  assign new_n9299_ = ~\all_features[815]  & (~\all_features[814]  | (~\all_features[812]  & ~\all_features[813]  & ~new_n9295_));
  assign new_n9300_ = ~new_n9299_ & (new_n9294_ | (~new_n9296_ & (new_n9298_ | new_n9301_)));
  assign new_n9301_ = new_n9293_ & (~new_n9292_ | (~new_n9302_ & new_n9287_));
  assign new_n9302_ = ~\all_features[813]  & \all_features[814]  & \all_features[815]  & (\all_features[812]  ? new_n9285_ : (new_n9286_ | ~new_n9285_));
  assign new_n9303_ = new_n9304_ & (~\all_features[813]  | (~\all_features[812]  & (~\all_features[811]  | (~\all_features[810]  & ~\all_features[809] ))));
  assign new_n9304_ = ~\all_features[814]  & ~\all_features[815] ;
  assign new_n9305_ = new_n9304_ & (~\all_features[811]  | ~new_n9288_ | (~\all_features[810]  & ~new_n9286_));
  assign new_n9306_ = ~\all_features[813]  & new_n9304_ & ((~\all_features[810]  & new_n9290_) | ~\all_features[812]  | ~\all_features[811] );
  assign new_n9307_ = ~\all_features[815]  & ~\all_features[814]  & ~\all_features[813]  & ~\all_features[811]  & ~\all_features[812] ;
  assign new_n9308_ = new_n9303_ | ~new_n9310_ | ((new_n9296_ | ~new_n9311_) & (new_n9309_ | new_n9305_));
  assign new_n9309_ = ~new_n9294_ & ~new_n9296_ & ~new_n9298_ & ~new_n9299_ & (~new_n9291_ | ~new_n9283_);
  assign new_n9310_ = ~new_n9306_ & ~new_n9307_;
  assign new_n9311_ = ~new_n9305_ & ~new_n9299_ & ~new_n9294_ & ~new_n9298_;
  assign new_n9312_ = ~new_n9341_ & new_n9313_;
  assign new_n9313_ = ~new_n9314_ & ~new_n9340_;
  assign new_n9314_ = new_n9327_ & (~new_n9315_ | (new_n9338_ & new_n9339_ & new_n9335_ & new_n9336_));
  assign new_n9315_ = new_n9316_ & new_n9323_;
  assign new_n9316_ = ~new_n9317_ & ~new_n9319_;
  assign new_n9317_ = ~new_n9318_ & ~\all_features[2175] ;
  assign new_n9318_ = \all_features[2173]  & \all_features[2174]  & (\all_features[2172]  | (\all_features[2170]  & \all_features[2171]  & \all_features[2169] ));
  assign new_n9319_ = ~\all_features[2175]  & (~\all_features[2174]  | ~new_n9320_ | ~new_n9321_ | ~new_n9322_);
  assign new_n9320_ = \all_features[2172]  & \all_features[2173] ;
  assign new_n9321_ = \all_features[2168]  & \all_features[2169] ;
  assign new_n9322_ = \all_features[2170]  & \all_features[2171] ;
  assign new_n9323_ = ~new_n9324_ & ~new_n9325_;
  assign new_n9324_ = ~\all_features[2175]  & (~\all_features[2174]  | (~\all_features[2172]  & ~\all_features[2173]  & ~new_n9322_));
  assign new_n9325_ = ~\all_features[2175]  & (~\all_features[2174]  | (~\all_features[2173]  & (new_n9326_ | ~new_n9322_ | ~\all_features[2172] )));
  assign new_n9326_ = ~\all_features[2168]  & ~\all_features[2169] ;
  assign new_n9327_ = new_n9328_ & new_n9332_;
  assign new_n9328_ = ~new_n9329_ & ~new_n9331_;
  assign new_n9329_ = new_n9330_ & (~\all_features[2173]  | (~\all_features[2172]  & (~\all_features[2171]  | (~\all_features[2170]  & ~\all_features[2169] ))));
  assign new_n9330_ = ~\all_features[2174]  & ~\all_features[2175] ;
  assign new_n9331_ = new_n9330_ & (~\all_features[2171]  | ~new_n9320_ | (~\all_features[2170]  & ~new_n9321_));
  assign new_n9332_ = ~new_n9333_ & ~new_n9334_;
  assign new_n9333_ = ~\all_features[2173]  & new_n9330_ & ((~\all_features[2170]  & new_n9326_) | ~\all_features[2172]  | ~\all_features[2171] );
  assign new_n9334_ = ~\all_features[2175]  & ~\all_features[2174]  & ~\all_features[2173]  & ~\all_features[2171]  & ~\all_features[2172] ;
  assign new_n9335_ = \all_features[2175]  & (\all_features[2174]  | (new_n9320_ & (\all_features[2170]  | \all_features[2171]  | \all_features[2169] )));
  assign new_n9336_ = \all_features[2174]  & \all_features[2175]  & (\all_features[2172]  | \all_features[2173]  | new_n9321_ | ~new_n9337_);
  assign new_n9337_ = ~\all_features[2170]  & ~\all_features[2171] ;
  assign new_n9338_ = \all_features[2175]  & (\all_features[2174]  | (\all_features[2173]  & (\all_features[2172]  | ~new_n9337_ | ~new_n9326_)));
  assign new_n9339_ = \all_features[2175]  & (\all_features[2173]  | \all_features[2174]  | \all_features[2172] );
  assign new_n9340_ = new_n9315_ & new_n9327_;
  assign new_n9341_ = new_n9332_ & (~new_n9328_ | (~new_n9342_ & new_n9323_));
  assign new_n9342_ = new_n9316_ & ((~new_n9343_ & new_n9336_ & new_n9335_) | ~new_n9339_ | ~new_n9338_);
  assign new_n9343_ = \all_features[2175]  & \all_features[2174]  & ~new_n9344_ & \all_features[2173] ;
  assign new_n9344_ = ~\all_features[2171]  & ~\all_features[2172]  & (~\all_features[2170]  | new_n9326_);
  assign new_n9345_ = ~new_n9346_ & new_n9375_;
  assign new_n9346_ = ~new_n9347_ & ~new_n9371_;
  assign new_n9347_ = new_n9362_ & (~new_n9367_ | (~new_n9365_ & ~new_n9348_ & ~new_n9370_));
  assign new_n9348_ = ~new_n9360_ & ~new_n9358_ & (~new_n9361_ | ~new_n9357_ | new_n9349_);
  assign new_n9349_ = new_n9350_ & new_n9352_ & (new_n9355_ | ~\all_features[1245]  | ~\all_features[1246]  | ~\all_features[1247] );
  assign new_n9350_ = \all_features[1247]  & (\all_features[1246]  | (new_n9351_ & (\all_features[1242]  | \all_features[1243]  | \all_features[1241] )));
  assign new_n9351_ = \all_features[1244]  & \all_features[1245] ;
  assign new_n9352_ = \all_features[1246]  & \all_features[1247]  & (\all_features[1244]  | \all_features[1245]  | new_n9354_ | ~new_n9353_);
  assign new_n9353_ = ~\all_features[1242]  & ~\all_features[1243] ;
  assign new_n9354_ = \all_features[1240]  & \all_features[1241] ;
  assign new_n9355_ = ~\all_features[1243]  & ~\all_features[1244]  & (~\all_features[1242]  | new_n9356_);
  assign new_n9356_ = ~\all_features[1240]  & ~\all_features[1241] ;
  assign new_n9357_ = \all_features[1247]  & (\all_features[1246]  | (\all_features[1245]  & (\all_features[1244]  | ~new_n9353_ | ~new_n9356_)));
  assign new_n9358_ = ~new_n9359_ & ~\all_features[1247] ;
  assign new_n9359_ = \all_features[1245]  & \all_features[1246]  & (\all_features[1244]  | (\all_features[1242]  & \all_features[1243]  & \all_features[1241] ));
  assign new_n9360_ = ~\all_features[1247]  & (~new_n9354_ | ~\all_features[1242]  | ~\all_features[1243]  | ~\all_features[1246]  | ~new_n9351_);
  assign new_n9361_ = \all_features[1247]  & (\all_features[1245]  | \all_features[1246]  | \all_features[1244] );
  assign new_n9362_ = ~new_n9363_ & (\all_features[1243]  | \all_features[1244]  | \all_features[1245]  | \all_features[1246]  | \all_features[1247] );
  assign new_n9363_ = ~\all_features[1245]  & new_n9364_ & ((~\all_features[1242]  & new_n9356_) | ~\all_features[1244]  | ~\all_features[1243] );
  assign new_n9364_ = ~\all_features[1246]  & ~\all_features[1247] ;
  assign new_n9365_ = ~\all_features[1247]  & (~\all_features[1246]  | new_n9366_);
  assign new_n9366_ = ~\all_features[1245]  & (new_n9356_ | ~\all_features[1243]  | ~\all_features[1244]  | ~\all_features[1242] );
  assign new_n9367_ = ~new_n9368_ & ~new_n9369_;
  assign new_n9368_ = new_n9364_ & (~\all_features[1245]  | (~\all_features[1244]  & (~\all_features[1243]  | (~\all_features[1242]  & ~\all_features[1241] ))));
  assign new_n9369_ = new_n9364_ & (~\all_features[1243]  | ~new_n9351_ | (~new_n9354_ & ~\all_features[1242] ));
  assign new_n9370_ = ~\all_features[1247]  & (~\all_features[1246]  | (~\all_features[1245]  & ~\all_features[1244]  & (~\all_features[1243]  | ~\all_features[1242] )));
  assign new_n9371_ = ~new_n9372_ & (\all_features[1243]  | \all_features[1244]  | \all_features[1245]  | \all_features[1246]  | \all_features[1247] );
  assign new_n9372_ = ~new_n9363_ & (new_n9368_ | (~new_n9369_ & (new_n9370_ | (~new_n9365_ & ~new_n9373_))));
  assign new_n9373_ = ~new_n9358_ & (new_n9360_ | (new_n9361_ & (~new_n9357_ | (~new_n9374_ & new_n9350_))));
  assign new_n9374_ = ~\all_features[1245]  & \all_features[1246]  & \all_features[1247]  & (\all_features[1244]  ? new_n9353_ : (new_n9354_ | ~new_n9353_));
  assign new_n9375_ = new_n9376_ & new_n9379_;
  assign new_n9376_ = new_n9367_ & ~new_n9377_ & new_n9362_;
  assign new_n9377_ = ~new_n9370_ & ~new_n9360_ & ~new_n9358_ & ~new_n9365_ & ~new_n9378_;
  assign new_n9378_ = new_n9361_ & new_n9357_ & new_n9350_ & new_n9352_;
  assign new_n9379_ = new_n9362_ & new_n9380_ & ~new_n9358_ & ~new_n9368_;
  assign new_n9380_ = ~new_n9370_ & ~new_n9369_ & ~new_n9365_ & ~new_n9360_;
  assign new_n9381_ = ~new_n9382_ & (~new_n9278_ | ~new_n9277_) & (~new_n9276_ | new_n9345_);
  assign new_n9382_ = new_n9208_ & (new_n9170_ ? new_n9247_ : ~new_n9245_);
  assign new_n9383_ = ~new_n9384_ & ~new_n9607_;
  assign new_n9384_ = ~new_n9546_ & new_n9385_ & (~new_n9545_ | (~new_n9549_ & ~new_n9583_));
  assign new_n9385_ = new_n9386_ & ((~new_n9518_ & new_n9544_) | new_n9485_ | new_n9387_);
  assign new_n9386_ = ~new_n9387_ | ((new_n9422_ | new_n9459_ | ~new_n9456_) & (new_n6662_ | ~new_n9457_ | new_n9456_));
  assign new_n9387_ = new_n9388_ & (~new_n9418_ | ~new_n9414_);
  assign new_n9388_ = ~new_n9389_ & ~new_n9411_;
  assign new_n9389_ = new_n9406_ & ~new_n9410_ & ~new_n9390_ & ~new_n9409_;
  assign new_n9390_ = new_n9391_ & ~new_n9404_ & (~new_n9399_ | ~new_n9405_ | ~new_n9402_ | ~new_n9403_);
  assign new_n9391_ = ~new_n9396_ & ~new_n9392_ & ~new_n9394_;
  assign new_n9392_ = ~new_n9393_ & ~\all_features[5319] ;
  assign new_n9393_ = \all_features[5317]  & \all_features[5318]  & (\all_features[5316]  | (\all_features[5314]  & \all_features[5315]  & \all_features[5313] ));
  assign new_n9394_ = ~\all_features[5319]  & (~\all_features[5318]  | (~\all_features[5316]  & ~\all_features[5317]  & ~new_n9395_));
  assign new_n9395_ = \all_features[5314]  & \all_features[5315] ;
  assign new_n9396_ = ~\all_features[5319]  & (~\all_features[5318]  | ~new_n9397_ | ~new_n9398_ | ~new_n9395_);
  assign new_n9397_ = \all_features[5316]  & \all_features[5317] ;
  assign new_n9398_ = \all_features[5312]  & \all_features[5313] ;
  assign new_n9399_ = \all_features[5319]  & (\all_features[5318]  | (\all_features[5317]  & (\all_features[5316]  | ~new_n9401_ | ~new_n9400_)));
  assign new_n9400_ = ~\all_features[5314]  & ~\all_features[5315] ;
  assign new_n9401_ = ~\all_features[5312]  & ~\all_features[5313] ;
  assign new_n9402_ = \all_features[5319]  & (\all_features[5318]  | (new_n9397_ & (\all_features[5314]  | \all_features[5315]  | \all_features[5313] )));
  assign new_n9403_ = \all_features[5318]  & \all_features[5319]  & (\all_features[5316]  | \all_features[5317]  | new_n9398_ | ~new_n9400_);
  assign new_n9404_ = ~\all_features[5319]  & (~\all_features[5318]  | (~\all_features[5317]  & (new_n9401_ | ~new_n9395_ | ~\all_features[5316] )));
  assign new_n9405_ = \all_features[5319]  & (\all_features[5317]  | \all_features[5318]  | \all_features[5316] );
  assign new_n9406_ = ~new_n9407_ & (\all_features[5315]  | \all_features[5316]  | \all_features[5317]  | \all_features[5318]  | \all_features[5319] );
  assign new_n9407_ = new_n9408_ & (~\all_features[5315]  | ~new_n9397_ | (~\all_features[5314]  & ~new_n9398_));
  assign new_n9408_ = ~\all_features[5318]  & ~\all_features[5319] ;
  assign new_n9409_ = new_n9408_ & (~\all_features[5317]  | (~\all_features[5316]  & (~\all_features[5315]  | (~\all_features[5314]  & ~\all_features[5313] ))));
  assign new_n9410_ = ~\all_features[5317]  & new_n9408_ & ((~\all_features[5314]  & new_n9401_) | ~\all_features[5316]  | ~\all_features[5315] );
  assign new_n9411_ = new_n9391_ & new_n9413_ & ~new_n9404_ & new_n9412_;
  assign new_n9412_ = ~new_n9410_ & (\all_features[5315]  | \all_features[5316]  | \all_features[5317]  | \all_features[5318]  | \all_features[5319] );
  assign new_n9413_ = ~new_n9409_ & ~new_n9407_;
  assign new_n9414_ = new_n9412_ & (~new_n9413_ | (~new_n9415_ & ~new_n9404_ & ~new_n9394_));
  assign new_n9415_ = ~new_n9396_ & ~new_n9392_ & (~new_n9405_ | ~new_n9399_ | new_n9416_);
  assign new_n9416_ = new_n9402_ & new_n9403_ & (new_n9417_ | ~\all_features[5317]  | ~\all_features[5318]  | ~\all_features[5319] );
  assign new_n9417_ = ~\all_features[5315]  & ~\all_features[5316]  & (~\all_features[5314]  | new_n9401_);
  assign new_n9418_ = ~new_n9419_ & (\all_features[5315]  | \all_features[5316]  | \all_features[5317]  | \all_features[5318]  | \all_features[5319] );
  assign new_n9419_ = ~new_n9410_ & (new_n9409_ | (~new_n9407_ & (new_n9394_ | (~new_n9404_ & ~new_n9420_))));
  assign new_n9420_ = ~new_n9392_ & (new_n9396_ | (new_n9405_ & (~new_n9399_ | (~new_n9421_ & new_n9402_))));
  assign new_n9421_ = ~\all_features[5317]  & \all_features[5318]  & \all_features[5319]  & (\all_features[5316]  ? new_n9400_ : (new_n9398_ | ~new_n9400_));
  assign new_n9422_ = new_n9423_ & ~new_n9452_ & ~new_n9455_;
  assign new_n9423_ = ~new_n9424_ & ~new_n9445_;
  assign new_n9424_ = ~new_n9425_ & (\all_features[3187]  | \all_features[3188]  | \all_features[3189]  | \all_features[3190]  | \all_features[3191] );
  assign new_n9425_ = ~new_n9439_ & (new_n9441_ | (~new_n9442_ & (new_n9443_ | (~new_n9426_ & ~new_n9444_))));
  assign new_n9426_ = ~new_n9427_ & (new_n9429_ | (new_n9438_ & (~new_n9433_ | (~new_n9437_ & new_n9436_))));
  assign new_n9427_ = ~new_n9428_ & ~\all_features[3191] ;
  assign new_n9428_ = \all_features[3189]  & \all_features[3190]  & (\all_features[3188]  | (\all_features[3186]  & \all_features[3187]  & \all_features[3185] ));
  assign new_n9429_ = ~\all_features[3191]  & (~\all_features[3190]  | ~new_n9430_ | ~new_n9431_ | ~new_n9432_);
  assign new_n9430_ = \all_features[3184]  & \all_features[3185] ;
  assign new_n9431_ = \all_features[3188]  & \all_features[3189] ;
  assign new_n9432_ = \all_features[3186]  & \all_features[3187] ;
  assign new_n9433_ = \all_features[3191]  & (\all_features[3190]  | (\all_features[3189]  & (\all_features[3188]  | ~new_n9435_ | ~new_n9434_)));
  assign new_n9434_ = ~\all_features[3184]  & ~\all_features[3185] ;
  assign new_n9435_ = ~\all_features[3186]  & ~\all_features[3187] ;
  assign new_n9436_ = \all_features[3191]  & (\all_features[3190]  | (new_n9431_ & (\all_features[3186]  | \all_features[3187]  | \all_features[3185] )));
  assign new_n9437_ = ~\all_features[3189]  & \all_features[3190]  & \all_features[3191]  & (\all_features[3188]  ? new_n9435_ : (new_n9430_ | ~new_n9435_));
  assign new_n9438_ = \all_features[3191]  & (\all_features[3189]  | \all_features[3190]  | \all_features[3188] );
  assign new_n9439_ = ~\all_features[3189]  & new_n9440_ & ((~\all_features[3186]  & new_n9434_) | ~\all_features[3188]  | ~\all_features[3187] );
  assign new_n9440_ = ~\all_features[3190]  & ~\all_features[3191] ;
  assign new_n9441_ = new_n9440_ & (~\all_features[3189]  | (~\all_features[3188]  & (~\all_features[3187]  | (~\all_features[3186]  & ~\all_features[3185] ))));
  assign new_n9442_ = new_n9440_ & (~\all_features[3187]  | ~new_n9431_ | (~\all_features[3186]  & ~new_n9430_));
  assign new_n9443_ = ~\all_features[3191]  & (~\all_features[3190]  | (~\all_features[3188]  & ~\all_features[3189]  & ~new_n9432_));
  assign new_n9444_ = ~\all_features[3191]  & (~\all_features[3190]  | (~\all_features[3189]  & (new_n9434_ | ~new_n9432_ | ~\all_features[3188] )));
  assign new_n9445_ = new_n9451_ & (~new_n9450_ | (~new_n9446_ & ~new_n9443_ & ~new_n9444_));
  assign new_n9446_ = ~new_n9427_ & ~new_n9429_ & (~new_n9438_ | ~new_n9433_ | new_n9447_);
  assign new_n9447_ = new_n9436_ & new_n9448_ & (new_n9449_ | ~\all_features[3189]  | ~\all_features[3190]  | ~\all_features[3191] );
  assign new_n9448_ = \all_features[3190]  & \all_features[3191]  & (\all_features[3188]  | \all_features[3189]  | new_n9430_ | ~new_n9435_);
  assign new_n9449_ = ~\all_features[3187]  & ~\all_features[3188]  & (~\all_features[3186]  | new_n9434_);
  assign new_n9450_ = ~new_n9441_ & ~new_n9442_;
  assign new_n9451_ = ~new_n9439_ & (\all_features[3187]  | \all_features[3188]  | \all_features[3189]  | \all_features[3190]  | \all_features[3191] );
  assign new_n9452_ = new_n9453_ & (~new_n9454_ | (new_n9448_ & new_n9438_ & new_n9433_ & new_n9436_));
  assign new_n9453_ = new_n9450_ & new_n9451_;
  assign new_n9454_ = ~new_n9429_ & ~new_n9427_ & ~new_n9443_ & ~new_n9444_;
  assign new_n9455_ = new_n9453_ & new_n9454_;
  assign new_n9456_ = new_n6426_ & new_n6456_;
  assign new_n9457_ = ~new_n9458_ & ~new_n9340_;
  assign new_n9458_ = new_n9341_ & new_n9314_;
  assign new_n9459_ = ~new_n9460_ & ~new_n9482_;
  assign new_n9460_ = ~new_n9481_ & ~new_n9480_ & ~new_n9479_ & ~new_n9461_ & ~new_n9477_;
  assign new_n9461_ = new_n9465_ & (~new_n9474_ | ~new_n9476_ | ~new_n9462_ | ~new_n9473_);
  assign new_n9462_ = \all_features[1215]  & (\all_features[1214]  | new_n9463_);
  assign new_n9463_ = \all_features[1213]  & (\all_features[1210]  | \all_features[1211]  | \all_features[1212]  | ~new_n9464_);
  assign new_n9464_ = ~\all_features[1208]  & ~\all_features[1209] ;
  assign new_n9465_ = ~new_n9471_ & ~new_n9470_ & ~new_n9466_ & ~new_n9468_;
  assign new_n9466_ = ~\all_features[1215]  & (~\all_features[1214]  | (~\all_features[1213]  & (new_n9464_ | ~new_n9467_ | ~\all_features[1212] )));
  assign new_n9467_ = \all_features[1210]  & \all_features[1211] ;
  assign new_n9468_ = ~new_n9469_ & ~\all_features[1215] ;
  assign new_n9469_ = \all_features[1213]  & \all_features[1214]  & (\all_features[1212]  | (\all_features[1210]  & \all_features[1211]  & \all_features[1209] ));
  assign new_n9470_ = ~\all_features[1215]  & (~\all_features[1214]  | (~\all_features[1212]  & ~\all_features[1213]  & ~new_n9467_));
  assign new_n9471_ = ~\all_features[1215]  & (~new_n9467_ | ~\all_features[1208]  | ~\all_features[1209]  | ~\all_features[1214]  | ~new_n9472_);
  assign new_n9472_ = \all_features[1212]  & \all_features[1213] ;
  assign new_n9473_ = \all_features[1215]  & (\all_features[1214]  | (new_n9472_ & (\all_features[1210]  | \all_features[1211]  | \all_features[1209] )));
  assign new_n9474_ = \all_features[1215]  & ~new_n9475_ & \all_features[1214] ;
  assign new_n9475_ = ~\all_features[1210]  & ~\all_features[1211]  & ~\all_features[1212]  & ~\all_features[1213]  & (~\all_features[1209]  | ~\all_features[1208] );
  assign new_n9476_ = \all_features[1215]  & (\all_features[1213]  | \all_features[1214]  | \all_features[1212] );
  assign new_n9477_ = new_n9478_ & (~\all_features[1213]  | (~\all_features[1212]  & (~\all_features[1211]  | (~\all_features[1210]  & ~\all_features[1209] ))));
  assign new_n9478_ = ~\all_features[1214]  & ~\all_features[1215] ;
  assign new_n9479_ = ~\all_features[1213]  & new_n9478_ & ((~\all_features[1210]  & new_n9464_) | ~\all_features[1212]  | ~\all_features[1211] );
  assign new_n9480_ = new_n9478_ & (~new_n9472_ | ~\all_features[1211]  | (~\all_features[1210]  & (~\all_features[1208]  | ~\all_features[1209] )));
  assign new_n9481_ = ~\all_features[1215]  & ~\all_features[1214]  & ~\all_features[1213]  & ~\all_features[1211]  & ~\all_features[1212] ;
  assign new_n9482_ = new_n9484_ & new_n9483_ & ~new_n9479_ & ~new_n9471_ & ~new_n9466_ & ~new_n9468_;
  assign new_n9483_ = ~new_n9470_ & ~new_n9481_;
  assign new_n9484_ = ~new_n9477_ & ~new_n9480_;
  assign new_n9485_ = ~new_n9514_ & (~new_n9516_ | (~new_n9507_ & ~new_n9486_));
  assign new_n9486_ = ~new_n9487_ & (\all_features[2283]  | \all_features[2284]  | \all_features[2285]  | \all_features[2286]  | \all_features[2287] );
  assign new_n9487_ = ~new_n9503_ & (new_n9501_ | (~new_n9505_ & (new_n9506_ | (~new_n9504_ & ~new_n9488_))));
  assign new_n9488_ = ~new_n9489_ & (new_n9491_ | (new_n9500_ & (~new_n9495_ | (~new_n9499_ & new_n9498_))));
  assign new_n9489_ = ~new_n9490_ & ~\all_features[2287] ;
  assign new_n9490_ = \all_features[2285]  & \all_features[2286]  & (\all_features[2284]  | (\all_features[2282]  & \all_features[2283]  & \all_features[2281] ));
  assign new_n9491_ = ~\all_features[2287]  & (~\all_features[2286]  | ~new_n9492_ | ~new_n9493_ | ~new_n9494_);
  assign new_n9492_ = \all_features[2282]  & \all_features[2283] ;
  assign new_n9493_ = \all_features[2280]  & \all_features[2281] ;
  assign new_n9494_ = \all_features[2284]  & \all_features[2285] ;
  assign new_n9495_ = \all_features[2287]  & (\all_features[2286]  | (\all_features[2285]  & (\all_features[2284]  | ~new_n9497_ | ~new_n9496_)));
  assign new_n9496_ = ~\all_features[2280]  & ~\all_features[2281] ;
  assign new_n9497_ = ~\all_features[2282]  & ~\all_features[2283] ;
  assign new_n9498_ = \all_features[2287]  & (\all_features[2286]  | (new_n9494_ & (\all_features[2282]  | \all_features[2283]  | \all_features[2281] )));
  assign new_n9499_ = ~\all_features[2285]  & \all_features[2286]  & \all_features[2287]  & (\all_features[2284]  ? new_n9497_ : (new_n9493_ | ~new_n9497_));
  assign new_n9500_ = \all_features[2287]  & (\all_features[2285]  | \all_features[2286]  | \all_features[2284] );
  assign new_n9501_ = new_n9502_ & (~\all_features[2285]  | (~\all_features[2284]  & (~\all_features[2283]  | (~\all_features[2282]  & ~\all_features[2281] ))));
  assign new_n9502_ = ~\all_features[2286]  & ~\all_features[2287] ;
  assign new_n9503_ = ~\all_features[2285]  & new_n9502_ & ((~\all_features[2282]  & new_n9496_) | ~\all_features[2284]  | ~\all_features[2283] );
  assign new_n9504_ = ~\all_features[2287]  & (~\all_features[2286]  | (~\all_features[2285]  & (new_n9496_ | ~new_n9492_ | ~\all_features[2284] )));
  assign new_n9505_ = new_n9502_ & (~\all_features[2283]  | ~new_n9494_ | (~\all_features[2282]  & ~new_n9493_));
  assign new_n9506_ = ~\all_features[2287]  & (~\all_features[2286]  | (~\all_features[2284]  & ~\all_features[2285]  & ~new_n9492_));
  assign new_n9507_ = new_n9512_ & (~new_n9513_ | (~new_n9508_ & ~new_n9504_ & ~new_n9506_));
  assign new_n9508_ = ~new_n9489_ & ~new_n9491_ & (~new_n9500_ | ~new_n9495_ | new_n9509_);
  assign new_n9509_ = new_n9498_ & new_n9510_ & (new_n9511_ | ~\all_features[2285]  | ~\all_features[2286]  | ~\all_features[2287] );
  assign new_n9510_ = \all_features[2286]  & \all_features[2287]  & (\all_features[2284]  | \all_features[2285]  | new_n9493_ | ~new_n9497_);
  assign new_n9511_ = ~\all_features[2283]  & ~\all_features[2284]  & (~\all_features[2282]  | new_n9496_);
  assign new_n9512_ = ~new_n9503_ & (\all_features[2283]  | \all_features[2284]  | \all_features[2285]  | \all_features[2286]  | \all_features[2287] );
  assign new_n9513_ = ~new_n9501_ & ~new_n9505_;
  assign new_n9514_ = new_n9515_ & new_n9512_ & ~new_n9505_ & ~new_n9504_ & ~new_n9489_ & ~new_n9501_;
  assign new_n9515_ = ~new_n9491_ & ~new_n9506_;
  assign new_n9516_ = new_n9512_ & new_n9513_ & (new_n9517_ | new_n9489_ | new_n9504_ | ~new_n9515_);
  assign new_n9517_ = new_n9500_ & new_n9510_ & new_n9495_ & new_n9498_;
  assign new_n9518_ = ~new_n9541_ | (~new_n9519_ & new_n9537_ & new_n9536_);
  assign new_n9519_ = new_n9520_ & (new_n9533_ | new_n9535_ | (new_n9525_ & (new_n9527_ | ~new_n9529_)));
  assign new_n9520_ = ~new_n9521_ & ~new_n9523_;
  assign new_n9521_ = ~\all_features[3999]  & (~\all_features[3998]  | (~\all_features[3996]  & ~\all_features[3997]  & ~new_n9522_));
  assign new_n9522_ = \all_features[3994]  & \all_features[3995] ;
  assign new_n9523_ = ~\all_features[3999]  & (~\all_features[3998]  | (~\all_features[3997]  & (new_n9524_ | ~\all_features[3996]  | ~new_n9522_)));
  assign new_n9524_ = ~\all_features[3992]  & ~\all_features[3993] ;
  assign new_n9525_ = \all_features[3999]  & (\all_features[3998]  | (~new_n9526_ & \all_features[3997] ));
  assign new_n9526_ = new_n9524_ & ~\all_features[3996]  & ~\all_features[3994]  & ~\all_features[3995] ;
  assign new_n9527_ = \all_features[3999]  & \all_features[3998]  & ~new_n9528_ & \all_features[3997] ;
  assign new_n9528_ = ~\all_features[3995]  & ~\all_features[3996]  & (~\all_features[3994]  | new_n9524_);
  assign new_n9529_ = \all_features[3999]  & \all_features[3998]  & ~new_n9532_ & new_n9530_;
  assign new_n9530_ = \all_features[3999]  & (\all_features[3998]  | (new_n9531_ & (\all_features[3994]  | \all_features[3995]  | \all_features[3993] )));
  assign new_n9531_ = \all_features[3996]  & \all_features[3997] ;
  assign new_n9532_ = ~\all_features[3994]  & ~\all_features[3995]  & ~\all_features[3996]  & ~\all_features[3997]  & (~\all_features[3993]  | ~\all_features[3992] );
  assign new_n9533_ = ~new_n9534_ & ~\all_features[3999] ;
  assign new_n9534_ = \all_features[3997]  & \all_features[3998]  & (\all_features[3996]  | (\all_features[3994]  & \all_features[3995]  & \all_features[3993] ));
  assign new_n9535_ = ~\all_features[3999]  & (~new_n9531_ | ~\all_features[3992]  | ~\all_features[3993]  | ~\all_features[3998]  | ~new_n9522_);
  assign new_n9536_ = ~new_n9521_ & ~new_n9523_ & ~new_n9533_ & ~new_n9535_ & (~new_n9529_ | ~new_n9525_);
  assign new_n9537_ = ~new_n9538_ & ~new_n9540_;
  assign new_n9538_ = new_n9539_ & (~new_n9531_ | ~\all_features[3995]  | (~\all_features[3994]  & (~\all_features[3992]  | ~\all_features[3993] )));
  assign new_n9539_ = ~\all_features[3998]  & ~\all_features[3999] ;
  assign new_n9540_ = new_n9539_ & (~\all_features[3997]  | (~\all_features[3996]  & (~\all_features[3995]  | (~\all_features[3994]  & ~\all_features[3993] ))));
  assign new_n9541_ = ~new_n9542_ & ~new_n9543_;
  assign new_n9542_ = ~\all_features[3997]  & new_n9539_ & ((~\all_features[3994]  & new_n9524_) | ~\all_features[3996]  | ~\all_features[3995] );
  assign new_n9543_ = ~\all_features[3999]  & ~\all_features[3998]  & ~\all_features[3997]  & ~\all_features[3995]  & ~\all_features[3996] ;
  assign new_n9544_ = new_n9537_ & new_n9520_ & new_n9541_ & ~new_n9533_ & ~new_n9535_;
  assign new_n9545_ = ~new_n9387_ & new_n9485_;
  assign new_n9546_ = new_n9387_ & ((~new_n9547_ & new_n9422_ & new_n9456_) | (~new_n9456_ & (new_n6662_ | ~new_n9457_)));
  assign new_n9547_ = new_n9548_ & new_n7475_;
  assign new_n9548_ = new_n7447_ & new_n7477_;
  assign new_n9549_ = new_n9579_ & (new_n9581_ | new_n9550_);
  assign new_n9550_ = new_n9551_ & new_n9572_;
  assign new_n9551_ = ~new_n9552_ & (\all_features[3659]  | \all_features[3660]  | \all_features[3661]  | \all_features[3662]  | \all_features[3663] );
  assign new_n9552_ = ~new_n9568_ & (new_n9566_ | (~new_n9570_ & (new_n9571_ | (~new_n9569_ & ~new_n9553_))));
  assign new_n9553_ = ~new_n9554_ & (new_n9556_ | (new_n9565_ & (~new_n9560_ | (~new_n9564_ & new_n9563_))));
  assign new_n9554_ = ~new_n9555_ & ~\all_features[3663] ;
  assign new_n9555_ = \all_features[3661]  & \all_features[3662]  & (\all_features[3660]  | (\all_features[3658]  & \all_features[3659]  & \all_features[3657] ));
  assign new_n9556_ = ~\all_features[3663]  & (~\all_features[3662]  | ~new_n9557_ | ~new_n9558_ | ~new_n9559_);
  assign new_n9557_ = \all_features[3658]  & \all_features[3659] ;
  assign new_n9558_ = \all_features[3656]  & \all_features[3657] ;
  assign new_n9559_ = \all_features[3660]  & \all_features[3661] ;
  assign new_n9560_ = \all_features[3663]  & (\all_features[3662]  | (\all_features[3661]  & (\all_features[3660]  | ~new_n9562_ | ~new_n9561_)));
  assign new_n9561_ = ~\all_features[3656]  & ~\all_features[3657] ;
  assign new_n9562_ = ~\all_features[3658]  & ~\all_features[3659] ;
  assign new_n9563_ = \all_features[3663]  & (\all_features[3662]  | (new_n9559_ & (\all_features[3658]  | \all_features[3659]  | \all_features[3657] )));
  assign new_n9564_ = ~\all_features[3661]  & \all_features[3662]  & \all_features[3663]  & (\all_features[3660]  ? new_n9562_ : (new_n9558_ | ~new_n9562_));
  assign new_n9565_ = \all_features[3663]  & (\all_features[3661]  | \all_features[3662]  | \all_features[3660] );
  assign new_n9566_ = new_n9567_ & (~\all_features[3661]  | (~\all_features[3660]  & (~\all_features[3659]  | (~\all_features[3658]  & ~\all_features[3657] ))));
  assign new_n9567_ = ~\all_features[3662]  & ~\all_features[3663] ;
  assign new_n9568_ = ~\all_features[3661]  & new_n9567_ & ((~\all_features[3658]  & new_n9561_) | ~\all_features[3660]  | ~\all_features[3659] );
  assign new_n9569_ = ~\all_features[3663]  & (~\all_features[3662]  | (~\all_features[3661]  & (new_n9561_ | ~new_n9557_ | ~\all_features[3660] )));
  assign new_n9570_ = new_n9567_ & (~\all_features[3659]  | ~new_n9559_ | (~\all_features[3658]  & ~new_n9558_));
  assign new_n9571_ = ~\all_features[3663]  & (~\all_features[3662]  | (~\all_features[3660]  & ~\all_features[3661]  & ~new_n9557_));
  assign new_n9572_ = new_n9577_ & (~new_n9578_ | (~new_n9573_ & ~new_n9569_ & ~new_n9571_));
  assign new_n9573_ = ~new_n9554_ & ~new_n9556_ & (~new_n9565_ | ~new_n9560_ | new_n9574_);
  assign new_n9574_ = new_n9563_ & new_n9575_ & (new_n9576_ | ~\all_features[3661]  | ~\all_features[3662]  | ~\all_features[3663] );
  assign new_n9575_ = \all_features[3662]  & \all_features[3663]  & (\all_features[3660]  | \all_features[3661]  | new_n9558_ | ~new_n9562_);
  assign new_n9576_ = ~\all_features[3659]  & ~\all_features[3660]  & (~\all_features[3658]  | new_n9561_);
  assign new_n9577_ = ~new_n9568_ & (\all_features[3659]  | \all_features[3660]  | \all_features[3661]  | \all_features[3662]  | \all_features[3663] );
  assign new_n9578_ = ~new_n9566_ & ~new_n9570_;
  assign new_n9579_ = new_n9580_ & new_n9577_ & ~new_n9570_ & ~new_n9569_ & ~new_n9554_ & ~new_n9566_;
  assign new_n9580_ = ~new_n9556_ & ~new_n9571_;
  assign new_n9581_ = new_n9577_ & new_n9578_ & (new_n9582_ | new_n9554_ | new_n9569_ | ~new_n9580_);
  assign new_n9582_ = new_n9565_ & new_n9575_ & new_n9560_ & new_n9563_;
  assign new_n9583_ = ~new_n9584_ & ~new_n9606_;
  assign new_n9584_ = new_n9585_ & (~new_n9594_ | (new_n9604_ & new_n9605_ & new_n9601_ & new_n9603_));
  assign new_n9585_ = new_n9586_ & ~new_n9590_ & ~new_n9591_;
  assign new_n9586_ = ~new_n9587_ & (\all_features[2627]  | \all_features[2628]  | \all_features[2629]  | \all_features[2630]  | \all_features[2631] );
  assign new_n9587_ = ~\all_features[2629]  & new_n9589_ & ((~\all_features[2626]  & new_n9588_) | ~\all_features[2628]  | ~\all_features[2627] );
  assign new_n9588_ = ~\all_features[2624]  & ~\all_features[2625] ;
  assign new_n9589_ = ~\all_features[2630]  & ~\all_features[2631] ;
  assign new_n9590_ = new_n9589_ & (~\all_features[2629]  | (~\all_features[2628]  & (~\all_features[2627]  | (~\all_features[2626]  & ~\all_features[2625] ))));
  assign new_n9591_ = new_n9589_ & (~\all_features[2627]  | ~new_n9592_ | (~\all_features[2626]  & ~new_n9593_));
  assign new_n9592_ = \all_features[2628]  & \all_features[2629] ;
  assign new_n9593_ = \all_features[2624]  & \all_features[2625] ;
  assign new_n9594_ = ~new_n9600_ & ~new_n9599_ & ~new_n9595_ & ~new_n9597_;
  assign new_n9595_ = ~\all_features[2631]  & (~\all_features[2630]  | (~\all_features[2629]  & (new_n9588_ | ~new_n9596_ | ~\all_features[2628] )));
  assign new_n9596_ = \all_features[2626]  & \all_features[2627] ;
  assign new_n9597_ = ~new_n9598_ & ~\all_features[2631] ;
  assign new_n9598_ = \all_features[2629]  & \all_features[2630]  & (\all_features[2628]  | (\all_features[2626]  & \all_features[2627]  & \all_features[2625] ));
  assign new_n9599_ = ~\all_features[2631]  & (~\all_features[2630]  | ~new_n9592_ | ~new_n9593_ | ~new_n9596_);
  assign new_n9600_ = ~\all_features[2631]  & (~\all_features[2630]  | (~\all_features[2628]  & ~\all_features[2629]  & ~new_n9596_));
  assign new_n9601_ = \all_features[2631]  & (\all_features[2630]  | (\all_features[2629]  & (\all_features[2628]  | ~new_n9588_ | ~new_n9602_)));
  assign new_n9602_ = ~\all_features[2626]  & ~\all_features[2627] ;
  assign new_n9603_ = \all_features[2631]  & (\all_features[2630]  | (new_n9592_ & (\all_features[2626]  | \all_features[2627]  | \all_features[2625] )));
  assign new_n9604_ = \all_features[2630]  & \all_features[2631]  & (\all_features[2628]  | \all_features[2629]  | new_n9593_ | ~new_n9602_);
  assign new_n9605_ = \all_features[2631]  & (\all_features[2629]  | \all_features[2630]  | \all_features[2628] );
  assign new_n9606_ = new_n9585_ & new_n9594_;
  assign new_n9607_ = new_n9545_ & ~new_n9549_ & ~new_n9583_;
  assign new_n9608_ = new_n9609_ & (new_n9832_ | new_n9688_ | new_n8701_);
  assign new_n9609_ = ~new_n9651_ & (new_n9687_ | ((new_n9797_ | ~new_n9759_ | ~new_n9761_) & (new_n9610_ | new_n9761_)));
  assign new_n9610_ = (~new_n9649_ & (~new_n9644_ | ~new_n9650_) & (~new_n9611_ | ~new_n9635_)) | (new_n9170_ & new_n9611_ & new_n9635_);
  assign new_n9611_ = ~new_n9612_ & ~new_n9634_;
  assign new_n9612_ = new_n9613_ & (~new_n9622_ | (new_n9632_ & new_n9633_ & new_n9629_ & new_n9631_));
  assign new_n9613_ = new_n9614_ & ~new_n9618_ & ~new_n9619_;
  assign new_n9614_ = ~new_n9615_ & (\all_features[5243]  | \all_features[5244]  | \all_features[5245]  | \all_features[5246]  | \all_features[5247] );
  assign new_n9615_ = ~\all_features[5245]  & new_n9617_ & ((~\all_features[5242]  & new_n9616_) | ~\all_features[5244]  | ~\all_features[5243] );
  assign new_n9616_ = ~\all_features[5240]  & ~\all_features[5241] ;
  assign new_n9617_ = ~\all_features[5246]  & ~\all_features[5247] ;
  assign new_n9618_ = new_n9617_ & (~\all_features[5245]  | (~\all_features[5244]  & (~\all_features[5243]  | (~\all_features[5242]  & ~\all_features[5241] ))));
  assign new_n9619_ = new_n9617_ & (~\all_features[5243]  | ~new_n9620_ | (~\all_features[5242]  & ~new_n9621_));
  assign new_n9620_ = \all_features[5244]  & \all_features[5245] ;
  assign new_n9621_ = \all_features[5240]  & \all_features[5241] ;
  assign new_n9622_ = ~new_n9628_ & ~new_n9627_ & ~new_n9623_ & ~new_n9625_;
  assign new_n9623_ = ~\all_features[5247]  & (~\all_features[5246]  | (~\all_features[5245]  & (new_n9616_ | ~new_n9624_ | ~\all_features[5244] )));
  assign new_n9624_ = \all_features[5242]  & \all_features[5243] ;
  assign new_n9625_ = ~new_n9626_ & ~\all_features[5247] ;
  assign new_n9626_ = \all_features[5245]  & \all_features[5246]  & (\all_features[5244]  | (\all_features[5242]  & \all_features[5243]  & \all_features[5241] ));
  assign new_n9627_ = ~\all_features[5247]  & (~\all_features[5246]  | ~new_n9620_ | ~new_n9621_ | ~new_n9624_);
  assign new_n9628_ = ~\all_features[5247]  & (~\all_features[5246]  | (~\all_features[5244]  & ~\all_features[5245]  & ~new_n9624_));
  assign new_n9629_ = \all_features[5247]  & (\all_features[5246]  | (\all_features[5245]  & (\all_features[5244]  | ~new_n9616_ | ~new_n9630_)));
  assign new_n9630_ = ~\all_features[5242]  & ~\all_features[5243] ;
  assign new_n9631_ = \all_features[5247]  & (\all_features[5246]  | (new_n9620_ & (\all_features[5242]  | \all_features[5243]  | \all_features[5241] )));
  assign new_n9632_ = \all_features[5246]  & \all_features[5247]  & (\all_features[5244]  | \all_features[5245]  | new_n9621_ | ~new_n9630_);
  assign new_n9633_ = \all_features[5247]  & (\all_features[5245]  | \all_features[5246]  | \all_features[5244] );
  assign new_n9634_ = new_n9613_ & new_n9622_;
  assign new_n9635_ = ~new_n9636_ & ~new_n9640_;
  assign new_n9636_ = ~new_n9637_ & (\all_features[5243]  | \all_features[5244]  | \all_features[5245]  | \all_features[5246]  | \all_features[5247] );
  assign new_n9637_ = ~new_n9615_ & (new_n9618_ | (~new_n9619_ & (new_n9628_ | (~new_n9623_ & ~new_n9638_))));
  assign new_n9638_ = ~new_n9625_ & (new_n9627_ | (new_n9633_ & (~new_n9629_ | (~new_n9639_ & new_n9631_))));
  assign new_n9639_ = ~\all_features[5245]  & \all_features[5246]  & \all_features[5247]  & (\all_features[5244]  ? new_n9630_ : (new_n9621_ | ~new_n9630_));
  assign new_n9640_ = new_n9614_ & (new_n9619_ | new_n9618_ | (~new_n9623_ & ~new_n9628_ & ~new_n9641_));
  assign new_n9641_ = ~new_n9627_ & ~new_n9625_ & (~new_n9633_ | ~new_n9629_ | new_n9642_);
  assign new_n9642_ = new_n9631_ & new_n9632_ & (new_n9643_ | ~\all_features[5245]  | ~\all_features[5246]  | ~\all_features[5247] );
  assign new_n9643_ = ~\all_features[5243]  & ~\all_features[5244]  & (~\all_features[5242]  | new_n9616_);
  assign new_n9644_ = new_n8031_ & new_n9645_;
  assign new_n9645_ = ~new_n9646_ & (\all_features[3923]  | \all_features[3924]  | \all_features[3925]  | \all_features[3926]  | \all_features[3927] );
  assign new_n9646_ = ~new_n8053_ & (new_n8049_ | (~new_n8047_ & (new_n8054_ | (~new_n8050_ & ~new_n9647_))));
  assign new_n9647_ = ~new_n8043_ & (new_n8042_ | (new_n8045_ & (~new_n8041_ | (~new_n9648_ & new_n8034_))));
  assign new_n9648_ = ~\all_features[3925]  & \all_features[3926]  & \all_features[3927]  & (\all_features[3924]  ? new_n8038_ : (new_n8037_ | ~new_n8038_));
  assign new_n9649_ = new_n8056_ & new_n8059_;
  assign new_n9650_ = ~new_n8056_ & new_n8059_;
  assign new_n9651_ = new_n9725_ & new_n9687_ & ~new_n9652_ & ~new_n9689_;
  assign new_n9652_ = ~new_n9653_ & ~new_n9686_;
  assign new_n9653_ = new_n9654_ & new_n9682_;
  assign new_n9654_ = new_n9655_ & new_n9679_;
  assign new_n9655_ = new_n9671_ & (~new_n9674_ | (~new_n9656_ & ~new_n9677_ & ~new_n9678_));
  assign new_n9656_ = ~new_n9665_ & ~new_n9667_ & (~new_n9670_ | ~new_n9669_ | new_n9657_);
  assign new_n9657_ = new_n9658_ & new_n9660_ & (new_n9663_ | ~\all_features[1909]  | ~\all_features[1910]  | ~\all_features[1911] );
  assign new_n9658_ = \all_features[1911]  & (\all_features[1910]  | (new_n9659_ & (\all_features[1906]  | \all_features[1907]  | \all_features[1905] )));
  assign new_n9659_ = \all_features[1908]  & \all_features[1909] ;
  assign new_n9660_ = \all_features[1910]  & \all_features[1911]  & (\all_features[1908]  | \all_features[1909]  | new_n9661_ | ~new_n9662_);
  assign new_n9661_ = \all_features[1904]  & \all_features[1905] ;
  assign new_n9662_ = ~\all_features[1906]  & ~\all_features[1907] ;
  assign new_n9663_ = ~\all_features[1907]  & ~\all_features[1908]  & (~\all_features[1906]  | new_n9664_);
  assign new_n9664_ = ~\all_features[1904]  & ~\all_features[1905] ;
  assign new_n9665_ = ~new_n9666_ & ~\all_features[1911] ;
  assign new_n9666_ = \all_features[1909]  & \all_features[1910]  & (\all_features[1908]  | (\all_features[1906]  & \all_features[1907]  & \all_features[1905] ));
  assign new_n9667_ = ~\all_features[1911]  & (~\all_features[1910]  | ~new_n9668_ | ~new_n9661_ | ~new_n9659_);
  assign new_n9668_ = \all_features[1906]  & \all_features[1907] ;
  assign new_n9669_ = \all_features[1911]  & (\all_features[1910]  | (\all_features[1909]  & (\all_features[1908]  | ~new_n9662_ | ~new_n9664_)));
  assign new_n9670_ = \all_features[1911]  & (\all_features[1909]  | \all_features[1910]  | \all_features[1908] );
  assign new_n9671_ = ~new_n9672_ & (\all_features[1907]  | \all_features[1908]  | \all_features[1909]  | \all_features[1910]  | \all_features[1911] );
  assign new_n9672_ = ~\all_features[1909]  & new_n9673_ & ((~\all_features[1906]  & new_n9664_) | ~\all_features[1908]  | ~\all_features[1907] );
  assign new_n9673_ = ~\all_features[1910]  & ~\all_features[1911] ;
  assign new_n9674_ = ~new_n9675_ & ~new_n9676_;
  assign new_n9675_ = new_n9673_ & (~\all_features[1909]  | (~\all_features[1908]  & (~\all_features[1907]  | (~\all_features[1906]  & ~\all_features[1905] ))));
  assign new_n9676_ = new_n9673_ & (~\all_features[1907]  | ~new_n9659_ | (~\all_features[1906]  & ~new_n9661_));
  assign new_n9677_ = ~\all_features[1911]  & (~\all_features[1910]  | (~\all_features[1909]  & (new_n9664_ | ~new_n9668_ | ~\all_features[1908] )));
  assign new_n9678_ = ~\all_features[1911]  & (~\all_features[1910]  | (~\all_features[1908]  & ~\all_features[1909]  & ~new_n9668_));
  assign new_n9679_ = new_n9671_ & new_n9674_ & (new_n9681_ | new_n9665_ | new_n9677_ | ~new_n9680_);
  assign new_n9680_ = ~new_n9667_ & ~new_n9678_;
  assign new_n9681_ = new_n9670_ & new_n9660_ & new_n9669_ & new_n9658_;
  assign new_n9682_ = ~new_n9683_ & (\all_features[1907]  | \all_features[1908]  | \all_features[1909]  | \all_features[1910]  | \all_features[1911] );
  assign new_n9683_ = ~new_n9672_ & (new_n9675_ | (~new_n9676_ & (new_n9678_ | (~new_n9677_ & ~new_n9684_))));
  assign new_n9684_ = ~new_n9665_ & (new_n9667_ | (new_n9670_ & (~new_n9669_ | (~new_n9685_ & new_n9658_))));
  assign new_n9685_ = ~\all_features[1909]  & \all_features[1910]  & \all_features[1911]  & (\all_features[1908]  ? new_n9662_ : (new_n9661_ | ~new_n9662_));
  assign new_n9686_ = new_n9680_ & new_n9671_ & ~new_n9676_ & ~new_n9677_ & ~new_n9665_ & ~new_n9675_;
  assign new_n9687_ = ~new_n9688_ & ~new_n8701_;
  assign new_n9688_ = new_n8669_ & new_n8698_;
  assign new_n9689_ = ~new_n9690_ & new_n9720_;
  assign new_n9690_ = new_n9691_ & new_n9712_;
  assign new_n9691_ = ~new_n9692_ & (\all_features[3019]  | \all_features[3020]  | \all_features[3021]  | \all_features[3022]  | \all_features[3023] );
  assign new_n9692_ = ~new_n9706_ & (new_n9711_ | (~new_n9708_ & (new_n9709_ | (~new_n9710_ & ~new_n9693_))));
  assign new_n9693_ = ~new_n9694_ & (new_n9703_ | (new_n9705_ & (~new_n9696_ | (~new_n9701_ & new_n9699_))));
  assign new_n9694_ = ~new_n9695_ & ~\all_features[3023] ;
  assign new_n9695_ = \all_features[3021]  & \all_features[3022]  & (\all_features[3020]  | (\all_features[3018]  & \all_features[3019]  & \all_features[3017] ));
  assign new_n9696_ = \all_features[3023]  & (\all_features[3022]  | (\all_features[3021]  & (\all_features[3020]  | ~new_n9698_ | ~new_n9697_)));
  assign new_n9697_ = ~\all_features[3016]  & ~\all_features[3017] ;
  assign new_n9698_ = ~\all_features[3018]  & ~\all_features[3019] ;
  assign new_n9699_ = \all_features[3023]  & (\all_features[3022]  | (new_n9700_ & (\all_features[3018]  | \all_features[3019]  | \all_features[3017] )));
  assign new_n9700_ = \all_features[3020]  & \all_features[3021] ;
  assign new_n9701_ = ~\all_features[3021]  & \all_features[3022]  & \all_features[3023]  & (\all_features[3020]  ? new_n9698_ : (new_n9702_ | ~new_n9698_));
  assign new_n9702_ = \all_features[3016]  & \all_features[3017] ;
  assign new_n9703_ = ~\all_features[3023]  & (~\all_features[3022]  | ~new_n9702_ | ~new_n9700_ | ~new_n9704_);
  assign new_n9704_ = \all_features[3018]  & \all_features[3019] ;
  assign new_n9705_ = \all_features[3023]  & (\all_features[3021]  | \all_features[3022]  | \all_features[3020] );
  assign new_n9706_ = ~\all_features[3021]  & new_n9707_ & ((~\all_features[3018]  & new_n9697_) | ~\all_features[3020]  | ~\all_features[3019] );
  assign new_n9707_ = ~\all_features[3022]  & ~\all_features[3023] ;
  assign new_n9708_ = new_n9707_ & (~\all_features[3019]  | ~new_n9700_ | (~\all_features[3018]  & ~new_n9702_));
  assign new_n9709_ = ~\all_features[3023]  & (~\all_features[3022]  | (~\all_features[3020]  & ~\all_features[3021]  & ~new_n9704_));
  assign new_n9710_ = ~\all_features[3023]  & (~\all_features[3022]  | (~\all_features[3021]  & (new_n9697_ | ~new_n9704_ | ~\all_features[3020] )));
  assign new_n9711_ = new_n9707_ & (~\all_features[3021]  | (~\all_features[3020]  & (~\all_features[3019]  | (~\all_features[3018]  & ~\all_features[3017] ))));
  assign new_n9712_ = new_n9718_ & (~new_n9719_ | (~new_n9713_ & ~new_n9709_ & ~new_n9710_));
  assign new_n9713_ = new_n9716_ & ((~new_n9714_ & new_n9699_ & new_n9717_) | ~new_n9705_ | ~new_n9696_);
  assign new_n9714_ = \all_features[3023]  & \all_features[3022]  & ~new_n9715_ & \all_features[3021] ;
  assign new_n9715_ = ~\all_features[3019]  & ~\all_features[3020]  & (~\all_features[3018]  | new_n9697_);
  assign new_n9716_ = ~new_n9694_ & ~new_n9703_;
  assign new_n9717_ = \all_features[3022]  & \all_features[3023]  & (\all_features[3020]  | \all_features[3021]  | new_n9702_ | ~new_n9698_);
  assign new_n9718_ = ~new_n9706_ & (\all_features[3019]  | \all_features[3020]  | \all_features[3021]  | \all_features[3022]  | \all_features[3023] );
  assign new_n9719_ = ~new_n9708_ & ~new_n9711_;
  assign new_n9720_ = ~new_n9721_ & ~new_n9724_;
  assign new_n9721_ = new_n9719_ & ~new_n9722_ & new_n9718_;
  assign new_n9722_ = new_n9723_ & (~new_n9717_ | ~new_n9705_ | ~new_n9696_ | ~new_n9699_);
  assign new_n9723_ = ~new_n9703_ & ~new_n9694_ & ~new_n9709_ & ~new_n9710_;
  assign new_n9724_ = new_n9716_ & new_n9718_ & ~new_n9711_ & ~new_n9710_ & ~new_n9708_ & ~new_n9709_;
  assign new_n9725_ = new_n9726_ & new_n9750_;
  assign new_n9726_ = ~new_n9727_ & ~new_n9749_;
  assign new_n9727_ = new_n9728_ & (~new_n9737_ | (new_n9747_ & new_n9748_ & new_n9744_ & new_n9746_));
  assign new_n9728_ = new_n9729_ & ~new_n9733_ & ~new_n9734_;
  assign new_n9729_ = ~new_n9730_ & (\all_features[1931]  | \all_features[1932]  | \all_features[1933]  | \all_features[1934]  | \all_features[1935] );
  assign new_n9730_ = ~\all_features[1933]  & new_n9732_ & ((~\all_features[1930]  & new_n9731_) | ~\all_features[1932]  | ~\all_features[1931] );
  assign new_n9731_ = ~\all_features[1928]  & ~\all_features[1929] ;
  assign new_n9732_ = ~\all_features[1934]  & ~\all_features[1935] ;
  assign new_n9733_ = new_n9732_ & (~\all_features[1933]  | (~\all_features[1932]  & (~\all_features[1931]  | (~\all_features[1930]  & ~\all_features[1929] ))));
  assign new_n9734_ = new_n9732_ & (~\all_features[1931]  | ~new_n9735_ | (~\all_features[1930]  & ~new_n9736_));
  assign new_n9735_ = \all_features[1932]  & \all_features[1933] ;
  assign new_n9736_ = \all_features[1928]  & \all_features[1929] ;
  assign new_n9737_ = ~new_n9743_ & ~new_n9742_ & ~new_n9738_ & ~new_n9740_;
  assign new_n9738_ = ~\all_features[1935]  & (~\all_features[1934]  | (~\all_features[1933]  & (new_n9731_ | ~new_n9739_ | ~\all_features[1932] )));
  assign new_n9739_ = \all_features[1930]  & \all_features[1931] ;
  assign new_n9740_ = ~new_n9741_ & ~\all_features[1935] ;
  assign new_n9741_ = \all_features[1933]  & \all_features[1934]  & (\all_features[1932]  | (\all_features[1930]  & \all_features[1931]  & \all_features[1929] ));
  assign new_n9742_ = ~\all_features[1935]  & (~\all_features[1934]  | ~new_n9735_ | ~new_n9736_ | ~new_n9739_);
  assign new_n9743_ = ~\all_features[1935]  & (~\all_features[1934]  | (~\all_features[1932]  & ~\all_features[1933]  & ~new_n9739_));
  assign new_n9744_ = \all_features[1935]  & (\all_features[1934]  | (\all_features[1933]  & (\all_features[1932]  | ~new_n9731_ | ~new_n9745_)));
  assign new_n9745_ = ~\all_features[1930]  & ~\all_features[1931] ;
  assign new_n9746_ = \all_features[1935]  & (\all_features[1934]  | (new_n9735_ & (\all_features[1930]  | \all_features[1931]  | \all_features[1929] )));
  assign new_n9747_ = \all_features[1934]  & \all_features[1935]  & (\all_features[1932]  | \all_features[1933]  | new_n9736_ | ~new_n9745_);
  assign new_n9748_ = \all_features[1935]  & (\all_features[1933]  | \all_features[1934]  | \all_features[1932] );
  assign new_n9749_ = new_n9728_ & new_n9737_;
  assign new_n9750_ = ~new_n9751_ & ~new_n9755_;
  assign new_n9751_ = ~new_n9752_ & (\all_features[1931]  | \all_features[1932]  | \all_features[1933]  | \all_features[1934]  | \all_features[1935] );
  assign new_n9752_ = ~new_n9730_ & (new_n9733_ | (~new_n9734_ & (new_n9743_ | (~new_n9738_ & ~new_n9753_))));
  assign new_n9753_ = ~new_n9740_ & (new_n9742_ | (new_n9748_ & (~new_n9744_ | (~new_n9754_ & new_n9746_))));
  assign new_n9754_ = ~\all_features[1933]  & \all_features[1934]  & \all_features[1935]  & (\all_features[1932]  ? new_n9745_ : (new_n9736_ | ~new_n9745_));
  assign new_n9755_ = new_n9729_ & (new_n9734_ | new_n9733_ | (~new_n9738_ & ~new_n9743_ & ~new_n9756_));
  assign new_n9756_ = ~new_n9742_ & ~new_n9740_ & (~new_n9748_ | ~new_n9744_ | new_n9757_);
  assign new_n9757_ = new_n9746_ & new_n9747_ & (new_n9758_ | ~\all_features[1933]  | ~\all_features[1934]  | ~\all_features[1935] );
  assign new_n9758_ = ~\all_features[1931]  & ~\all_features[1932]  & (~\all_features[1930]  | new_n9731_);
  assign new_n9759_ = ~new_n9760_ & ~new_n7407_;
  assign new_n9760_ = new_n7375_ & new_n7405_;
  assign new_n9761_ = new_n9762_ & new_n9789_;
  assign new_n9762_ = ~new_n9763_ & ~new_n9787_;
  assign new_n9763_ = new_n9781_ & ~new_n9786_ & ~new_n9764_ & ~new_n9785_;
  assign new_n9764_ = ~new_n9779_ & ~new_n9780_ & new_n9774_ & (~new_n9768_ | ~new_n9765_);
  assign new_n9765_ = \all_features[4839]  & (\all_features[4838]  | new_n9766_);
  assign new_n9766_ = \all_features[4837]  & (\all_features[4834]  | \all_features[4835]  | \all_features[4836]  | ~new_n9767_);
  assign new_n9767_ = ~\all_features[4832]  & ~\all_features[4833] ;
  assign new_n9768_ = new_n9773_ & new_n9769_ & new_n9771_;
  assign new_n9769_ = \all_features[4839]  & (\all_features[4838]  | (new_n9770_ & (\all_features[4834]  | \all_features[4835]  | \all_features[4833] )));
  assign new_n9770_ = \all_features[4836]  & \all_features[4837] ;
  assign new_n9771_ = \all_features[4839]  & ~new_n9772_ & \all_features[4838] ;
  assign new_n9772_ = ~\all_features[4834]  & ~\all_features[4835]  & ~\all_features[4836]  & ~\all_features[4837]  & (~\all_features[4833]  | ~\all_features[4832] );
  assign new_n9773_ = \all_features[4839]  & (\all_features[4837]  | \all_features[4838]  | \all_features[4836] );
  assign new_n9774_ = ~new_n9775_ & ~new_n9777_;
  assign new_n9775_ = ~new_n9776_ & ~\all_features[4839] ;
  assign new_n9776_ = \all_features[4837]  & \all_features[4838]  & (\all_features[4836]  | (\all_features[4834]  & \all_features[4835]  & \all_features[4833] ));
  assign new_n9777_ = ~\all_features[4839]  & (~\all_features[4838]  | (~\all_features[4836]  & ~\all_features[4837]  & ~new_n9778_));
  assign new_n9778_ = \all_features[4834]  & \all_features[4835] ;
  assign new_n9779_ = ~\all_features[4839]  & (~\all_features[4838]  | (~\all_features[4837]  & (new_n9767_ | ~new_n9778_ | ~\all_features[4836] )));
  assign new_n9780_ = ~\all_features[4839]  & (~new_n9778_ | ~\all_features[4832]  | ~\all_features[4833]  | ~\all_features[4838]  | ~new_n9770_);
  assign new_n9781_ = ~new_n9782_ & ~new_n9784_;
  assign new_n9782_ = ~\all_features[4837]  & new_n9783_ & ((~\all_features[4834]  & new_n9767_) | ~\all_features[4836]  | ~\all_features[4835] );
  assign new_n9783_ = ~\all_features[4838]  & ~\all_features[4839] ;
  assign new_n9784_ = ~\all_features[4839]  & ~\all_features[4838]  & ~\all_features[4837]  & ~\all_features[4835]  & ~\all_features[4836] ;
  assign new_n9785_ = new_n9783_ & (~\all_features[4837]  | (~\all_features[4836]  & (~\all_features[4835]  | (~\all_features[4834]  & ~\all_features[4833] ))));
  assign new_n9786_ = new_n9783_ & (~new_n9770_ | ~\all_features[4835]  | (~\all_features[4834]  & (~\all_features[4832]  | ~\all_features[4833] )));
  assign new_n9787_ = new_n9781_ & new_n9774_ & new_n9788_ & ~new_n9779_ & ~new_n9780_;
  assign new_n9788_ = ~new_n9785_ & ~new_n9786_;
  assign new_n9789_ = ~new_n9790_ & (new_n9784_ | (~new_n9794_ & ~new_n9782_));
  assign new_n9790_ = new_n9781_ & (~new_n9788_ | (~new_n9791_ & ~new_n9777_ & ~new_n9779_));
  assign new_n9791_ = ~new_n9780_ & ~new_n9775_ & (~new_n9773_ | new_n9792_ | ~new_n9765_);
  assign new_n9792_ = ~new_n9772_ & new_n9769_ & \all_features[4838]  & \all_features[4839]  & (~\all_features[4837]  | new_n9793_);
  assign new_n9793_ = ~\all_features[4835]  & ~\all_features[4836]  & (~\all_features[4834]  | new_n9767_);
  assign new_n9794_ = ~new_n9785_ & (new_n9786_ | (~new_n9777_ & (new_n9779_ | (~new_n9775_ & ~new_n9795_))));
  assign new_n9795_ = ~new_n9780_ & (~new_n9773_ | (new_n9765_ & (~new_n9769_ | (~new_n9796_ & new_n9771_))));
  assign new_n9796_ = \all_features[4838]  & \all_features[4839]  & (\all_features[4837]  | (\all_features[4836]  & (\all_features[4835]  | \all_features[4834] )));
  assign new_n9797_ = new_n9830_ & ~new_n9798_ & new_n9827_;
  assign new_n9798_ = ~new_n9799_ & ~new_n9823_;
  assign new_n9799_ = new_n9820_ & (~new_n9814_ | (~new_n9800_ & ~new_n9818_ & ~new_n9822_));
  assign new_n9800_ = ~new_n9811_ & ~new_n9810_ & (~new_n9813_ | ~new_n9809_ | new_n9801_);
  assign new_n9801_ = new_n9802_ & new_n9804_ & (new_n9807_ | ~\all_features[4525]  | ~\all_features[4526]  | ~\all_features[4527] );
  assign new_n9802_ = \all_features[4527]  & (\all_features[4526]  | (new_n9803_ & (\all_features[4522]  | \all_features[4523]  | \all_features[4521] )));
  assign new_n9803_ = \all_features[4524]  & \all_features[4525] ;
  assign new_n9804_ = \all_features[4526]  & \all_features[4527]  & (\all_features[4524]  | \all_features[4525]  | new_n9805_ | ~new_n9806_);
  assign new_n9805_ = \all_features[4520]  & \all_features[4521] ;
  assign new_n9806_ = ~\all_features[4522]  & ~\all_features[4523] ;
  assign new_n9807_ = ~\all_features[4523]  & ~\all_features[4524]  & (~\all_features[4522]  | new_n9808_);
  assign new_n9808_ = ~\all_features[4520]  & ~\all_features[4521] ;
  assign new_n9809_ = \all_features[4527]  & (\all_features[4526]  | (\all_features[4525]  & (\all_features[4524]  | ~new_n9808_ | ~new_n9806_)));
  assign new_n9810_ = ~\all_features[4527]  & (~new_n9803_ | ~\all_features[4522]  | ~\all_features[4523]  | ~\all_features[4526]  | ~new_n9805_);
  assign new_n9811_ = ~new_n9812_ & ~\all_features[4527] ;
  assign new_n9812_ = \all_features[4525]  & \all_features[4526]  & (\all_features[4524]  | (\all_features[4522]  & \all_features[4523]  & \all_features[4521] ));
  assign new_n9813_ = \all_features[4527]  & (\all_features[4525]  | \all_features[4526]  | \all_features[4524] );
  assign new_n9814_ = ~new_n9815_ & ~new_n9817_;
  assign new_n9815_ = new_n9816_ & (~\all_features[4523]  | ~new_n9803_ | (~\all_features[4522]  & ~new_n9805_));
  assign new_n9816_ = ~\all_features[4526]  & ~\all_features[4527] ;
  assign new_n9817_ = new_n9816_ & (~\all_features[4525]  | (~\all_features[4524]  & (~\all_features[4523]  | (~\all_features[4522]  & ~\all_features[4521] ))));
  assign new_n9818_ = ~\all_features[4527]  & (~\all_features[4526]  | new_n9819_);
  assign new_n9819_ = ~\all_features[4525]  & (new_n9808_ | ~\all_features[4523]  | ~\all_features[4524]  | ~\all_features[4522] );
  assign new_n9820_ = ~new_n9821_ & (\all_features[4523]  | \all_features[4524]  | \all_features[4525]  | \all_features[4526]  | \all_features[4527] );
  assign new_n9821_ = ~\all_features[4525]  & new_n9816_ & ((~\all_features[4522]  & new_n9808_) | ~\all_features[4524]  | ~\all_features[4523] );
  assign new_n9822_ = ~\all_features[4527]  & (~\all_features[4526]  | (~\all_features[4525]  & ~\all_features[4524]  & (~\all_features[4523]  | ~\all_features[4522] )));
  assign new_n9823_ = ~new_n9824_ & (\all_features[4523]  | \all_features[4524]  | \all_features[4525]  | \all_features[4526]  | \all_features[4527] );
  assign new_n9824_ = ~new_n9821_ & (new_n9817_ | (~new_n9815_ & (new_n9822_ | (~new_n9818_ & ~new_n9825_))));
  assign new_n9825_ = ~new_n9811_ & (new_n9810_ | (new_n9813_ & (~new_n9809_ | (~new_n9826_ & new_n9802_))));
  assign new_n9826_ = ~\all_features[4525]  & \all_features[4526]  & \all_features[4527]  & (\all_features[4524]  ? new_n9806_ : (new_n9805_ | ~new_n9806_));
  assign new_n9827_ = new_n9814_ & new_n9829_ & new_n9828_ & ~new_n9818_ & ~new_n9821_;
  assign new_n9828_ = ~new_n9810_ & (\all_features[4523]  | \all_features[4524]  | \all_features[4525]  | \all_features[4526]  | \all_features[4527] );
  assign new_n9829_ = ~new_n9811_ & ~new_n9822_;
  assign new_n9830_ = new_n9814_ & new_n9820_ & (new_n9818_ | new_n9831_ | new_n9810_ | ~new_n9829_);
  assign new_n9831_ = new_n9813_ & new_n9809_ & new_n9802_ & new_n9804_;
  assign new_n9832_ = (~new_n9652_ | new_n9833_ | new_n9689_) & (new_n9869_ | new_n9870_ | new_n9893_ | ~new_n9689_);
  assign new_n9833_ = new_n9834_ & new_n9867_;
  assign new_n9834_ = new_n9835_ & new_n9864_;
  assign new_n9835_ = new_n9836_ & new_n9860_;
  assign new_n9836_ = new_n9857_ & (~new_n9851_ | (~new_n9837_ & ~new_n9855_ & ~new_n9859_));
  assign new_n9837_ = ~new_n9846_ & ~new_n9847_ & (~new_n9850_ | ~new_n9849_ | new_n9838_);
  assign new_n9838_ = new_n9839_ & new_n9841_ & (new_n9844_ | ~\all_features[3949]  | ~\all_features[3950]  | ~\all_features[3951] );
  assign new_n9839_ = \all_features[3951]  & (\all_features[3950]  | (new_n9840_ & (\all_features[3946]  | \all_features[3947]  | \all_features[3945] )));
  assign new_n9840_ = \all_features[3948]  & \all_features[3949] ;
  assign new_n9841_ = \all_features[3950]  & \all_features[3951]  & (\all_features[3948]  | \all_features[3949]  | new_n9842_ | ~new_n9843_);
  assign new_n9842_ = \all_features[3944]  & \all_features[3945] ;
  assign new_n9843_ = ~\all_features[3946]  & ~\all_features[3947] ;
  assign new_n9844_ = ~\all_features[3947]  & ~\all_features[3948]  & (~\all_features[3946]  | new_n9845_);
  assign new_n9845_ = ~\all_features[3944]  & ~\all_features[3945] ;
  assign new_n9846_ = ~\all_features[3951]  & (~new_n9840_ | ~\all_features[3946]  | ~\all_features[3947]  | ~\all_features[3950]  | ~new_n9842_);
  assign new_n9847_ = ~new_n9848_ & ~\all_features[3951] ;
  assign new_n9848_ = \all_features[3949]  & \all_features[3950]  & (\all_features[3948]  | (\all_features[3946]  & \all_features[3947]  & \all_features[3945] ));
  assign new_n9849_ = \all_features[3951]  & (\all_features[3950]  | (\all_features[3949]  & (\all_features[3948]  | ~new_n9843_ | ~new_n9845_)));
  assign new_n9850_ = \all_features[3951]  & (\all_features[3949]  | \all_features[3950]  | \all_features[3948] );
  assign new_n9851_ = ~new_n9852_ & ~new_n9854_;
  assign new_n9852_ = new_n9853_ & (~\all_features[3947]  | ~new_n9840_ | (~\all_features[3946]  & ~new_n9842_));
  assign new_n9853_ = ~\all_features[3950]  & ~\all_features[3951] ;
  assign new_n9854_ = new_n9853_ & (~\all_features[3949]  | (~\all_features[3948]  & (~\all_features[3947]  | (~\all_features[3946]  & ~\all_features[3945] ))));
  assign new_n9855_ = ~\all_features[3951]  & (~\all_features[3950]  | new_n9856_);
  assign new_n9856_ = ~\all_features[3949]  & (new_n9845_ | ~\all_features[3947]  | ~\all_features[3948]  | ~\all_features[3946] );
  assign new_n9857_ = ~new_n9858_ & (\all_features[3947]  | \all_features[3948]  | \all_features[3949]  | \all_features[3950]  | \all_features[3951] );
  assign new_n9858_ = ~\all_features[3949]  & new_n9853_ & ((~\all_features[3946]  & new_n9845_) | ~\all_features[3948]  | ~\all_features[3947] );
  assign new_n9859_ = ~\all_features[3951]  & (~\all_features[3950]  | (~\all_features[3949]  & ~\all_features[3948]  & (~\all_features[3947]  | ~\all_features[3946] )));
  assign new_n9860_ = ~new_n9861_ & (\all_features[3947]  | \all_features[3948]  | \all_features[3949]  | \all_features[3950]  | \all_features[3951] );
  assign new_n9861_ = ~new_n9858_ & (new_n9854_ | (~new_n9852_ & (new_n9859_ | (~new_n9855_ & ~new_n9862_))));
  assign new_n9862_ = ~new_n9847_ & (new_n9846_ | (new_n9850_ & (~new_n9849_ | (~new_n9863_ & new_n9839_))));
  assign new_n9863_ = ~\all_features[3949]  & \all_features[3950]  & \all_features[3951]  & (\all_features[3948]  ? new_n9843_ : (new_n9842_ | ~new_n9843_));
  assign new_n9864_ = new_n9851_ & new_n9857_ & (new_n9855_ | new_n9866_ | new_n9846_ | ~new_n9865_);
  assign new_n9865_ = ~new_n9847_ & ~new_n9859_;
  assign new_n9866_ = new_n9850_ & new_n9849_ & new_n9839_ & new_n9841_;
  assign new_n9867_ = new_n9868_ & new_n9865_ & new_n9851_ & ~new_n9855_ & ~new_n9858_;
  assign new_n9868_ = ~new_n9846_ & (\all_features[3947]  | \all_features[3948]  | \all_features[3949]  | \all_features[3950]  | \all_features[3951] );
  assign new_n9869_ = ~new_n6806_ & new_n6837_;
  assign new_n9870_ = ~new_n9892_ & ~new_n9891_ & ~new_n9890_ & ~new_n9871_ & ~new_n9888_;
  assign new_n9871_ = ~new_n9872_ & ~new_n9886_ & new_n9875_ & (~new_n9887_ | ~new_n9879_);
  assign new_n9872_ = ~\all_features[4183]  & (~\all_features[4182]  | new_n9873_);
  assign new_n9873_ = ~\all_features[4181]  & (new_n9874_ | ~\all_features[4179]  | ~\all_features[4180]  | ~\all_features[4178] );
  assign new_n9874_ = ~\all_features[4176]  & ~\all_features[4177] ;
  assign new_n9875_ = ~new_n9876_ & ~new_n9878_;
  assign new_n9876_ = ~new_n9877_ & ~\all_features[4183] ;
  assign new_n9877_ = \all_features[4181]  & \all_features[4182]  & (\all_features[4180]  | (\all_features[4178]  & \all_features[4179]  & \all_features[4177] ));
  assign new_n9878_ = ~\all_features[4183]  & (~\all_features[4182]  | (~\all_features[4181]  & ~\all_features[4180]  & (~\all_features[4179]  | ~\all_features[4178] )));
  assign new_n9879_ = new_n9885_ & new_n9880_ & new_n9882_;
  assign new_n9880_ = \all_features[4183]  & (\all_features[4182]  | (new_n9881_ & (\all_features[4178]  | \all_features[4179]  | \all_features[4177] )));
  assign new_n9881_ = \all_features[4180]  & \all_features[4181] ;
  assign new_n9882_ = \all_features[4182]  & \all_features[4183]  & (\all_features[4180]  | \all_features[4181]  | new_n9883_ | ~new_n9884_);
  assign new_n9883_ = \all_features[4176]  & \all_features[4177] ;
  assign new_n9884_ = ~\all_features[4178]  & ~\all_features[4179] ;
  assign new_n9885_ = \all_features[4183]  & (\all_features[4181]  | \all_features[4182]  | \all_features[4180] );
  assign new_n9886_ = ~\all_features[4183]  & (~new_n9881_ | ~\all_features[4178]  | ~\all_features[4179]  | ~\all_features[4182]  | ~new_n9883_);
  assign new_n9887_ = \all_features[4183]  & (\all_features[4182]  | (\all_features[4181]  & (\all_features[4180]  | ~new_n9884_ | ~new_n9874_)));
  assign new_n9888_ = new_n9889_ & (~\all_features[4179]  | ~new_n9881_ | (~\all_features[4178]  & ~new_n9883_));
  assign new_n9889_ = ~\all_features[4182]  & ~\all_features[4183] ;
  assign new_n9890_ = new_n9889_ & (~\all_features[4181]  | (~\all_features[4180]  & (~\all_features[4179]  | (~\all_features[4178]  & ~\all_features[4177] ))));
  assign new_n9891_ = ~\all_features[4181]  & new_n9889_ & ((~\all_features[4178]  & new_n9874_) | ~\all_features[4180]  | ~\all_features[4179] );
  assign new_n9892_ = ~\all_features[4183]  & ~\all_features[4182]  & ~\all_features[4181]  & ~\all_features[4179]  & ~\all_features[4180] ;
  assign new_n9893_ = new_n9894_ & new_n9875_ & ~new_n9892_ & ~new_n9886_ & ~new_n9872_ & ~new_n9891_;
  assign new_n9894_ = ~new_n9888_ & ~new_n9890_;
  assign new_n9895_ = new_n9997_ & (new_n9998_ ? (~new_n10000_ | (new_n7603_ & new_n7625_)) : new_n9896_);
  assign new_n9896_ = (~new_n9966_ | ~new_n9897_ | (new_n9634_ & (new_n9996_ | new_n9612_))) & (~new_n9933_ | new_n9897_);
  assign new_n9897_ = new_n9932_ & (new_n9930_ | new_n9898_);
  assign new_n9898_ = new_n9899_ & (new_n9913_ | new_n9926_);
  assign new_n9899_ = new_n9900_ & (\all_features[3955]  | \all_features[3956]  | \all_features[3957]  | \all_features[3958]  | \all_features[3959] );
  assign new_n9900_ = new_n9912_ & (~new_n9915_ | (new_n9923_ & (~new_n9918_ | new_n9901_)));
  assign new_n9901_ = new_n9911_ & ~new_n9905_ & new_n9902_;
  assign new_n9902_ = \all_features[3959]  & (\all_features[3958]  | new_n9903_);
  assign new_n9903_ = \all_features[3957]  & (\all_features[3954]  | \all_features[3955]  | \all_features[3956]  | ~new_n9904_);
  assign new_n9904_ = ~\all_features[3952]  & ~\all_features[3953] ;
  assign new_n9905_ = ~new_n9908_ & new_n9906_ & \all_features[3958]  & \all_features[3959]  & (~\all_features[3957]  | new_n9910_);
  assign new_n9906_ = \all_features[3959]  & (\all_features[3958]  | (new_n9907_ & (\all_features[3954]  | \all_features[3955]  | \all_features[3953] )));
  assign new_n9907_ = \all_features[3956]  & \all_features[3957] ;
  assign new_n9908_ = ~\all_features[3957]  & ~\all_features[3956]  & ~\all_features[3955]  & ~new_n9909_ & ~\all_features[3954] ;
  assign new_n9909_ = \all_features[3952]  & \all_features[3953] ;
  assign new_n9910_ = ~\all_features[3955]  & ~\all_features[3956]  & (~\all_features[3954]  | new_n9904_);
  assign new_n9911_ = \all_features[3959]  & (\all_features[3957]  | \all_features[3958]  | \all_features[3956] );
  assign new_n9912_ = ~new_n9913_ & (\all_features[3955]  | \all_features[3956]  | \all_features[3957]  | \all_features[3958]  | \all_features[3959] );
  assign new_n9913_ = ~\all_features[3957]  & new_n9914_ & ((~\all_features[3954]  & new_n9904_) | ~\all_features[3956]  | ~\all_features[3955] );
  assign new_n9914_ = ~\all_features[3958]  & ~\all_features[3959] ;
  assign new_n9915_ = ~new_n9916_ & ~new_n9917_;
  assign new_n9916_ = new_n9914_ & (~\all_features[3957]  | (~\all_features[3956]  & (~\all_features[3955]  | (~\all_features[3954]  & ~\all_features[3953] ))));
  assign new_n9917_ = new_n9914_ & (~\all_features[3955]  | ~new_n9907_ | (~\all_features[3954]  & ~new_n9909_));
  assign new_n9918_ = ~new_n9919_ & ~new_n9921_;
  assign new_n9919_ = ~new_n9920_ & ~\all_features[3959] ;
  assign new_n9920_ = \all_features[3957]  & \all_features[3958]  & (\all_features[3956]  | (\all_features[3954]  & \all_features[3955]  & \all_features[3953] ));
  assign new_n9921_ = ~\all_features[3959]  & (~\all_features[3958]  | ~new_n9909_ | ~new_n9907_ | ~new_n9922_);
  assign new_n9922_ = \all_features[3954]  & \all_features[3955] ;
  assign new_n9923_ = ~new_n9924_ & ~new_n9925_;
  assign new_n9924_ = ~\all_features[3959]  & (~\all_features[3958]  | (~\all_features[3956]  & ~\all_features[3957]  & ~new_n9922_));
  assign new_n9925_ = ~\all_features[3959]  & (~\all_features[3958]  | (~\all_features[3957]  & (new_n9904_ | ~new_n9922_ | ~\all_features[3956] )));
  assign new_n9926_ = ~new_n9916_ & (new_n9917_ | (~new_n9924_ & (new_n9925_ | (~new_n9927_ & ~new_n9919_))));
  assign new_n9927_ = ~new_n9921_ & (~new_n9911_ | (new_n9902_ & (~new_n9906_ | (~new_n9929_ & new_n9928_))));
  assign new_n9928_ = \all_features[3959]  & ~new_n9908_ & \all_features[3958] ;
  assign new_n9929_ = \all_features[3958]  & \all_features[3959]  & (\all_features[3957]  | (\all_features[3956]  & (\all_features[3955]  | \all_features[3954] )));
  assign new_n9930_ = new_n9915_ & new_n9912_ & (~new_n9923_ | ~new_n9918_ | (new_n9902_ & new_n9931_));
  assign new_n9931_ = new_n9911_ & new_n9928_ & new_n9906_;
  assign new_n9932_ = new_n9915_ & new_n9912_ & ~new_n9925_ & ~new_n9924_ & ~new_n9919_ & ~new_n9921_;
  assign new_n9933_ = new_n9936_ & new_n9934_ & (new_n9958_ | (~new_n9963_ & ~new_n9959_));
  assign new_n9934_ = ~new_n9935_ & ~new_n9932_;
  assign new_n9935_ = new_n9930_ & new_n9900_;
  assign new_n9936_ = new_n9959_ | ((new_n9958_ | (~new_n9937_ & ~new_n9961_ & ~new_n9962_)) & (new_n9958_ | new_n9961_ | new_n9962_));
  assign new_n9937_ = ~new_n9949_ & ~new_n9951_ & (new_n9954_ | new_n9952_ | new_n9938_);
  assign new_n9938_ = new_n9948_ & ~new_n9942_ & new_n9939_;
  assign new_n9939_ = \all_features[3975]  & (\all_features[3974]  | new_n9940_);
  assign new_n9940_ = \all_features[3973]  & (\all_features[3970]  | \all_features[3971]  | \all_features[3972]  | ~new_n9941_);
  assign new_n9941_ = ~\all_features[3968]  & ~\all_features[3969] ;
  assign new_n9942_ = ~new_n9945_ & new_n9943_ & \all_features[3974]  & \all_features[3975]  & (~\all_features[3973]  | new_n9947_);
  assign new_n9943_ = \all_features[3975]  & (\all_features[3974]  | (new_n9944_ & (\all_features[3970]  | \all_features[3971]  | \all_features[3969] )));
  assign new_n9944_ = \all_features[3972]  & \all_features[3973] ;
  assign new_n9945_ = ~\all_features[3973]  & ~\all_features[3972]  & ~\all_features[3971]  & ~new_n9946_ & ~\all_features[3970] ;
  assign new_n9946_ = \all_features[3968]  & \all_features[3969] ;
  assign new_n9947_ = ~\all_features[3971]  & ~\all_features[3972]  & (~\all_features[3970]  | new_n9941_);
  assign new_n9948_ = \all_features[3975]  & (\all_features[3973]  | \all_features[3974]  | \all_features[3972] );
  assign new_n9949_ = ~\all_features[3975]  & (~\all_features[3974]  | (~\all_features[3972]  & ~\all_features[3973]  & ~new_n9950_));
  assign new_n9950_ = \all_features[3970]  & \all_features[3971] ;
  assign new_n9951_ = ~\all_features[3975]  & (~\all_features[3974]  | (~\all_features[3973]  & (new_n9941_ | ~new_n9950_ | ~\all_features[3972] )));
  assign new_n9952_ = ~new_n9953_ & ~\all_features[3975] ;
  assign new_n9953_ = \all_features[3973]  & \all_features[3974]  & (\all_features[3972]  | (\all_features[3970]  & \all_features[3971]  & \all_features[3969] ));
  assign new_n9954_ = ~\all_features[3975]  & (~\all_features[3974]  | ~new_n9946_ | ~new_n9944_ | ~new_n9950_);
  assign new_n9956_ = \all_features[3975]  & ~new_n9945_ & \all_features[3974] ;
  assign new_n9958_ = ~\all_features[3975]  & ~\all_features[3974]  & ~\all_features[3973]  & ~\all_features[3971]  & ~\all_features[3972] ;
  assign new_n9959_ = ~\all_features[3973]  & new_n9960_ & ((~\all_features[3970]  & new_n9941_) | ~\all_features[3972]  | ~\all_features[3971] );
  assign new_n9960_ = ~\all_features[3974]  & ~\all_features[3975] ;
  assign new_n9961_ = new_n9960_ & (~\all_features[3973]  | (~\all_features[3972]  & (~\all_features[3971]  | (~\all_features[3970]  & ~\all_features[3969] ))));
  assign new_n9962_ = new_n9960_ & (~\all_features[3971]  | ~new_n9944_ | (~\all_features[3970]  & ~new_n9946_));
  assign new_n9963_ = ~new_n9961_ & (new_n9962_ | (~new_n9949_ & (new_n9951_ | (~new_n9964_ & ~new_n9952_))));
  assign new_n9964_ = ~new_n9954_ & (~new_n9948_ | (new_n9939_ & (~new_n9943_ | (~new_n9965_ & new_n9956_))));
  assign new_n9965_ = \all_features[3974]  & \all_features[3975]  & (\all_features[3973]  | (\all_features[3972]  & (\all_features[3971]  | \all_features[3970] )));
  assign new_n9966_ = ~new_n9995_ & new_n9967_;
  assign new_n9967_ = ~new_n9968_ & ~new_n9993_;
  assign new_n9968_ = new_n9969_ & (~new_n9987_ | (new_n9983_ & (new_n9975_ | new_n9990_ | new_n9992_)));
  assign new_n9969_ = ~new_n9970_ & ~new_n9974_;
  assign new_n9970_ = new_n9971_ & ((~\all_features[2986]  & new_n9973_) | ~\all_features[2988]  | ~\all_features[2987] );
  assign new_n9971_ = ~\all_features[2989]  & new_n9972_;
  assign new_n9972_ = ~\all_features[2990]  & ~\all_features[2991] ;
  assign new_n9973_ = ~\all_features[2984]  & ~\all_features[2985] ;
  assign new_n9974_ = new_n9971_ & ~\all_features[2987]  & ~\all_features[2988] ;
  assign new_n9975_ = new_n9976_ & (~new_n9978_ | (~new_n9982_ & \all_features[2989]  & \all_features[2990]  & \all_features[2991] ));
  assign new_n9976_ = \all_features[2991]  & (\all_features[2990]  | (~new_n9977_ & \all_features[2989] ));
  assign new_n9977_ = new_n9973_ & ~\all_features[2988]  & ~\all_features[2986]  & ~\all_features[2987] ;
  assign new_n9978_ = \all_features[2991]  & \all_features[2990]  & ~new_n9981_ & new_n9979_;
  assign new_n9979_ = \all_features[2991]  & (\all_features[2990]  | (new_n9980_ & (\all_features[2986]  | \all_features[2987]  | \all_features[2985] )));
  assign new_n9980_ = \all_features[2988]  & \all_features[2989] ;
  assign new_n9981_ = ~\all_features[2986]  & ~\all_features[2987]  & ~\all_features[2988]  & ~\all_features[2989]  & (~\all_features[2985]  | ~\all_features[2984] );
  assign new_n9982_ = ~\all_features[2987]  & ~\all_features[2988]  & (~\all_features[2986]  | new_n9973_);
  assign new_n9983_ = ~new_n9984_ & ~new_n9986_;
  assign new_n9984_ = ~\all_features[2991]  & (~\all_features[2990]  | (~\all_features[2988]  & ~\all_features[2989]  & ~new_n9985_));
  assign new_n9985_ = \all_features[2986]  & \all_features[2987] ;
  assign new_n9986_ = ~\all_features[2991]  & (~\all_features[2990]  | (~\all_features[2989]  & (new_n9973_ | ~\all_features[2988]  | ~new_n9985_)));
  assign new_n9987_ = ~new_n9988_ & ~new_n9989_;
  assign new_n9988_ = new_n9972_ & (~new_n9980_ | ~\all_features[2987]  | (~\all_features[2986]  & (~\all_features[2984]  | ~\all_features[2985] )));
  assign new_n9989_ = new_n9972_ & (~\all_features[2989]  | (~\all_features[2988]  & (~\all_features[2987]  | (~\all_features[2986]  & ~\all_features[2985] ))));
  assign new_n9990_ = ~new_n9991_ & ~\all_features[2991] ;
  assign new_n9991_ = \all_features[2989]  & \all_features[2990]  & (\all_features[2988]  | (\all_features[2986]  & \all_features[2987]  & \all_features[2985] ));
  assign new_n9992_ = ~\all_features[2991]  & (~new_n9980_ | ~\all_features[2984]  | ~\all_features[2985]  | ~\all_features[2990]  | ~new_n9985_);
  assign new_n9993_ = new_n9987_ & ~new_n9994_ & new_n9969_;
  assign new_n9994_ = ~new_n9984_ & ~new_n9986_ & ~new_n9990_ & ~new_n9992_ & (~new_n9978_ | ~new_n9976_);
  assign new_n9995_ = new_n9987_ & new_n9983_ & ~new_n9992_ & ~new_n9990_ & ~new_n9970_ & ~new_n9974_;
  assign new_n9996_ = new_n9636_ & new_n9640_;
  assign new_n9997_ = (new_n10036_ | new_n10000_ | ~new_n9998_) & (new_n9934_ | new_n9897_ | new_n10128_ | new_n9998_);
  assign new_n9998_ = new_n7479_ & new_n9999_;
  assign new_n9999_ = new_n7510_ & new_n7513_;
  assign new_n10000_ = new_n10001_ & new_n10027_;
  assign new_n10001_ = ~new_n10002_ & ~new_n10024_;
  assign new_n10002_ = ~new_n10023_ & ~new_n10022_ & ~new_n10021_ & ~new_n10003_ & ~new_n10019_;
  assign new_n10003_ = new_n10004_ & (~new_n10017_ | ~new_n10018_ | ~new_n10014_ | ~new_n10016_);
  assign new_n10004_ = ~new_n10011_ & ~new_n10010_ & ~new_n10005_ & ~new_n10008_;
  assign new_n10005_ = ~\all_features[3711]  & (~\all_features[3710]  | (~\all_features[3709]  & (new_n10006_ | ~new_n10007_ | ~\all_features[3708] )));
  assign new_n10006_ = ~\all_features[3704]  & ~\all_features[3705] ;
  assign new_n10007_ = \all_features[3706]  & \all_features[3707] ;
  assign new_n10008_ = ~new_n10009_ & ~\all_features[3711] ;
  assign new_n10009_ = \all_features[3709]  & \all_features[3710]  & (\all_features[3708]  | (\all_features[3706]  & \all_features[3707]  & \all_features[3705] ));
  assign new_n10010_ = ~\all_features[3711]  & (~\all_features[3710]  | (~\all_features[3708]  & ~\all_features[3709]  & ~new_n10007_));
  assign new_n10011_ = ~\all_features[3711]  & (~\all_features[3710]  | ~new_n10012_ | ~new_n10013_ | ~new_n10007_);
  assign new_n10012_ = \all_features[3708]  & \all_features[3709] ;
  assign new_n10013_ = \all_features[3704]  & \all_features[3705] ;
  assign new_n10014_ = \all_features[3711]  & (\all_features[3710]  | (\all_features[3709]  & (\all_features[3708]  | ~new_n10006_ | ~new_n10015_)));
  assign new_n10015_ = ~\all_features[3706]  & ~\all_features[3707] ;
  assign new_n10016_ = \all_features[3711]  & (\all_features[3710]  | (new_n10012_ & (\all_features[3706]  | \all_features[3707]  | \all_features[3705] )));
  assign new_n10017_ = \all_features[3710]  & \all_features[3711]  & (\all_features[3708]  | \all_features[3709]  | new_n10013_ | ~new_n10015_);
  assign new_n10018_ = \all_features[3711]  & (\all_features[3709]  | \all_features[3710]  | \all_features[3708] );
  assign new_n10019_ = new_n10020_ & (~\all_features[3709]  | (~\all_features[3708]  & (~\all_features[3707]  | (~\all_features[3706]  & ~\all_features[3705] ))));
  assign new_n10020_ = ~\all_features[3710]  & ~\all_features[3711] ;
  assign new_n10021_ = ~\all_features[3709]  & new_n10020_ & ((~\all_features[3706]  & new_n10006_) | ~\all_features[3708]  | ~\all_features[3707] );
  assign new_n10022_ = new_n10020_ & (~\all_features[3707]  | ~new_n10012_ | (~\all_features[3706]  & ~new_n10013_));
  assign new_n10023_ = ~\all_features[3711]  & ~\all_features[3710]  & ~\all_features[3709]  & ~\all_features[3707]  & ~\all_features[3708] ;
  assign new_n10024_ = new_n10026_ & new_n10025_ & ~new_n10021_ & ~new_n10011_ & ~new_n10005_ & ~new_n10008_;
  assign new_n10025_ = ~new_n10010_ & ~new_n10023_;
  assign new_n10026_ = ~new_n10019_ & ~new_n10022_;
  assign new_n10027_ = ~new_n10028_ & ~new_n10032_;
  assign new_n10028_ = ~new_n10029_ & ~new_n10023_;
  assign new_n10029_ = ~new_n10021_ & (new_n10019_ | (~new_n10022_ & (new_n10010_ | (~new_n10005_ & ~new_n10030_))));
  assign new_n10030_ = ~new_n10008_ & (new_n10011_ | (new_n10018_ & (~new_n10014_ | (~new_n10031_ & new_n10016_))));
  assign new_n10031_ = ~\all_features[3709]  & \all_features[3710]  & \all_features[3711]  & (\all_features[3708]  ? new_n10015_ : (new_n10013_ | ~new_n10015_));
  assign new_n10032_ = ~new_n10021_ & ~new_n10023_ & (~new_n10026_ | (~new_n10033_ & ~new_n10005_ & ~new_n10010_));
  assign new_n10033_ = ~new_n10011_ & ~new_n10008_ & (~new_n10018_ | ~new_n10014_ | new_n10034_);
  assign new_n10034_ = new_n10016_ & new_n10017_ & (new_n10035_ | ~\all_features[3709]  | ~\all_features[3710]  | ~\all_features[3711] );
  assign new_n10035_ = ~\all_features[3707]  & ~\all_features[3708]  & (~\all_features[3706]  | new_n10006_);
  assign new_n10036_ = (new_n10071_ & new_n10037_) | (new_n10100_ & new_n10125_ & new_n10127_ & ~new_n10037_);
  assign new_n10037_ = new_n10069_ & new_n10066_ & new_n10038_ & new_n10060_;
  assign new_n10038_ = ~new_n10039_ & ~new_n10059_;
  assign new_n10039_ = ~new_n10053_ & (new_n10055_ | (~new_n10056_ & (new_n10057_ | (~new_n10040_ & ~new_n10058_))));
  assign new_n10040_ = ~new_n10041_ & (new_n10043_ | (new_n10052_ & (~new_n10047_ | (~new_n10051_ & new_n10050_))));
  assign new_n10041_ = ~new_n10042_ & ~\all_features[3319] ;
  assign new_n10042_ = \all_features[3317]  & \all_features[3318]  & (\all_features[3316]  | (\all_features[3314]  & \all_features[3315]  & \all_features[3313] ));
  assign new_n10043_ = ~\all_features[3319]  & (~\all_features[3318]  | ~new_n10044_ | ~new_n10045_ | ~new_n10046_);
  assign new_n10044_ = \all_features[3312]  & \all_features[3313] ;
  assign new_n10045_ = \all_features[3316]  & \all_features[3317] ;
  assign new_n10046_ = \all_features[3314]  & \all_features[3315] ;
  assign new_n10047_ = \all_features[3319]  & (\all_features[3318]  | (\all_features[3317]  & (\all_features[3316]  | ~new_n10049_ | ~new_n10048_)));
  assign new_n10048_ = ~\all_features[3312]  & ~\all_features[3313] ;
  assign new_n10049_ = ~\all_features[3314]  & ~\all_features[3315] ;
  assign new_n10050_ = \all_features[3319]  & (\all_features[3318]  | (new_n10045_ & (\all_features[3314]  | \all_features[3315]  | \all_features[3313] )));
  assign new_n10051_ = ~\all_features[3317]  & \all_features[3318]  & \all_features[3319]  & (\all_features[3316]  ? new_n10049_ : (new_n10044_ | ~new_n10049_));
  assign new_n10052_ = \all_features[3319]  & (\all_features[3317]  | \all_features[3318]  | \all_features[3316] );
  assign new_n10053_ = ~\all_features[3317]  & new_n10054_ & ((~\all_features[3314]  & new_n10048_) | ~\all_features[3316]  | ~\all_features[3315] );
  assign new_n10054_ = ~\all_features[3318]  & ~\all_features[3319] ;
  assign new_n10055_ = new_n10054_ & (~\all_features[3317]  | (~\all_features[3316]  & (~\all_features[3315]  | (~\all_features[3314]  & ~\all_features[3313] ))));
  assign new_n10056_ = new_n10054_ & (~\all_features[3315]  | ~new_n10045_ | (~\all_features[3314]  & ~new_n10044_));
  assign new_n10057_ = ~\all_features[3319]  & (~\all_features[3318]  | (~\all_features[3316]  & ~\all_features[3317]  & ~new_n10046_));
  assign new_n10058_ = ~\all_features[3319]  & (~\all_features[3318]  | (~\all_features[3317]  & (new_n10048_ | ~new_n10046_ | ~\all_features[3316] )));
  assign new_n10059_ = ~\all_features[3319]  & ~\all_features[3318]  & ~\all_features[3317]  & ~\all_features[3315]  & ~\all_features[3316] ;
  assign new_n10060_ = ~new_n10053_ & ~new_n10059_ & (~new_n10065_ | (~new_n10061_ & ~new_n10057_ & ~new_n10058_));
  assign new_n10061_ = ~new_n10041_ & ~new_n10043_ & (~new_n10052_ | ~new_n10047_ | new_n10062_);
  assign new_n10062_ = new_n10050_ & new_n10063_ & (new_n10064_ | ~\all_features[3317]  | ~\all_features[3318]  | ~\all_features[3319] );
  assign new_n10063_ = \all_features[3318]  & \all_features[3319]  & (\all_features[3316]  | \all_features[3317]  | new_n10044_ | ~new_n10049_);
  assign new_n10064_ = ~\all_features[3315]  & ~\all_features[3316]  & (~\all_features[3314]  | new_n10048_);
  assign new_n10065_ = ~new_n10055_ & ~new_n10056_;
  assign new_n10066_ = ~new_n10059_ & ~new_n10056_ & ~new_n10055_ & ~new_n10067_ & ~new_n10053_;
  assign new_n10067_ = new_n10068_ & (~new_n10063_ | ~new_n10052_ | ~new_n10047_ | ~new_n10050_);
  assign new_n10068_ = ~new_n10043_ & ~new_n10041_ & ~new_n10057_ & ~new_n10058_;
  assign new_n10069_ = new_n10070_ & new_n10065_ & ~new_n10041_ & ~new_n10058_ & ~new_n10053_ & ~new_n10057_;
  assign new_n10070_ = ~new_n10043_ & ~new_n10059_;
  assign new_n10071_ = new_n10099_ & new_n10072_ & new_n10097_;
  assign new_n10072_ = new_n10073_ & (~new_n10087_ | (new_n10090_ & (new_n10079_ | new_n10094_ | new_n10095_)));
  assign new_n10073_ = ~new_n10074_ & ~new_n10077_;
  assign new_n10074_ = new_n10075_ & ~\all_features[4539]  & ~\all_features[4540] ;
  assign new_n10075_ = ~\all_features[4541]  & new_n10076_;
  assign new_n10076_ = ~\all_features[4542]  & ~\all_features[4543] ;
  assign new_n10077_ = new_n10075_ & ((~\all_features[4538]  & new_n10078_) | ~\all_features[4540]  | ~\all_features[4539] );
  assign new_n10078_ = ~\all_features[4536]  & ~\all_features[4537] ;
  assign new_n10079_ = new_n10080_ & (~new_n10082_ | (~new_n10086_ & \all_features[4541]  & \all_features[4542]  & \all_features[4543] ));
  assign new_n10080_ = \all_features[4543]  & (\all_features[4542]  | (~new_n10081_ & \all_features[4541] ));
  assign new_n10081_ = new_n10078_ & ~\all_features[4540]  & ~\all_features[4538]  & ~\all_features[4539] ;
  assign new_n10082_ = \all_features[4543]  & \all_features[4542]  & ~new_n10085_ & new_n10083_;
  assign new_n10083_ = \all_features[4543]  & (\all_features[4542]  | (new_n10084_ & (\all_features[4538]  | \all_features[4539]  | \all_features[4537] )));
  assign new_n10084_ = \all_features[4540]  & \all_features[4541] ;
  assign new_n10085_ = ~\all_features[4538]  & ~\all_features[4539]  & ~\all_features[4540]  & ~\all_features[4541]  & (~\all_features[4537]  | ~\all_features[4536] );
  assign new_n10086_ = ~\all_features[4539]  & ~\all_features[4540]  & (~\all_features[4538]  | new_n10078_);
  assign new_n10087_ = ~new_n10088_ & ~new_n10089_;
  assign new_n10088_ = new_n10076_ & (~new_n10084_ | ~\all_features[4539]  | (~\all_features[4538]  & (~\all_features[4536]  | ~\all_features[4537] )));
  assign new_n10089_ = new_n10076_ & (~\all_features[4541]  | (~\all_features[4540]  & (~\all_features[4539]  | (~\all_features[4538]  & ~\all_features[4537] ))));
  assign new_n10090_ = ~new_n10091_ & ~new_n10093_;
  assign new_n10091_ = ~\all_features[4543]  & (~\all_features[4542]  | (~\all_features[4540]  & ~\all_features[4541]  & ~new_n10092_));
  assign new_n10092_ = \all_features[4538]  & \all_features[4539] ;
  assign new_n10093_ = ~\all_features[4543]  & (~\all_features[4542]  | (~\all_features[4541]  & (new_n10078_ | ~new_n10092_ | ~\all_features[4540] )));
  assign new_n10094_ = ~\all_features[4543]  & (~new_n10092_ | ~\all_features[4536]  | ~\all_features[4537]  | ~\all_features[4542]  | ~new_n10084_);
  assign new_n10095_ = ~new_n10096_ & ~\all_features[4543] ;
  assign new_n10096_ = \all_features[4541]  & \all_features[4542]  & (\all_features[4540]  | (\all_features[4538]  & \all_features[4539]  & \all_features[4537] ));
  assign new_n10097_ = new_n10087_ & ~new_n10098_ & new_n10073_;
  assign new_n10098_ = ~new_n10091_ & ~new_n10093_ & ~new_n10094_ & ~new_n10095_ & (~new_n10082_ | ~new_n10080_);
  assign new_n10099_ = new_n10090_ & new_n10087_ & ~new_n10095_ & ~new_n10094_ & ~new_n10074_ & ~new_n10077_;
  assign new_n10100_ = new_n10101_ & (~new_n10115_ | (new_n10118_ & (new_n10107_ | new_n10122_ | new_n10123_)));
  assign new_n10101_ = ~new_n10102_ & ~new_n10105_;
  assign new_n10102_ = new_n10103_ & ~\all_features[1027]  & ~\all_features[1028] ;
  assign new_n10103_ = ~\all_features[1029]  & new_n10104_;
  assign new_n10104_ = ~\all_features[1030]  & ~\all_features[1031] ;
  assign new_n10105_ = new_n10103_ & ((~\all_features[1026]  & new_n10106_) | ~\all_features[1028]  | ~\all_features[1027] );
  assign new_n10106_ = ~\all_features[1024]  & ~\all_features[1025] ;
  assign new_n10107_ = new_n10108_ & (~new_n10110_ | (~new_n10114_ & \all_features[1029]  & \all_features[1030]  & \all_features[1031] ));
  assign new_n10108_ = \all_features[1031]  & (\all_features[1030]  | (~new_n10109_ & \all_features[1029] ));
  assign new_n10109_ = new_n10106_ & ~\all_features[1028]  & ~\all_features[1026]  & ~\all_features[1027] ;
  assign new_n10110_ = \all_features[1031]  & \all_features[1030]  & ~new_n10113_ & new_n10111_;
  assign new_n10111_ = \all_features[1031]  & (\all_features[1030]  | (new_n10112_ & (\all_features[1026]  | \all_features[1027]  | \all_features[1025] )));
  assign new_n10112_ = \all_features[1028]  & \all_features[1029] ;
  assign new_n10113_ = ~\all_features[1026]  & ~\all_features[1027]  & ~\all_features[1028]  & ~\all_features[1029]  & (~\all_features[1025]  | ~\all_features[1024] );
  assign new_n10114_ = ~\all_features[1027]  & ~\all_features[1028]  & (~\all_features[1026]  | new_n10106_);
  assign new_n10115_ = ~new_n10116_ & ~new_n10117_;
  assign new_n10116_ = new_n10104_ & (~new_n10112_ | ~\all_features[1027]  | (~\all_features[1026]  & (~\all_features[1024]  | ~\all_features[1025] )));
  assign new_n10117_ = new_n10104_ & (~\all_features[1029]  | (~\all_features[1028]  & (~\all_features[1027]  | (~\all_features[1026]  & ~\all_features[1025] ))));
  assign new_n10118_ = ~new_n10119_ & ~new_n10121_;
  assign new_n10119_ = ~\all_features[1031]  & (~\all_features[1030]  | (~\all_features[1028]  & ~\all_features[1029]  & ~new_n10120_));
  assign new_n10120_ = \all_features[1026]  & \all_features[1027] ;
  assign new_n10121_ = ~\all_features[1031]  & (~\all_features[1030]  | (~\all_features[1029]  & (new_n10106_ | ~new_n10120_ | ~\all_features[1028] )));
  assign new_n10122_ = ~\all_features[1031]  & (~new_n10120_ | ~\all_features[1024]  | ~\all_features[1025]  | ~\all_features[1030]  | ~new_n10112_);
  assign new_n10123_ = ~new_n10124_ & ~\all_features[1031] ;
  assign new_n10124_ = \all_features[1029]  & \all_features[1030]  & (\all_features[1028]  | (\all_features[1026]  & \all_features[1027]  & \all_features[1025] ));
  assign new_n10125_ = new_n10115_ & ~new_n10126_ & new_n10101_;
  assign new_n10126_ = ~new_n10119_ & ~new_n10121_ & ~new_n10122_ & ~new_n10123_ & (~new_n10110_ | ~new_n10108_);
  assign new_n10127_ = new_n10118_ & new_n10115_ & ~new_n10123_ & ~new_n10122_ & ~new_n10102_ & ~new_n10105_;
  assign new_n10128_ = new_n10129_ & ~new_n10155_ & ~new_n10159_;
  assign new_n10129_ = ~new_n10130_ & ~new_n10153_;
  assign new_n10130_ = new_n10148_ & ~new_n10152_ & ~new_n10131_ & ~new_n10151_;
  assign new_n10131_ = ~new_n10144_ & ~new_n10146_ & new_n10139_ & (~new_n10147_ | ~new_n10132_);
  assign new_n10132_ = new_n10138_ & new_n10133_ & new_n10135_;
  assign new_n10133_ = \all_features[4999]  & (\all_features[4998]  | (new_n10134_ & (\all_features[4994]  | \all_features[4995]  | \all_features[4993] )));
  assign new_n10134_ = \all_features[4996]  & \all_features[4997] ;
  assign new_n10135_ = \all_features[4998]  & \all_features[4999]  & (\all_features[4996]  | \all_features[4997]  | new_n10136_ | ~new_n10137_);
  assign new_n10136_ = \all_features[4992]  & \all_features[4993] ;
  assign new_n10137_ = ~\all_features[4994]  & ~\all_features[4995] ;
  assign new_n10138_ = \all_features[4999]  & (\all_features[4997]  | \all_features[4998]  | \all_features[4996] );
  assign new_n10139_ = ~new_n10140_ & ~new_n10142_;
  assign new_n10140_ = ~\all_features[4999]  & (~\all_features[4998]  | (~\all_features[4996]  & ~\all_features[4997]  & ~new_n10141_));
  assign new_n10141_ = \all_features[4994]  & \all_features[4995] ;
  assign new_n10142_ = ~new_n10143_ & ~\all_features[4999] ;
  assign new_n10143_ = \all_features[4997]  & \all_features[4998]  & (\all_features[4996]  | (\all_features[4994]  & \all_features[4995]  & \all_features[4993] ));
  assign new_n10144_ = ~\all_features[4999]  & (~\all_features[4998]  | (~\all_features[4997]  & (new_n10145_ | ~new_n10141_ | ~\all_features[4996] )));
  assign new_n10145_ = ~\all_features[4992]  & ~\all_features[4993] ;
  assign new_n10146_ = ~\all_features[4999]  & (~\all_features[4998]  | ~new_n10136_ | ~new_n10134_ | ~new_n10141_);
  assign new_n10147_ = \all_features[4999]  & (\all_features[4998]  | (\all_features[4997]  & (\all_features[4996]  | ~new_n10137_ | ~new_n10145_)));
  assign new_n10148_ = ~new_n10149_ & (\all_features[4995]  | \all_features[4996]  | \all_features[4997]  | \all_features[4998]  | \all_features[4999] );
  assign new_n10149_ = ~\all_features[4997]  & new_n10150_ & ((~\all_features[4994]  & new_n10145_) | ~\all_features[4996]  | ~\all_features[4995] );
  assign new_n10150_ = ~\all_features[4998]  & ~\all_features[4999] ;
  assign new_n10151_ = new_n10150_ & (~\all_features[4997]  | (~\all_features[4996]  & (~\all_features[4995]  | (~\all_features[4994]  & ~\all_features[4993] ))));
  assign new_n10152_ = new_n10150_ & (~\all_features[4995]  | ~new_n10134_ | (~\all_features[4994]  & ~new_n10136_));
  assign new_n10153_ = new_n10148_ & new_n10139_ & new_n10154_ & ~new_n10144_ & ~new_n10146_;
  assign new_n10154_ = ~new_n10151_ & ~new_n10152_;
  assign new_n10155_ = ~new_n10156_ & (\all_features[4995]  | \all_features[4996]  | \all_features[4997]  | \all_features[4998]  | \all_features[4999] );
  assign new_n10156_ = ~new_n10149_ & (new_n10151_ | (~new_n10152_ & (new_n10140_ | (~new_n10157_ & ~new_n10144_))));
  assign new_n10157_ = ~new_n10142_ & (new_n10146_ | (new_n10138_ & (~new_n10147_ | (~new_n10158_ & new_n10133_))));
  assign new_n10158_ = ~\all_features[4997]  & \all_features[4998]  & \all_features[4999]  & (\all_features[4996]  ? new_n10137_ : (new_n10136_ | ~new_n10137_));
  assign new_n10159_ = new_n10148_ & (~new_n10154_ | (~new_n10160_ & ~new_n10140_ & ~new_n10144_));
  assign new_n10160_ = ~new_n10142_ & ~new_n10146_ & (~new_n10138_ | ~new_n10147_ | new_n10161_);
  assign new_n10161_ = new_n10133_ & new_n10135_ & (new_n10162_ | ~\all_features[4997]  | ~\all_features[4998]  | ~\all_features[4999] );
  assign new_n10162_ = ~\all_features[4995]  & ~\all_features[4996]  & (~\all_features[4994]  | new_n10145_);
  assign new_n10163_ = ~new_n10164_ & new_n10369_;
  assign new_n10164_ = new_n10165_ & ((~new_n10241_ & new_n10205_) | ~new_n10167_ | (new_n10367_ & ~new_n8434_));
  assign new_n10165_ = ~new_n10166_ & (new_n10167_ | (~new_n10281_ & new_n10343_ & ~new_n9387_) | (new_n10283_ & new_n9387_));
  assign new_n10166_ = new_n10247_ & new_n10167_ & ~new_n10241_ & new_n10205_;
  assign new_n10167_ = ~new_n10168_ & new_n10200_;
  assign new_n10168_ = ~new_n10169_ & ~new_n10190_;
  assign new_n10169_ = ~new_n10170_ & (\all_features[2875]  | \all_features[2876]  | \all_features[2877]  | \all_features[2878]  | \all_features[2879] );
  assign new_n10170_ = ~new_n10184_ & (new_n10186_ | (~new_n10187_ & (new_n10188_ | (~new_n10171_ & ~new_n10189_))));
  assign new_n10171_ = ~new_n10179_ & (new_n10181_ | (~new_n10172_ & new_n10183_));
  assign new_n10172_ = \all_features[2879]  & ((~new_n10177_ & ~\all_features[2877]  & \all_features[2878] ) | (~new_n10175_ & (\all_features[2878]  | (~new_n10173_ & \all_features[2877] ))));
  assign new_n10173_ = new_n10174_ & ~\all_features[2876]  & ~\all_features[2874]  & ~\all_features[2875] ;
  assign new_n10174_ = ~\all_features[2872]  & ~\all_features[2873] ;
  assign new_n10175_ = \all_features[2879]  & (\all_features[2878]  | (new_n10176_ & (\all_features[2874]  | \all_features[2875]  | \all_features[2873] )));
  assign new_n10176_ = \all_features[2876]  & \all_features[2877] ;
  assign new_n10177_ = (\all_features[2876]  & (\all_features[2874]  | \all_features[2875] )) | (~new_n10178_ & ~\all_features[2874]  & ~\all_features[2875]  & ~\all_features[2876] );
  assign new_n10178_ = \all_features[2872]  & \all_features[2873] ;
  assign new_n10179_ = ~new_n10180_ & ~\all_features[2879] ;
  assign new_n10180_ = \all_features[2877]  & \all_features[2878]  & (\all_features[2876]  | (\all_features[2874]  & \all_features[2875]  & \all_features[2873] ));
  assign new_n10181_ = ~\all_features[2879]  & (~\all_features[2878]  | ~new_n10178_ | ~new_n10176_ | ~new_n10182_);
  assign new_n10182_ = \all_features[2874]  & \all_features[2875] ;
  assign new_n10183_ = \all_features[2879]  & (\all_features[2877]  | \all_features[2878]  | \all_features[2876] );
  assign new_n10184_ = ~\all_features[2877]  & new_n10185_ & ((~\all_features[2874]  & new_n10174_) | ~\all_features[2876]  | ~\all_features[2875] );
  assign new_n10185_ = ~\all_features[2878]  & ~\all_features[2879] ;
  assign new_n10186_ = new_n10185_ & (~\all_features[2877]  | (~\all_features[2876]  & (~\all_features[2875]  | (~\all_features[2874]  & ~\all_features[2873] ))));
  assign new_n10187_ = new_n10185_ & (~\all_features[2875]  | ~new_n10176_ | (~\all_features[2874]  & ~new_n10178_));
  assign new_n10188_ = ~\all_features[2879]  & (~\all_features[2878]  | (~\all_features[2876]  & ~\all_features[2877]  & ~new_n10182_));
  assign new_n10189_ = ~\all_features[2879]  & (~\all_features[2878]  | (~\all_features[2877]  & (new_n10174_ | ~new_n10182_ | ~\all_features[2876] )));
  assign new_n10190_ = new_n10196_ & (~new_n10197_ | (new_n10198_ & (~new_n10199_ | new_n10191_)));
  assign new_n10191_ = new_n10192_ & (~new_n10193_ | (~new_n10195_ & \all_features[2877]  & \all_features[2878]  & \all_features[2879] ));
  assign new_n10192_ = \all_features[2879]  & (\all_features[2878]  | (~new_n10173_ & \all_features[2877] ));
  assign new_n10193_ = \all_features[2879]  & \all_features[2878]  & ~new_n10194_ & new_n10175_;
  assign new_n10194_ = ~\all_features[2877]  & ~\all_features[2876]  & ~\all_features[2875]  & ~new_n10178_ & ~\all_features[2874] ;
  assign new_n10195_ = ~\all_features[2875]  & ~\all_features[2876]  & (~\all_features[2874]  | new_n10174_);
  assign new_n10196_ = ~new_n10184_ & (\all_features[2875]  | \all_features[2876]  | \all_features[2877]  | \all_features[2878]  | \all_features[2879] );
  assign new_n10197_ = ~new_n10186_ & ~new_n10187_;
  assign new_n10198_ = ~new_n10188_ & ~new_n10189_;
  assign new_n10199_ = ~new_n10179_ & ~new_n10181_;
  assign new_n10200_ = new_n10201_ & new_n10204_;
  assign new_n10201_ = new_n10202_ & (new_n10189_ | new_n10179_ | ~new_n10203_ | (new_n10193_ & new_n10192_));
  assign new_n10202_ = new_n10196_ & new_n10197_;
  assign new_n10203_ = ~new_n10188_ & ~new_n10181_;
  assign new_n10204_ = new_n10199_ & new_n10202_ & new_n10198_;
  assign new_n10205_ = ~new_n10206_ & ~new_n10240_;
  assign new_n10206_ = ~new_n10207_ & new_n10238_;
  assign new_n10207_ = ~new_n10208_ & ~new_n10229_;
  assign new_n10208_ = ~new_n10225_ & (new_n10222_ | (~new_n10228_ & (new_n10227_ | (~new_n10226_ & ~new_n10209_))));
  assign new_n10209_ = ~new_n10216_ & (new_n10218_ | (~new_n10220_ & (~new_n10221_ | new_n10210_)));
  assign new_n10210_ = \all_features[2839]  & ((~new_n10215_ & ~\all_features[2837]  & \all_features[2838] ) | (~new_n10213_ & (\all_features[2838]  | (~new_n10211_ & \all_features[2837] ))));
  assign new_n10211_ = new_n10212_ & ~\all_features[2836]  & ~\all_features[2834]  & ~\all_features[2835] ;
  assign new_n10212_ = ~\all_features[2832]  & ~\all_features[2833] ;
  assign new_n10213_ = \all_features[2839]  & (\all_features[2838]  | (new_n10214_ & (\all_features[2834]  | \all_features[2835]  | \all_features[2833] )));
  assign new_n10214_ = \all_features[2836]  & \all_features[2837] ;
  assign new_n10215_ = (~\all_features[2834]  & ~\all_features[2835]  & ~\all_features[2836]  & (~\all_features[2833]  | ~\all_features[2832] )) | (\all_features[2836]  & (\all_features[2834]  | \all_features[2835] ));
  assign new_n10216_ = ~\all_features[2839]  & (~\all_features[2838]  | (~\all_features[2837]  & (new_n10212_ | ~\all_features[2836]  | ~new_n10217_)));
  assign new_n10217_ = \all_features[2834]  & \all_features[2835] ;
  assign new_n10218_ = ~new_n10219_ & ~\all_features[2839] ;
  assign new_n10219_ = \all_features[2837]  & \all_features[2838]  & (\all_features[2836]  | (\all_features[2834]  & \all_features[2835]  & \all_features[2833] ));
  assign new_n10220_ = ~\all_features[2839]  & (~new_n10214_ | ~\all_features[2832]  | ~\all_features[2833]  | ~\all_features[2838]  | ~new_n10217_);
  assign new_n10221_ = \all_features[2839]  & (\all_features[2837]  | \all_features[2838]  | \all_features[2836] );
  assign new_n10222_ = new_n10223_ & ((~\all_features[2834]  & new_n10212_) | ~\all_features[2836]  | ~\all_features[2835] );
  assign new_n10223_ = ~\all_features[2837]  & new_n10224_;
  assign new_n10224_ = ~\all_features[2838]  & ~\all_features[2839] ;
  assign new_n10225_ = new_n10223_ & ~\all_features[2835]  & ~\all_features[2836] ;
  assign new_n10226_ = ~\all_features[2839]  & (~\all_features[2838]  | (~\all_features[2836]  & ~\all_features[2837]  & ~new_n10217_));
  assign new_n10227_ = new_n10224_ & (~new_n10214_ | ~\all_features[2835]  | (~\all_features[2834]  & (~\all_features[2832]  | ~\all_features[2833] )));
  assign new_n10228_ = new_n10224_ & (~\all_features[2837]  | (~\all_features[2836]  & (~\all_features[2835]  | (~\all_features[2834]  & ~\all_features[2833] ))));
  assign new_n10229_ = new_n10230_ & (~new_n10237_ | (new_n10236_ & (new_n10231_ | new_n10218_ | new_n10220_)));
  assign new_n10230_ = ~new_n10222_ & ~new_n10225_;
  assign new_n10231_ = new_n10232_ & (~new_n10233_ | (~new_n10235_ & \all_features[2837]  & \all_features[2838]  & \all_features[2839] ));
  assign new_n10232_ = \all_features[2839]  & (\all_features[2838]  | (~new_n10211_ & \all_features[2837] ));
  assign new_n10233_ = \all_features[2839]  & \all_features[2838]  & ~new_n10234_ & new_n10213_;
  assign new_n10234_ = ~\all_features[2834]  & ~\all_features[2835]  & ~\all_features[2836]  & ~\all_features[2837]  & (~\all_features[2833]  | ~\all_features[2832] );
  assign new_n10235_ = ~\all_features[2835]  & ~\all_features[2836]  & (~\all_features[2834]  | new_n10212_);
  assign new_n10236_ = ~new_n10226_ & ~new_n10216_;
  assign new_n10237_ = ~new_n10227_ & ~new_n10228_;
  assign new_n10238_ = new_n10237_ & ~new_n10239_ & new_n10230_;
  assign new_n10239_ = ~new_n10226_ & ~new_n10216_ & ~new_n10218_ & ~new_n10220_ & (~new_n10233_ | ~new_n10232_);
  assign new_n10240_ = new_n10237_ & new_n10236_ & ~new_n10220_ & ~new_n10218_ & ~new_n10222_ & ~new_n10225_;
  assign new_n10241_ = new_n10242_ & ~new_n6760_ & ~new_n10243_;
  assign new_n10242_ = ~new_n6738_ & ~new_n6766_;
  assign new_n10243_ = ~new_n10244_ & (\all_features[3867]  | \all_features[3868]  | \all_features[3869]  | \all_features[3870]  | \all_features[3871] );
  assign new_n10244_ = ~new_n6759_ & (new_n6758_ | (~new_n6756_ & (new_n6743_ | (~new_n6753_ & ~new_n10245_))));
  assign new_n10245_ = ~new_n6741_ & (new_n6745_ | (new_n6754_ & (~new_n6748_ | (~new_n10246_ & new_n6751_))));
  assign new_n10246_ = ~\all_features[3869]  & \all_features[3870]  & \all_features[3871]  & (\all_features[3868]  ? new_n6749_ : (new_n6747_ | ~new_n6749_));
  assign new_n10247_ = new_n10248_ & new_n10272_;
  assign new_n10248_ = ~new_n10249_ & ~new_n10271_;
  assign new_n10249_ = new_n10250_ & (~new_n10259_ | (new_n10269_ & new_n10270_ & new_n10266_ & new_n10268_));
  assign new_n10250_ = new_n10251_ & ~new_n10255_ & ~new_n10256_;
  assign new_n10251_ = ~new_n10252_ & (\all_features[2755]  | \all_features[2756]  | \all_features[2757]  | \all_features[2758]  | \all_features[2759] );
  assign new_n10252_ = ~\all_features[2757]  & new_n10254_ & ((~\all_features[2754]  & new_n10253_) | ~\all_features[2756]  | ~\all_features[2755] );
  assign new_n10253_ = ~\all_features[2752]  & ~\all_features[2753] ;
  assign new_n10254_ = ~\all_features[2758]  & ~\all_features[2759] ;
  assign new_n10255_ = new_n10254_ & (~\all_features[2757]  | (~\all_features[2756]  & (~\all_features[2755]  | (~\all_features[2754]  & ~\all_features[2753] ))));
  assign new_n10256_ = new_n10254_ & (~\all_features[2755]  | ~new_n10257_ | (~\all_features[2754]  & ~new_n10258_));
  assign new_n10257_ = \all_features[2756]  & \all_features[2757] ;
  assign new_n10258_ = \all_features[2752]  & \all_features[2753] ;
  assign new_n10259_ = ~new_n10265_ & ~new_n10264_ & ~new_n10260_ & ~new_n10262_;
  assign new_n10260_ = ~\all_features[2759]  & (~\all_features[2758]  | (~\all_features[2757]  & (new_n10253_ | ~new_n10261_ | ~\all_features[2756] )));
  assign new_n10261_ = \all_features[2754]  & \all_features[2755] ;
  assign new_n10262_ = ~new_n10263_ & ~\all_features[2759] ;
  assign new_n10263_ = \all_features[2757]  & \all_features[2758]  & (\all_features[2756]  | (\all_features[2754]  & \all_features[2755]  & \all_features[2753] ));
  assign new_n10264_ = ~\all_features[2759]  & (~\all_features[2758]  | ~new_n10257_ | ~new_n10258_ | ~new_n10261_);
  assign new_n10265_ = ~\all_features[2759]  & (~\all_features[2758]  | (~\all_features[2756]  & ~\all_features[2757]  & ~new_n10261_));
  assign new_n10266_ = \all_features[2759]  & (\all_features[2758]  | (\all_features[2757]  & (\all_features[2756]  | ~new_n10253_ | ~new_n10267_)));
  assign new_n10267_ = ~\all_features[2754]  & ~\all_features[2755] ;
  assign new_n10268_ = \all_features[2759]  & (\all_features[2758]  | (new_n10257_ & (\all_features[2754]  | \all_features[2755]  | \all_features[2753] )));
  assign new_n10269_ = \all_features[2758]  & \all_features[2759]  & (\all_features[2756]  | \all_features[2757]  | new_n10258_ | ~new_n10267_);
  assign new_n10270_ = \all_features[2759]  & (\all_features[2757]  | \all_features[2758]  | \all_features[2756] );
  assign new_n10271_ = new_n10250_ & new_n10259_;
  assign new_n10272_ = ~new_n10273_ & ~new_n10277_;
  assign new_n10273_ = new_n10251_ & (new_n10256_ | new_n10255_ | (~new_n10260_ & ~new_n10265_ & ~new_n10274_));
  assign new_n10274_ = ~new_n10264_ & ~new_n10262_ & (~new_n10270_ | ~new_n10266_ | new_n10275_);
  assign new_n10275_ = new_n10268_ & new_n10269_ & (new_n10276_ | ~\all_features[2757]  | ~\all_features[2758]  | ~\all_features[2759] );
  assign new_n10276_ = ~\all_features[2755]  & ~\all_features[2756]  & (~\all_features[2754]  | new_n10253_);
  assign new_n10277_ = ~new_n10278_ & (\all_features[2755]  | \all_features[2756]  | \all_features[2757]  | \all_features[2758]  | \all_features[2759] );
  assign new_n10278_ = ~new_n10252_ & (new_n10255_ | (~new_n10256_ & (new_n10265_ | (~new_n10260_ & ~new_n10279_))));
  assign new_n10279_ = ~new_n10262_ & (new_n10264_ | (new_n10270_ & (~new_n10266_ | (~new_n10280_ & new_n10268_))));
  assign new_n10280_ = ~\all_features[2757]  & \all_features[2758]  & \all_features[2759]  & (\all_features[2756]  ? new_n10267_ : (new_n10258_ | ~new_n10267_));
  assign new_n10281_ = new_n8264_ & ~new_n10282_ & new_n8232_;
  assign new_n10282_ = ~new_n8255_ & ~new_n8260_;
  assign new_n10283_ = new_n10284_ & (new_n10335_ | new_n10339_ | ~new_n10310_);
  assign new_n10284_ = ~new_n10285_ & ~new_n10308_;
  assign new_n10285_ = new_n10303_ & ~new_n10307_ & ~new_n10286_ & ~new_n10306_;
  assign new_n10286_ = ~new_n10301_ & ~new_n10302_ & new_n10294_ & (~new_n10299_ | ~new_n10287_);
  assign new_n10287_ = new_n10293_ & new_n10288_ & new_n10290_;
  assign new_n10288_ = \all_features[5471]  & (\all_features[5470]  | (new_n10289_ & (\all_features[5466]  | \all_features[5467]  | \all_features[5465] )));
  assign new_n10289_ = \all_features[5468]  & \all_features[5469] ;
  assign new_n10290_ = \all_features[5470]  & \all_features[5471]  & (\all_features[5468]  | \all_features[5469]  | new_n10292_ | ~new_n10291_);
  assign new_n10291_ = ~\all_features[5466]  & ~\all_features[5467] ;
  assign new_n10292_ = \all_features[5464]  & \all_features[5465] ;
  assign new_n10293_ = \all_features[5471]  & (\all_features[5469]  | \all_features[5470]  | \all_features[5468] );
  assign new_n10294_ = ~new_n10295_ & ~new_n10297_;
  assign new_n10295_ = ~new_n10296_ & ~\all_features[5471] ;
  assign new_n10296_ = \all_features[5469]  & \all_features[5470]  & (\all_features[5468]  | (\all_features[5466]  & \all_features[5467]  & \all_features[5465] ));
  assign new_n10297_ = ~\all_features[5471]  & (~\all_features[5470]  | (~\all_features[5468]  & ~\all_features[5469]  & ~new_n10298_));
  assign new_n10298_ = \all_features[5466]  & \all_features[5467] ;
  assign new_n10299_ = \all_features[5471]  & (\all_features[5470]  | (\all_features[5469]  & (\all_features[5468]  | ~new_n10300_ | ~new_n10291_)));
  assign new_n10300_ = ~\all_features[5464]  & ~\all_features[5465] ;
  assign new_n10301_ = ~\all_features[5471]  & (~\all_features[5470]  | (~\all_features[5469]  & (new_n10300_ | ~new_n10298_ | ~\all_features[5468] )));
  assign new_n10302_ = ~\all_features[5471]  & (~\all_features[5470]  | ~new_n10289_ | ~new_n10292_ | ~new_n10298_);
  assign new_n10303_ = ~new_n10304_ & (\all_features[5467]  | \all_features[5468]  | \all_features[5469]  | \all_features[5470]  | \all_features[5471] );
  assign new_n10304_ = ~\all_features[5469]  & new_n10305_ & ((~\all_features[5466]  & new_n10300_) | ~\all_features[5468]  | ~\all_features[5467] );
  assign new_n10305_ = ~\all_features[5470]  & ~\all_features[5471] ;
  assign new_n10306_ = new_n10305_ & (~\all_features[5469]  | (~\all_features[5468]  & (~\all_features[5467]  | (~\all_features[5466]  & ~\all_features[5465] ))));
  assign new_n10307_ = new_n10305_ & (~\all_features[5467]  | ~new_n10289_ | (~\all_features[5466]  & ~new_n10292_));
  assign new_n10308_ = new_n10303_ & new_n10294_ & new_n10309_ & ~new_n10301_ & ~new_n10302_;
  assign new_n10309_ = ~new_n10306_ & ~new_n10307_;
  assign new_n10310_ = ~new_n10311_ & ~new_n10333_;
  assign new_n10311_ = new_n10328_ & ~new_n10332_ & ~new_n10312_ & ~new_n10331_;
  assign new_n10312_ = new_n10313_ & (~new_n10326_ | ~new_n10327_ | ~new_n10323_ | ~new_n10325_);
  assign new_n10313_ = ~new_n10320_ & ~new_n10318_ & ~new_n10314_ & ~new_n10316_;
  assign new_n10314_ = ~\all_features[5727]  & (~\all_features[5726]  | (~\all_features[5724]  & ~\all_features[5725]  & ~new_n10315_));
  assign new_n10315_ = \all_features[5722]  & \all_features[5723] ;
  assign new_n10316_ = ~\all_features[5727]  & (~\all_features[5726]  | (~\all_features[5725]  & (new_n10317_ | ~new_n10315_ | ~\all_features[5724] )));
  assign new_n10317_ = ~\all_features[5720]  & ~\all_features[5721] ;
  assign new_n10318_ = ~new_n10319_ & ~\all_features[5727] ;
  assign new_n10319_ = \all_features[5725]  & \all_features[5726]  & (\all_features[5724]  | (\all_features[5722]  & \all_features[5723]  & \all_features[5721] ));
  assign new_n10320_ = ~\all_features[5727]  & (~\all_features[5726]  | ~new_n10321_ | ~new_n10322_ | ~new_n10315_);
  assign new_n10321_ = \all_features[5720]  & \all_features[5721] ;
  assign new_n10322_ = \all_features[5724]  & \all_features[5725] ;
  assign new_n10323_ = \all_features[5727]  & (\all_features[5726]  | (\all_features[5725]  & (\all_features[5724]  | ~new_n10324_ | ~new_n10317_)));
  assign new_n10324_ = ~\all_features[5722]  & ~\all_features[5723] ;
  assign new_n10325_ = \all_features[5727]  & (\all_features[5726]  | (new_n10322_ & (\all_features[5722]  | \all_features[5723]  | \all_features[5721] )));
  assign new_n10326_ = \all_features[5726]  & \all_features[5727]  & (\all_features[5724]  | \all_features[5725]  | new_n10321_ | ~new_n10324_);
  assign new_n10327_ = \all_features[5727]  & (\all_features[5725]  | \all_features[5726]  | \all_features[5724] );
  assign new_n10328_ = ~new_n10329_ & (\all_features[5723]  | \all_features[5724]  | \all_features[5725]  | \all_features[5726]  | \all_features[5727] );
  assign new_n10329_ = ~\all_features[5725]  & new_n10330_ & ((~\all_features[5722]  & new_n10317_) | ~\all_features[5724]  | ~\all_features[5723] );
  assign new_n10330_ = ~\all_features[5726]  & ~\all_features[5727] ;
  assign new_n10331_ = new_n10330_ & (~\all_features[5725]  | (~\all_features[5724]  & (~\all_features[5723]  | (~\all_features[5722]  & ~\all_features[5721] ))));
  assign new_n10332_ = new_n10330_ & (~\all_features[5723]  | ~new_n10322_ | (~\all_features[5722]  & ~new_n10321_));
  assign new_n10333_ = new_n10334_ & new_n10328_ & ~new_n10331_ & ~new_n10318_;
  assign new_n10334_ = ~new_n10320_ & ~new_n10316_ & ~new_n10332_ & ~new_n10314_;
  assign new_n10335_ = ~new_n10336_ & (\all_features[5723]  | \all_features[5724]  | \all_features[5725]  | \all_features[5726]  | \all_features[5727] );
  assign new_n10336_ = ~new_n10329_ & (new_n10331_ | (~new_n10332_ & (new_n10314_ | (~new_n10337_ & ~new_n10316_))));
  assign new_n10337_ = ~new_n10318_ & (new_n10320_ | (new_n10327_ & (~new_n10323_ | (~new_n10338_ & new_n10325_))));
  assign new_n10338_ = ~\all_features[5725]  & \all_features[5726]  & \all_features[5727]  & (\all_features[5724]  ? new_n10324_ : (new_n10321_ | ~new_n10324_));
  assign new_n10339_ = new_n10328_ & (new_n10332_ | new_n10331_ | (~new_n10340_ & ~new_n10314_ & ~new_n10316_));
  assign new_n10340_ = ~new_n10318_ & ~new_n10320_ & (~new_n10327_ | ~new_n10323_ | new_n10341_);
  assign new_n10341_ = new_n10325_ & new_n10326_ & (new_n10342_ | ~\all_features[5725]  | ~\all_features[5726]  | ~\all_features[5727] );
  assign new_n10342_ = ~\all_features[5723]  & ~\all_features[5724]  & (~\all_features[5722]  | new_n10317_);
  assign new_n10343_ = new_n10351_ | ~new_n10361_ | (~new_n10360_ & new_n10344_);
  assign new_n10344_ = ~new_n10345_ & ~new_n10351_ & new_n10354_ & (\all_features[3991]  | new_n10357_);
  assign new_n10345_ = \all_features[3991]  & \all_features[3990]  & ~new_n10346_ & new_n10348_;
  assign new_n10346_ = ~\all_features[3989]  & ~\all_features[3988]  & ~\all_features[3987]  & ~new_n10347_ & ~\all_features[3986] ;
  assign new_n10347_ = \all_features[3984]  & \all_features[3985] ;
  assign new_n10348_ = \all_features[3991]  & (\all_features[3990]  | (~new_n10349_ & \all_features[3989]  & \all_features[3988] ));
  assign new_n10349_ = ~\all_features[3987]  & ~\all_features[3985]  & ~\all_features[3986] ;
  assign new_n10351_ = ~\all_features[3991]  & (~\all_features[3990]  | new_n10352_);
  assign new_n10352_ = ~\all_features[3989]  & (~\all_features[3988]  | ~new_n10353_ | (~\all_features[3985]  & ~\all_features[3984] ));
  assign new_n10353_ = \all_features[3986]  & \all_features[3987] ;
  assign new_n10354_ = \all_features[3991]  | (~new_n10355_ & new_n10347_ & \all_features[3990]  & new_n10356_);
  assign new_n10355_ = ~\all_features[3989]  & ~new_n10353_ & ~\all_features[3988] ;
  assign new_n10356_ = \all_features[3989]  & new_n10353_ & \all_features[3988] ;
  assign new_n10357_ = \all_features[3989]  & \all_features[3990]  & (\all_features[3988]  | (\all_features[3986]  & \all_features[3987]  & \all_features[3985] ));
  assign new_n10360_ = \all_features[3991]  | (\all_features[3990]  & new_n10356_ & new_n10347_ & new_n10357_);
  assign new_n10361_ = new_n10362_ & (\all_features[3991]  | (~new_n10355_ & \all_features[3990] ));
  assign new_n10362_ = \all_features[3989]  | \all_features[3990]  | \all_features[3991]  | (\all_features[3988]  & \all_features[3987]  & ~new_n10363_);
  assign new_n10363_ = ~\all_features[3986]  & ~\all_features[3984]  & ~\all_features[3985] ;
  assign new_n10367_ = new_n10241_ & (~new_n8097_ | (~new_n8094_ & new_n10368_));
  assign new_n10368_ = ~new_n8062_ & ~new_n8083_;
  assign new_n10369_ = new_n10370_ & (new_n8434_ | ~new_n10167_ | ~new_n10367_);
  assign new_n10370_ = new_n10167_ | ((new_n10281_ | ~new_n10343_ | new_n9387_) & (~new_n10283_ | ~new_n9387_));
  assign new_n10371_ = new_n10372_ ? (~new_n12043_ ^ new_n12260_) : (new_n12043_ ^ new_n12260_);
  assign new_n10372_ = new_n10373_ ? (~new_n11126_ ^ new_n11721_) : (new_n11126_ ^ new_n11721_);
  assign new_n10373_ = new_n10374_ ? (~new_n10641_ ^ new_n10835_) : (new_n10641_ ^ new_n10835_);
  assign new_n10374_ = ~new_n10375_ & new_n10638_;
  assign new_n10375_ = new_n10376_ & new_n10535_ & (~new_n10637_ | ~new_n10636_);
  assign new_n10376_ = new_n10397_ & (~new_n10377_ | (~new_n10524_ & new_n10454_) | (~new_n10489_ & ~new_n10454_));
  assign new_n10377_ = ~new_n10378_ & new_n8892_;
  assign new_n10378_ = ~new_n10379_ & ~new_n8391_;
  assign new_n10379_ = new_n10380_ & new_n10395_;
  assign new_n10380_ = new_n10381_ & new_n10389_;
  assign new_n10381_ = ~new_n10382_ & (\all_features[1419]  | \all_features[1420]  | \all_features[1421]  | \all_features[1422]  | \all_features[1423] );
  assign new_n10382_ = ~new_n8393_ & (new_n8404_ | (~new_n8406_ & (new_n8401_ | (~new_n8405_ & ~new_n10383_))));
  assign new_n10383_ = ~new_n8402_ & (new_n8397_ | (new_n10388_ & (~new_n10384_ | (~new_n10387_ & new_n10386_))));
  assign new_n10384_ = \all_features[1423]  & (\all_features[1422]  | (\all_features[1421]  & (\all_features[1420]  | ~new_n10385_ | ~new_n8395_)));
  assign new_n10385_ = ~\all_features[1418]  & ~\all_features[1419] ;
  assign new_n10386_ = \all_features[1423]  & (\all_features[1422]  | (new_n8400_ & (\all_features[1418]  | \all_features[1419]  | \all_features[1417] )));
  assign new_n10387_ = ~\all_features[1421]  & \all_features[1422]  & \all_features[1423]  & (\all_features[1420]  ? new_n10385_ : (new_n8399_ | ~new_n10385_));
  assign new_n10388_ = \all_features[1423]  & (\all_features[1421]  | \all_features[1422]  | \all_features[1420] );
  assign new_n10389_ = new_n8392_ & (~new_n10394_ | (~new_n10390_ & ~new_n8405_ & ~new_n8401_));
  assign new_n10390_ = ~new_n8402_ & ~new_n8397_ & (~new_n10388_ | ~new_n10384_ | new_n10391_);
  assign new_n10391_ = new_n10386_ & new_n10392_ & (new_n10393_ | ~\all_features[1421]  | ~\all_features[1422]  | ~\all_features[1423] );
  assign new_n10392_ = \all_features[1422]  & \all_features[1423]  & (\all_features[1420]  | \all_features[1421]  | new_n8399_ | ~new_n10385_);
  assign new_n10393_ = ~\all_features[1419]  & ~\all_features[1420]  & (~\all_features[1418]  | new_n8395_);
  assign new_n10394_ = ~new_n8404_ & ~new_n8406_;
  assign new_n10395_ = new_n8392_ & new_n10394_ & (new_n10396_ | new_n8402_ | new_n8405_ | ~new_n8396_);
  assign new_n10396_ = new_n10388_ & new_n10392_ & new_n10384_ & new_n10386_;
  assign new_n10397_ = ~new_n10378_ | ((new_n10407_ | new_n10398_) & (new_n10438_ | ~new_n7698_ | ~new_n10398_));
  assign new_n10398_ = new_n10399_ & new_n8483_;
  assign new_n10399_ = ~new_n10400_ & (\all_features[3323]  | \all_features[3324]  | \all_features[3325]  | \all_features[3326]  | \all_features[3327] );
  assign new_n10400_ = new_n10406_ & (new_n8499_ | (~new_n8494_ & new_n10401_ & (new_n8496_ | new_n10404_)));
  assign new_n10401_ = ~new_n8496_ & ~new_n8498_ & (~new_n8505_ | ~new_n8500_ | new_n10402_);
  assign new_n10402_ = new_n8502_ & ~new_n10403_ & new_n8503_;
  assign new_n10403_ = new_n8504_ & \all_features[3325]  & ((~new_n8487_ & \all_features[3322] ) | \all_features[3324]  | \all_features[3323] );
  assign new_n10404_ = ~new_n8498_ & (~new_n8505_ | (new_n8500_ & (~new_n8502_ | (~new_n10405_ & new_n8503_))));
  assign new_n10405_ = new_n8504_ & (\all_features[3325]  | (~new_n8501_ & \all_features[3324] ));
  assign new_n10406_ = ~new_n8486_ & ~new_n8489_ & ~new_n8490_;
  assign new_n10407_ = ~new_n10434_ & new_n10408_;
  assign new_n10408_ = ~new_n10409_ & ~new_n10432_;
  assign new_n10409_ = new_n10429_ & ~new_n10410_ & new_n10426_;
  assign new_n10410_ = ~new_n10425_ & ~new_n10423_ & ~new_n10422_ & ~new_n10411_ & ~new_n10414_;
  assign new_n10411_ = ~\all_features[2783]  & (~\all_features[2782]  | new_n10412_);
  assign new_n10412_ = ~\all_features[2781]  & (new_n10413_ | ~\all_features[2779]  | ~\all_features[2780]  | ~\all_features[2778] );
  assign new_n10413_ = ~\all_features[2776]  & ~\all_features[2777] ;
  assign new_n10414_ = new_n10421_ & new_n10420_ & new_n10415_ & new_n10417_;
  assign new_n10415_ = \all_features[2783]  & (\all_features[2782]  | (new_n10416_ & (\all_features[2778]  | \all_features[2779]  | \all_features[2777] )));
  assign new_n10416_ = \all_features[2780]  & \all_features[2781] ;
  assign new_n10417_ = \all_features[2782]  & \all_features[2783]  & (\all_features[2780]  | \all_features[2781]  | new_n10419_ | ~new_n10418_);
  assign new_n10418_ = ~\all_features[2778]  & ~\all_features[2779] ;
  assign new_n10419_ = \all_features[2776]  & \all_features[2777] ;
  assign new_n10420_ = \all_features[2783]  & (\all_features[2782]  | (\all_features[2781]  & (\all_features[2780]  | ~new_n10418_ | ~new_n10413_)));
  assign new_n10421_ = \all_features[2783]  & (\all_features[2781]  | \all_features[2782]  | \all_features[2780] );
  assign new_n10422_ = ~\all_features[2783]  & (~new_n10419_ | ~\all_features[2778]  | ~\all_features[2779]  | ~\all_features[2782]  | ~new_n10416_);
  assign new_n10423_ = ~new_n10424_ & ~\all_features[2783] ;
  assign new_n10424_ = \all_features[2781]  & \all_features[2782]  & (\all_features[2780]  | (\all_features[2778]  & \all_features[2779]  & \all_features[2777] ));
  assign new_n10425_ = ~\all_features[2783]  & (~\all_features[2782]  | (~\all_features[2781]  & ~\all_features[2780]  & (~\all_features[2779]  | ~\all_features[2778] )));
  assign new_n10426_ = ~new_n10427_ & (\all_features[2779]  | \all_features[2780]  | \all_features[2781]  | \all_features[2782]  | \all_features[2783] );
  assign new_n10427_ = ~\all_features[2781]  & new_n10428_ & ((~\all_features[2778]  & new_n10413_) | ~\all_features[2780]  | ~\all_features[2779] );
  assign new_n10428_ = ~\all_features[2782]  & ~\all_features[2783] ;
  assign new_n10429_ = ~new_n10430_ & ~new_n10431_;
  assign new_n10430_ = new_n10428_ & (~\all_features[2779]  | ~new_n10416_ | (~new_n10419_ & ~\all_features[2778] ));
  assign new_n10431_ = new_n10428_ & (~\all_features[2781]  | (~\all_features[2780]  & (~\all_features[2779]  | (~\all_features[2778]  & ~\all_features[2777] ))));
  assign new_n10432_ = new_n10426_ & new_n10433_ & ~new_n10423_ & ~new_n10431_;
  assign new_n10433_ = ~new_n10425_ & ~new_n10430_ & ~new_n10411_ & ~new_n10422_;
  assign new_n10434_ = new_n10426_ & (~new_n10429_ | (~new_n10411_ & ~new_n10435_ & ~new_n10425_));
  assign new_n10435_ = ~new_n10423_ & ~new_n10422_ & (~new_n10421_ | ~new_n10420_ | new_n10436_);
  assign new_n10436_ = new_n10415_ & new_n10417_ & (new_n10437_ | ~\all_features[2781]  | ~\all_features[2782]  | ~\all_features[2783] );
  assign new_n10437_ = ~\all_features[2779]  & ~\all_features[2780]  & (~\all_features[2778]  | new_n10413_);
  assign new_n10438_ = new_n10439_ & ~new_n10453_ & ~new_n10452_ & ~new_n10449_ & ~new_n10451_;
  assign new_n10439_ = ~new_n10448_ & ~new_n10444_ & ~new_n10440_ & ~new_n10442_;
  assign new_n10440_ = ~new_n10441_ & ~\all_features[4799] ;
  assign new_n10441_ = \all_features[4797]  & \all_features[4798]  & (\all_features[4796]  | (\all_features[4794]  & \all_features[4795]  & \all_features[4793] ));
  assign new_n10442_ = new_n10443_ & (~\all_features[4797]  | (~\all_features[4796]  & (~\all_features[4795]  | (~\all_features[4794]  & ~\all_features[4793] ))));
  assign new_n10443_ = ~\all_features[4798]  & ~\all_features[4799] ;
  assign new_n10444_ = ~\all_features[4799]  & (~\all_features[4798]  | ~new_n10445_ | ~new_n10446_ | ~new_n10447_);
  assign new_n10445_ = \all_features[4792]  & \all_features[4793] ;
  assign new_n10446_ = \all_features[4796]  & \all_features[4797] ;
  assign new_n10447_ = \all_features[4794]  & \all_features[4795] ;
  assign new_n10448_ = ~\all_features[4799]  & ~\all_features[4798]  & ~\all_features[4797]  & ~\all_features[4795]  & ~\all_features[4796] ;
  assign new_n10449_ = ~\all_features[4799]  & (~\all_features[4798]  | (~\all_features[4797]  & (new_n10450_ | ~\all_features[4796]  | ~new_n10447_)));
  assign new_n10450_ = ~\all_features[4792]  & ~\all_features[4793] ;
  assign new_n10451_ = ~\all_features[4799]  & (~\all_features[4798]  | (~\all_features[4796]  & ~\all_features[4797]  & ~new_n10447_));
  assign new_n10452_ = ~\all_features[4797]  & new_n10443_ & ((~\all_features[4794]  & new_n10450_) | ~\all_features[4796]  | ~\all_features[4795] );
  assign new_n10453_ = new_n10443_ & (~\all_features[4795]  | ~new_n10446_ | (~\all_features[4794]  & ~new_n10445_));
  assign new_n10454_ = new_n10455_ & (new_n10485_ | new_n10481_);
  assign new_n10455_ = new_n10456_ & new_n10478_;
  assign new_n10456_ = new_n10473_ & ~new_n10477_ & ~new_n10457_ & ~new_n10476_;
  assign new_n10457_ = new_n10458_ & ~new_n10471_ & (~new_n10466_ | ~new_n10472_ | ~new_n10469_ | ~new_n10470_);
  assign new_n10458_ = ~new_n10463_ & ~new_n10459_ & ~new_n10461_;
  assign new_n10459_ = ~new_n10460_ & ~\all_features[4383] ;
  assign new_n10460_ = \all_features[4381]  & \all_features[4382]  & (\all_features[4380]  | (\all_features[4378]  & \all_features[4379]  & \all_features[4377] ));
  assign new_n10461_ = ~\all_features[4383]  & (~\all_features[4382]  | (~\all_features[4380]  & ~\all_features[4381]  & ~new_n10462_));
  assign new_n10462_ = \all_features[4378]  & \all_features[4379] ;
  assign new_n10463_ = ~\all_features[4383]  & (~\all_features[4382]  | ~new_n10464_ | ~new_n10465_ | ~new_n10462_);
  assign new_n10464_ = \all_features[4380]  & \all_features[4381] ;
  assign new_n10465_ = \all_features[4376]  & \all_features[4377] ;
  assign new_n10466_ = \all_features[4383]  & (\all_features[4382]  | (\all_features[4381]  & (\all_features[4380]  | ~new_n10468_ | ~new_n10467_)));
  assign new_n10467_ = ~\all_features[4378]  & ~\all_features[4379] ;
  assign new_n10468_ = ~\all_features[4376]  & ~\all_features[4377] ;
  assign new_n10469_ = \all_features[4383]  & (\all_features[4382]  | (new_n10464_ & (\all_features[4378]  | \all_features[4379]  | \all_features[4377] )));
  assign new_n10470_ = \all_features[4382]  & \all_features[4383]  & (\all_features[4380]  | \all_features[4381]  | new_n10465_ | ~new_n10467_);
  assign new_n10471_ = ~\all_features[4383]  & (~\all_features[4382]  | (~\all_features[4381]  & (new_n10468_ | ~new_n10462_ | ~\all_features[4380] )));
  assign new_n10472_ = \all_features[4383]  & (\all_features[4381]  | \all_features[4382]  | \all_features[4380] );
  assign new_n10473_ = ~new_n10474_ & (\all_features[4379]  | \all_features[4380]  | \all_features[4381]  | \all_features[4382]  | \all_features[4383] );
  assign new_n10474_ = new_n10475_ & (~\all_features[4379]  | ~new_n10464_ | (~\all_features[4378]  & ~new_n10465_));
  assign new_n10475_ = ~\all_features[4382]  & ~\all_features[4383] ;
  assign new_n10476_ = new_n10475_ & (~\all_features[4381]  | (~\all_features[4380]  & (~\all_features[4379]  | (~\all_features[4378]  & ~\all_features[4377] ))));
  assign new_n10477_ = ~\all_features[4381]  & new_n10475_ & ((~\all_features[4378]  & new_n10468_) | ~\all_features[4380]  | ~\all_features[4379] );
  assign new_n10478_ = new_n10458_ & new_n10480_ & ~new_n10471_ & new_n10479_;
  assign new_n10479_ = ~new_n10477_ & (\all_features[4379]  | \all_features[4380]  | \all_features[4381]  | \all_features[4382]  | \all_features[4383] );
  assign new_n10480_ = ~new_n10476_ & ~new_n10474_;
  assign new_n10481_ = new_n10479_ & (~new_n10480_ | (~new_n10482_ & ~new_n10471_ & ~new_n10461_));
  assign new_n10482_ = ~new_n10463_ & ~new_n10459_ & (~new_n10472_ | ~new_n10466_ | new_n10483_);
  assign new_n10483_ = new_n10469_ & new_n10470_ & (new_n10484_ | ~\all_features[4381]  | ~\all_features[4382]  | ~\all_features[4383] );
  assign new_n10484_ = ~\all_features[4379]  & ~\all_features[4380]  & (~\all_features[4378]  | new_n10468_);
  assign new_n10485_ = ~new_n10486_ & (\all_features[4379]  | \all_features[4380]  | \all_features[4381]  | \all_features[4382]  | \all_features[4383] );
  assign new_n10486_ = ~new_n10477_ & (new_n10476_ | (~new_n10474_ & (new_n10461_ | (~new_n10471_ & ~new_n10487_))));
  assign new_n10487_ = ~new_n10459_ & (new_n10463_ | (new_n10472_ & (~new_n10466_ | (~new_n10488_ & new_n10469_))));
  assign new_n10488_ = ~\all_features[4381]  & \all_features[4382]  & \all_features[4383]  & (\all_features[4380]  ? new_n10467_ : (new_n10465_ | ~new_n10467_));
  assign new_n10489_ = new_n10490_ & (~new_n10520_ | ~new_n10516_);
  assign new_n10490_ = ~new_n10491_ & ~new_n10513_;
  assign new_n10491_ = new_n10508_ & ~new_n10512_ & ~new_n10492_ & ~new_n10511_;
  assign new_n10492_ = new_n10493_ & ~new_n10506_ & (~new_n10501_ | ~new_n10507_ | ~new_n10504_ | ~new_n10505_);
  assign new_n10493_ = ~new_n10498_ & ~new_n10494_ & ~new_n10496_;
  assign new_n10494_ = ~new_n10495_ & ~\all_features[3247] ;
  assign new_n10495_ = \all_features[3245]  & \all_features[3246]  & (\all_features[3244]  | (\all_features[3242]  & \all_features[3243]  & \all_features[3241] ));
  assign new_n10496_ = ~\all_features[3247]  & (~\all_features[3246]  | (~\all_features[3244]  & ~\all_features[3245]  & ~new_n10497_));
  assign new_n10497_ = \all_features[3242]  & \all_features[3243] ;
  assign new_n10498_ = ~\all_features[3247]  & (~\all_features[3246]  | ~new_n10499_ | ~new_n10500_ | ~new_n10497_);
  assign new_n10499_ = \all_features[3244]  & \all_features[3245] ;
  assign new_n10500_ = \all_features[3240]  & \all_features[3241] ;
  assign new_n10501_ = \all_features[3247]  & (\all_features[3246]  | (\all_features[3245]  & (\all_features[3244]  | ~new_n10503_ | ~new_n10502_)));
  assign new_n10502_ = ~\all_features[3242]  & ~\all_features[3243] ;
  assign new_n10503_ = ~\all_features[3240]  & ~\all_features[3241] ;
  assign new_n10504_ = \all_features[3247]  & (\all_features[3246]  | (new_n10499_ & (\all_features[3242]  | \all_features[3243]  | \all_features[3241] )));
  assign new_n10505_ = \all_features[3246]  & \all_features[3247]  & (\all_features[3244]  | \all_features[3245]  | new_n10500_ | ~new_n10502_);
  assign new_n10506_ = ~\all_features[3247]  & (~\all_features[3246]  | (~\all_features[3245]  & (new_n10503_ | ~new_n10497_ | ~\all_features[3244] )));
  assign new_n10507_ = \all_features[3247]  & (\all_features[3245]  | \all_features[3246]  | \all_features[3244] );
  assign new_n10508_ = ~new_n10509_ & (\all_features[3243]  | \all_features[3244]  | \all_features[3245]  | \all_features[3246]  | \all_features[3247] );
  assign new_n10509_ = new_n10510_ & (~\all_features[3243]  | ~new_n10499_ | (~\all_features[3242]  & ~new_n10500_));
  assign new_n10510_ = ~\all_features[3246]  & ~\all_features[3247] ;
  assign new_n10511_ = new_n10510_ & (~\all_features[3245]  | (~\all_features[3244]  & (~\all_features[3243]  | (~\all_features[3242]  & ~\all_features[3241] ))));
  assign new_n10512_ = ~\all_features[3245]  & new_n10510_ & ((~\all_features[3242]  & new_n10503_) | ~\all_features[3244]  | ~\all_features[3243] );
  assign new_n10513_ = new_n10493_ & new_n10515_ & ~new_n10506_ & new_n10514_;
  assign new_n10514_ = ~new_n10512_ & (\all_features[3243]  | \all_features[3244]  | \all_features[3245]  | \all_features[3246]  | \all_features[3247] );
  assign new_n10515_ = ~new_n10511_ & ~new_n10509_;
  assign new_n10516_ = new_n10514_ & (~new_n10515_ | (~new_n10517_ & ~new_n10506_ & ~new_n10496_));
  assign new_n10517_ = ~new_n10498_ & ~new_n10494_ & (~new_n10507_ | ~new_n10501_ | new_n10518_);
  assign new_n10518_ = new_n10504_ & new_n10505_ & (new_n10519_ | ~\all_features[3245]  | ~\all_features[3246]  | ~\all_features[3247] );
  assign new_n10519_ = ~\all_features[3243]  & ~\all_features[3244]  & (~\all_features[3242]  | new_n10503_);
  assign new_n10520_ = ~new_n10521_ & (\all_features[3243]  | \all_features[3244]  | \all_features[3245]  | \all_features[3246]  | \all_features[3247] );
  assign new_n10521_ = ~new_n10512_ & (new_n10511_ | (~new_n10509_ & (new_n10496_ | (~new_n10506_ & ~new_n10522_))));
  assign new_n10522_ = ~new_n10494_ & (new_n10498_ | (new_n10507_ & (~new_n10501_ | (~new_n10523_ & new_n10504_))));
  assign new_n10523_ = ~\all_features[3245]  & \all_features[3246]  & \all_features[3247]  & (\all_features[3244]  ? new_n10502_ : (new_n10500_ | ~new_n10502_));
  assign new_n10524_ = new_n10525_ & new_n10526_;
  assign new_n10525_ = new_n9584_ & new_n9606_;
  assign new_n10526_ = new_n10527_ & new_n10531_;
  assign new_n10527_ = ~new_n10528_ & (\all_features[2627]  | \all_features[2628]  | \all_features[2629]  | \all_features[2630]  | \all_features[2631] );
  assign new_n10528_ = ~new_n9587_ & (new_n9590_ | (~new_n9591_ & (new_n9600_ | (~new_n9595_ & ~new_n10529_))));
  assign new_n10529_ = ~new_n9597_ & (new_n9599_ | (new_n9605_ & (~new_n9601_ | (~new_n10530_ & new_n9603_))));
  assign new_n10530_ = ~\all_features[2629]  & \all_features[2630]  & \all_features[2631]  & (\all_features[2628]  ? new_n9602_ : (new_n9593_ | ~new_n9602_));
  assign new_n10531_ = new_n9586_ & (new_n9591_ | new_n9590_ | (~new_n9595_ & ~new_n9600_ & ~new_n10532_));
  assign new_n10532_ = ~new_n9599_ & ~new_n9597_ & (~new_n9605_ | ~new_n9601_ | new_n10533_);
  assign new_n10533_ = new_n9603_ & new_n9604_ & (new_n10534_ | ~\all_features[2629]  | ~\all_features[2630]  | ~\all_features[2631] );
  assign new_n10534_ = ~\all_features[2627]  & ~\all_features[2628]  & (~\all_features[2626]  | new_n9588_);
  assign new_n10535_ = (~new_n10536_ | new_n10538_) & (~new_n10537_ | (new_n10573_ ? new_n10608_ : ~new_n10610_));
  assign new_n10536_ = new_n10438_ & new_n10378_ & new_n10398_;
  assign new_n10537_ = ~new_n10378_ & ~new_n8892_;
  assign new_n10538_ = new_n10539_ & ~new_n10565_ & ~new_n10569_;
  assign new_n10539_ = ~new_n10540_ & ~new_n10562_;
  assign new_n10540_ = new_n10557_ & ~new_n10561_ & ~new_n10541_ & ~new_n10560_;
  assign new_n10541_ = new_n10542_ & ~new_n10550_ & (~new_n10555_ | ~new_n10556_ | ~new_n10552_ | ~new_n10554_);
  assign new_n10542_ = ~new_n10547_ & ~new_n10543_ & ~new_n10545_;
  assign new_n10543_ = ~\all_features[2655]  & (~\all_features[2654]  | (~\all_features[2652]  & ~\all_features[2653]  & ~new_n10544_));
  assign new_n10544_ = \all_features[2650]  & \all_features[2651] ;
  assign new_n10545_ = ~new_n10546_ & ~\all_features[2655] ;
  assign new_n10546_ = \all_features[2653]  & \all_features[2654]  & (\all_features[2652]  | (\all_features[2650]  & \all_features[2651]  & \all_features[2649] ));
  assign new_n10547_ = ~\all_features[2655]  & (~\all_features[2654]  | ~new_n10548_ | ~new_n10549_ | ~new_n10544_);
  assign new_n10548_ = \all_features[2648]  & \all_features[2649] ;
  assign new_n10549_ = \all_features[2652]  & \all_features[2653] ;
  assign new_n10550_ = ~\all_features[2655]  & (~\all_features[2654]  | (~\all_features[2653]  & (new_n10551_ | ~new_n10544_ | ~\all_features[2652] )));
  assign new_n10551_ = ~\all_features[2648]  & ~\all_features[2649] ;
  assign new_n10552_ = \all_features[2655]  & (\all_features[2654]  | (\all_features[2653]  & (\all_features[2652]  | ~new_n10553_ | ~new_n10551_)));
  assign new_n10553_ = ~\all_features[2650]  & ~\all_features[2651] ;
  assign new_n10554_ = \all_features[2655]  & (\all_features[2654]  | (new_n10549_ & (\all_features[2650]  | \all_features[2651]  | \all_features[2649] )));
  assign new_n10555_ = \all_features[2654]  & \all_features[2655]  & (\all_features[2652]  | \all_features[2653]  | new_n10548_ | ~new_n10553_);
  assign new_n10556_ = \all_features[2655]  & (\all_features[2653]  | \all_features[2654]  | \all_features[2652] );
  assign new_n10557_ = ~new_n10558_ & (\all_features[2651]  | \all_features[2652]  | \all_features[2653]  | \all_features[2654]  | \all_features[2655] );
  assign new_n10558_ = new_n10559_ & (~\all_features[2651]  | ~new_n10549_ | (~\all_features[2650]  & ~new_n10548_));
  assign new_n10559_ = ~\all_features[2654]  & ~\all_features[2655] ;
  assign new_n10560_ = ~\all_features[2653]  & new_n10559_ & ((~\all_features[2650]  & new_n10551_) | ~\all_features[2652]  | ~\all_features[2651] );
  assign new_n10561_ = new_n10559_ & (~\all_features[2653]  | (~\all_features[2652]  & (~\all_features[2651]  | (~\all_features[2650]  & ~\all_features[2649] ))));
  assign new_n10562_ = new_n10542_ & new_n10564_ & ~new_n10550_ & new_n10563_;
  assign new_n10563_ = ~new_n10560_ & (\all_features[2651]  | \all_features[2652]  | \all_features[2653]  | \all_features[2654]  | \all_features[2655] );
  assign new_n10564_ = ~new_n10561_ & ~new_n10558_;
  assign new_n10565_ = ~new_n10566_ & (\all_features[2651]  | \all_features[2652]  | \all_features[2653]  | \all_features[2654]  | \all_features[2655] );
  assign new_n10566_ = ~new_n10560_ & (new_n10561_ | (~new_n10558_ & (new_n10543_ | (~new_n10567_ & ~new_n10550_))));
  assign new_n10567_ = ~new_n10545_ & (new_n10547_ | (new_n10556_ & (~new_n10552_ | (~new_n10568_ & new_n10554_))));
  assign new_n10568_ = ~\all_features[2653]  & \all_features[2654]  & \all_features[2655]  & (\all_features[2652]  ? new_n10553_ : (new_n10548_ | ~new_n10553_));
  assign new_n10569_ = new_n10563_ & (~new_n10564_ | (~new_n10570_ & ~new_n10543_ & ~new_n10550_));
  assign new_n10570_ = ~new_n10545_ & ~new_n10547_ & (~new_n10556_ | ~new_n10552_ | new_n10571_);
  assign new_n10571_ = new_n10554_ & new_n10555_ & (new_n10572_ | ~\all_features[2653]  | ~\all_features[2654]  | ~\all_features[2655] );
  assign new_n10572_ = ~\all_features[2651]  & ~\all_features[2652]  & (~\all_features[2650]  | new_n10551_);
  assign new_n10573_ = new_n10574_ & new_n10603_;
  assign new_n10574_ = new_n10575_ & new_n10596_;
  assign new_n10575_ = ~new_n10576_ & (\all_features[1883]  | \all_features[1884]  | \all_features[1885]  | \all_features[1886]  | \all_features[1887] );
  assign new_n10576_ = ~new_n10590_ & (new_n10592_ | (~new_n10593_ & (new_n10594_ | (~new_n10577_ & ~new_n10595_))));
  assign new_n10577_ = ~new_n10578_ & (new_n10587_ | (new_n10589_ & (~new_n10580_ | (~new_n10585_ & new_n10583_))));
  assign new_n10578_ = ~new_n10579_ & ~\all_features[1887] ;
  assign new_n10579_ = \all_features[1885]  & \all_features[1886]  & (\all_features[1884]  | (\all_features[1882]  & \all_features[1883]  & \all_features[1881] ));
  assign new_n10580_ = \all_features[1887]  & (\all_features[1886]  | (\all_features[1885]  & (\all_features[1884]  | ~new_n10582_ | ~new_n10581_)));
  assign new_n10581_ = ~\all_features[1880]  & ~\all_features[1881] ;
  assign new_n10582_ = ~\all_features[1882]  & ~\all_features[1883] ;
  assign new_n10583_ = \all_features[1887]  & (\all_features[1886]  | (new_n10584_ & (\all_features[1882]  | \all_features[1883]  | \all_features[1881] )));
  assign new_n10584_ = \all_features[1884]  & \all_features[1885] ;
  assign new_n10585_ = ~\all_features[1885]  & \all_features[1886]  & \all_features[1887]  & (\all_features[1884]  ? new_n10582_ : (new_n10586_ | ~new_n10582_));
  assign new_n10586_ = \all_features[1880]  & \all_features[1881] ;
  assign new_n10587_ = ~\all_features[1887]  & (~\all_features[1886]  | ~new_n10586_ | ~new_n10584_ | ~new_n10588_);
  assign new_n10588_ = \all_features[1882]  & \all_features[1883] ;
  assign new_n10589_ = \all_features[1887]  & (\all_features[1885]  | \all_features[1886]  | \all_features[1884] );
  assign new_n10590_ = ~\all_features[1885]  & new_n10591_ & ((~\all_features[1882]  & new_n10581_) | ~\all_features[1884]  | ~\all_features[1883] );
  assign new_n10591_ = ~\all_features[1886]  & ~\all_features[1887] ;
  assign new_n10592_ = new_n10591_ & (~\all_features[1885]  | (~\all_features[1884]  & (~\all_features[1883]  | (~\all_features[1882]  & ~\all_features[1881] ))));
  assign new_n10593_ = new_n10591_ & (~\all_features[1883]  | ~new_n10584_ | (~\all_features[1882]  & ~new_n10586_));
  assign new_n10594_ = ~\all_features[1887]  & (~\all_features[1886]  | (~\all_features[1884]  & ~\all_features[1885]  & ~new_n10588_));
  assign new_n10595_ = ~\all_features[1887]  & (~\all_features[1886]  | (~\all_features[1885]  & (new_n10581_ | ~new_n10588_ | ~\all_features[1884] )));
  assign new_n10596_ = new_n10602_ & (~new_n10601_ | (~new_n10597_ & ~new_n10594_ & ~new_n10595_));
  assign new_n10597_ = ~new_n10587_ & ~new_n10578_ & (~new_n10589_ | ~new_n10580_ | new_n10598_);
  assign new_n10598_ = new_n10583_ & new_n10599_ & (new_n10600_ | ~\all_features[1885]  | ~\all_features[1886]  | ~\all_features[1887] );
  assign new_n10599_ = \all_features[1886]  & \all_features[1887]  & (\all_features[1884]  | \all_features[1885]  | new_n10586_ | ~new_n10582_);
  assign new_n10600_ = ~\all_features[1883]  & ~\all_features[1884]  & (~\all_features[1882]  | new_n10581_);
  assign new_n10601_ = ~new_n10592_ & ~new_n10593_;
  assign new_n10602_ = ~new_n10590_ & (\all_features[1883]  | \all_features[1884]  | \all_features[1885]  | \all_features[1886]  | \all_features[1887] );
  assign new_n10603_ = new_n10604_ & new_n10607_;
  assign new_n10604_ = new_n10601_ & new_n10602_ & (new_n10605_ | new_n10595_ | new_n10587_ | ~new_n10606_);
  assign new_n10605_ = new_n10589_ & new_n10599_ & new_n10580_ & new_n10583_;
  assign new_n10606_ = ~new_n10594_ & ~new_n10578_;
  assign new_n10607_ = new_n10602_ & new_n10601_ & new_n10606_ & ~new_n10595_ & ~new_n10587_;
  assign new_n10608_ = new_n7101_ & (new_n7098_ | ~new_n10609_);
  assign new_n10609_ = ~new_n7068_ & ~new_n7089_;
  assign new_n10610_ = new_n10611_ & new_n10634_;
  assign new_n10611_ = new_n10629_ & ~new_n10633_ & ~new_n10612_ & ~new_n10632_;
  assign new_n10612_ = ~new_n10627_ & ~new_n10628_ & new_n10620_ & (~new_n10625_ | ~new_n10613_);
  assign new_n10613_ = new_n10619_ & new_n10614_ & new_n10616_;
  assign new_n10614_ = \all_features[3415]  & (\all_features[3414]  | (new_n10615_ & (\all_features[3410]  | \all_features[3411]  | \all_features[3409] )));
  assign new_n10615_ = \all_features[3412]  & \all_features[3413] ;
  assign new_n10616_ = \all_features[3414]  & \all_features[3415]  & (\all_features[3412]  | \all_features[3413]  | new_n10618_ | ~new_n10617_);
  assign new_n10617_ = ~\all_features[3410]  & ~\all_features[3411] ;
  assign new_n10618_ = \all_features[3408]  & \all_features[3409] ;
  assign new_n10619_ = \all_features[3415]  & (\all_features[3413]  | \all_features[3414]  | \all_features[3412] );
  assign new_n10620_ = ~new_n10621_ & ~new_n10623_;
  assign new_n10621_ = ~new_n10622_ & ~\all_features[3415] ;
  assign new_n10622_ = \all_features[3413]  & \all_features[3414]  & (\all_features[3412]  | (\all_features[3410]  & \all_features[3411]  & \all_features[3409] ));
  assign new_n10623_ = ~\all_features[3415]  & (~\all_features[3414]  | (~\all_features[3412]  & ~\all_features[3413]  & ~new_n10624_));
  assign new_n10624_ = \all_features[3410]  & \all_features[3411] ;
  assign new_n10625_ = \all_features[3415]  & (\all_features[3414]  | (\all_features[3413]  & (\all_features[3412]  | ~new_n10626_ | ~new_n10617_)));
  assign new_n10626_ = ~\all_features[3408]  & ~\all_features[3409] ;
  assign new_n10627_ = ~\all_features[3415]  & (~\all_features[3414]  | (~\all_features[3413]  & (new_n10626_ | ~new_n10624_ | ~\all_features[3412] )));
  assign new_n10628_ = ~\all_features[3415]  & (~\all_features[3414]  | ~new_n10615_ | ~new_n10618_ | ~new_n10624_);
  assign new_n10629_ = ~new_n10630_ & (\all_features[3411]  | \all_features[3412]  | \all_features[3413]  | \all_features[3414]  | \all_features[3415] );
  assign new_n10630_ = ~\all_features[3413]  & new_n10631_ & ((~\all_features[3410]  & new_n10626_) | ~\all_features[3412]  | ~\all_features[3411] );
  assign new_n10631_ = ~\all_features[3414]  & ~\all_features[3415] ;
  assign new_n10632_ = new_n10631_ & (~\all_features[3413]  | (~\all_features[3412]  & (~\all_features[3411]  | (~\all_features[3410]  & ~\all_features[3409] ))));
  assign new_n10633_ = new_n10631_ & (~\all_features[3411]  | ~new_n10615_ | (~\all_features[3410]  & ~new_n10618_));
  assign new_n10634_ = new_n10629_ & new_n10620_ & new_n10635_ & ~new_n10627_ & ~new_n10628_;
  assign new_n10635_ = ~new_n10632_ & ~new_n10633_;
  assign new_n10636_ = new_n10407_ & ~new_n10398_ & new_n10378_;
  assign new_n10637_ = ~new_n9867_ & ~new_n9864_;
  assign new_n10638_ = new_n10639_ & new_n10640_;
  assign new_n10639_ = (~new_n10636_ | new_n10637_) & (~new_n10377_ | (new_n10454_ ? new_n10524_ : new_n10489_));
  assign new_n10640_ = (~new_n10538_ | ~new_n10536_) & (~new_n10537_ | (new_n10573_ ? ~new_n10608_ : new_n10610_));
  assign new_n10641_ = new_n10772_ & ~new_n10642_ & ~new_n10699_;
  assign new_n10642_ = ~new_n10643_ & (new_n10682_ ? (new_n10647_ ? ~new_n10645_ : new_n7602_) : ~new_n10681_);
  assign new_n10643_ = ~new_n10644_ & new_n6384_;
  assign new_n10644_ = new_n6356_ & new_n6378_;
  assign new_n10645_ = new_n9720_ & new_n10646_;
  assign new_n10646_ = ~new_n9691_ & ~new_n9712_;
  assign new_n10647_ = ~new_n10677_ & (~new_n10679_ | new_n10648_);
  assign new_n10648_ = ~new_n10649_ & ~new_n10670_;
  assign new_n10649_ = ~new_n10650_ & (\all_features[3899]  | \all_features[3900]  | \all_features[3901]  | \all_features[3902]  | \all_features[3903] );
  assign new_n10650_ = ~new_n10666_ & (new_n10664_ | (~new_n10668_ & (new_n10669_ | (~new_n10667_ & ~new_n10651_))));
  assign new_n10651_ = ~new_n10652_ & (new_n10654_ | (new_n10663_ & (~new_n10658_ | (~new_n10662_ & new_n10661_))));
  assign new_n10652_ = ~new_n10653_ & ~\all_features[3903] ;
  assign new_n10653_ = \all_features[3901]  & \all_features[3902]  & (\all_features[3900]  | (\all_features[3898]  & \all_features[3899]  & \all_features[3897] ));
  assign new_n10654_ = ~\all_features[3903]  & (~\all_features[3902]  | ~new_n10655_ | ~new_n10656_ | ~new_n10657_);
  assign new_n10655_ = \all_features[3898]  & \all_features[3899] ;
  assign new_n10656_ = \all_features[3896]  & \all_features[3897] ;
  assign new_n10657_ = \all_features[3900]  & \all_features[3901] ;
  assign new_n10658_ = \all_features[3903]  & (\all_features[3902]  | (\all_features[3901]  & (\all_features[3900]  | ~new_n10660_ | ~new_n10659_)));
  assign new_n10659_ = ~\all_features[3896]  & ~\all_features[3897] ;
  assign new_n10660_ = ~\all_features[3898]  & ~\all_features[3899] ;
  assign new_n10661_ = \all_features[3903]  & (\all_features[3902]  | (new_n10657_ & (\all_features[3898]  | \all_features[3899]  | \all_features[3897] )));
  assign new_n10662_ = ~\all_features[3901]  & \all_features[3902]  & \all_features[3903]  & (\all_features[3900]  ? new_n10660_ : (new_n10656_ | ~new_n10660_));
  assign new_n10663_ = \all_features[3903]  & (\all_features[3901]  | \all_features[3902]  | \all_features[3900] );
  assign new_n10664_ = new_n10665_ & (~\all_features[3901]  | (~\all_features[3900]  & (~\all_features[3899]  | (~\all_features[3898]  & ~\all_features[3897] ))));
  assign new_n10665_ = ~\all_features[3902]  & ~\all_features[3903] ;
  assign new_n10666_ = ~\all_features[3901]  & new_n10665_ & ((~\all_features[3898]  & new_n10659_) | ~\all_features[3900]  | ~\all_features[3899] );
  assign new_n10667_ = ~\all_features[3903]  & (~\all_features[3902]  | (~\all_features[3901]  & (new_n10659_ | ~new_n10655_ | ~\all_features[3900] )));
  assign new_n10668_ = new_n10665_ & (~\all_features[3899]  | ~new_n10657_ | (~\all_features[3898]  & ~new_n10656_));
  assign new_n10669_ = ~\all_features[3903]  & (~\all_features[3902]  | (~\all_features[3900]  & ~\all_features[3901]  & ~new_n10655_));
  assign new_n10670_ = new_n10675_ & (~new_n10676_ | (~new_n10671_ & ~new_n10667_ & ~new_n10669_));
  assign new_n10671_ = ~new_n10652_ & ~new_n10654_ & (~new_n10663_ | ~new_n10658_ | new_n10672_);
  assign new_n10672_ = new_n10661_ & new_n10673_ & (new_n10674_ | ~\all_features[3901]  | ~\all_features[3902]  | ~\all_features[3903] );
  assign new_n10673_ = \all_features[3902]  & \all_features[3903]  & (\all_features[3900]  | \all_features[3901]  | new_n10656_ | ~new_n10660_);
  assign new_n10674_ = ~\all_features[3899]  & ~\all_features[3900]  & (~\all_features[3898]  | new_n10659_);
  assign new_n10675_ = ~new_n10666_ & (\all_features[3899]  | \all_features[3900]  | \all_features[3901]  | \all_features[3902]  | \all_features[3903] );
  assign new_n10676_ = ~new_n10664_ & ~new_n10668_;
  assign new_n10677_ = new_n10678_ & new_n10675_ & ~new_n10668_ & ~new_n10667_ & ~new_n10652_ & ~new_n10664_;
  assign new_n10678_ = ~new_n10654_ & ~new_n10669_;
  assign new_n10679_ = new_n10675_ & new_n10676_ & (new_n10680_ | new_n10652_ | new_n10667_ | ~new_n10678_);
  assign new_n10680_ = new_n10663_ & new_n10673_ & new_n10658_ & new_n10661_;
  assign new_n10681_ = ~new_n9129_ & ~new_n9131_;
  assign new_n10682_ = new_n10694_ & new_n10686_ & ~new_n10698_ & ~new_n10697_ & ~new_n10683_ & ~new_n10692_;
  assign new_n10683_ = ~\all_features[2383]  & (~\all_features[2382]  | new_n10684_);
  assign new_n10684_ = ~\all_features[2381]  & (new_n10685_ | ~\all_features[2379]  | ~\all_features[2380]  | ~\all_features[2378] );
  assign new_n10685_ = ~\all_features[2376]  & ~\all_features[2377] ;
  assign new_n10686_ = ~new_n10687_ & ~new_n10691_;
  assign new_n10687_ = new_n10688_ & (~\all_features[2379]  | ~new_n10690_ | (~\all_features[2378]  & ~new_n10689_));
  assign new_n10688_ = ~\all_features[2382]  & ~\all_features[2383] ;
  assign new_n10689_ = \all_features[2376]  & \all_features[2377] ;
  assign new_n10690_ = \all_features[2380]  & \all_features[2381] ;
  assign new_n10691_ = new_n10688_ & (~\all_features[2381]  | (~\all_features[2380]  & (~\all_features[2379]  | (~\all_features[2378]  & ~\all_features[2377] ))));
  assign new_n10692_ = ~new_n10693_ & ~\all_features[2383] ;
  assign new_n10693_ = \all_features[2381]  & \all_features[2382]  & (\all_features[2380]  | (\all_features[2378]  & \all_features[2379]  & \all_features[2377] ));
  assign new_n10694_ = ~new_n10695_ & ~new_n10696_;
  assign new_n10695_ = ~\all_features[2383]  & ~\all_features[2382]  & ~\all_features[2381]  & ~\all_features[2379]  & ~\all_features[2380] ;
  assign new_n10696_ = ~\all_features[2383]  & (~\all_features[2382]  | (~\all_features[2381]  & ~\all_features[2380]  & (~\all_features[2379]  | ~\all_features[2378] )));
  assign new_n10697_ = ~\all_features[2381]  & new_n10688_ & ((~\all_features[2378]  & new_n10685_) | ~\all_features[2380]  | ~\all_features[2379] );
  assign new_n10698_ = ~\all_features[2383]  & (~new_n10690_ | ~\all_features[2378]  | ~\all_features[2379]  | ~\all_features[2382]  | ~new_n10689_);
  assign new_n10699_ = new_n10737_ & new_n10643_ & (new_n10700_ ? ~new_n10701_ : ~new_n10771_);
  assign new_n10700_ = ~new_n7101_ & (~new_n7098_ | ~new_n7067_);
  assign new_n10701_ = new_n10702_ & new_n10728_;
  assign new_n10702_ = ~new_n10703_ & ~new_n10726_;
  assign new_n10703_ = new_n10721_ & ~new_n10725_ & ~new_n10704_ & ~new_n10724_;
  assign new_n10704_ = ~new_n10719_ & ~new_n10720_ & new_n10712_ & (~new_n10717_ | ~new_n10705_);
  assign new_n10705_ = new_n10711_ & new_n10706_ & new_n10708_;
  assign new_n10706_ = \all_features[1479]  & (\all_features[1478]  | (new_n10707_ & (\all_features[1474]  | \all_features[1475]  | \all_features[1473] )));
  assign new_n10707_ = \all_features[1476]  & \all_features[1477] ;
  assign new_n10708_ = \all_features[1478]  & \all_features[1479]  & (\all_features[1476]  | \all_features[1477]  | new_n10710_ | ~new_n10709_);
  assign new_n10709_ = ~\all_features[1474]  & ~\all_features[1475] ;
  assign new_n10710_ = \all_features[1472]  & \all_features[1473] ;
  assign new_n10711_ = \all_features[1479]  & (\all_features[1477]  | \all_features[1478]  | \all_features[1476] );
  assign new_n10712_ = ~new_n10713_ & ~new_n10715_;
  assign new_n10713_ = ~new_n10714_ & ~\all_features[1479] ;
  assign new_n10714_ = \all_features[1477]  & \all_features[1478]  & (\all_features[1476]  | (\all_features[1474]  & \all_features[1475]  & \all_features[1473] ));
  assign new_n10715_ = ~\all_features[1479]  & (~\all_features[1478]  | (~\all_features[1476]  & ~\all_features[1477]  & ~new_n10716_));
  assign new_n10716_ = \all_features[1474]  & \all_features[1475] ;
  assign new_n10717_ = \all_features[1479]  & (\all_features[1478]  | (\all_features[1477]  & (\all_features[1476]  | ~new_n10718_ | ~new_n10709_)));
  assign new_n10718_ = ~\all_features[1472]  & ~\all_features[1473] ;
  assign new_n10719_ = ~\all_features[1479]  & (~\all_features[1478]  | (~\all_features[1477]  & (new_n10718_ | ~new_n10716_ | ~\all_features[1476] )));
  assign new_n10720_ = ~\all_features[1479]  & (~\all_features[1478]  | ~new_n10707_ | ~new_n10710_ | ~new_n10716_);
  assign new_n10721_ = ~new_n10722_ & (\all_features[1475]  | \all_features[1476]  | \all_features[1477]  | \all_features[1478]  | \all_features[1479] );
  assign new_n10722_ = ~\all_features[1477]  & new_n10723_ & ((~\all_features[1474]  & new_n10718_) | ~\all_features[1476]  | ~\all_features[1475] );
  assign new_n10723_ = ~\all_features[1478]  & ~\all_features[1479] ;
  assign new_n10724_ = new_n10723_ & (~\all_features[1477]  | (~\all_features[1476]  & (~\all_features[1475]  | (~\all_features[1474]  & ~\all_features[1473] ))));
  assign new_n10725_ = new_n10723_ & (~\all_features[1475]  | ~new_n10707_ | (~\all_features[1474]  & ~new_n10710_));
  assign new_n10726_ = new_n10721_ & new_n10712_ & new_n10727_ & ~new_n10719_ & ~new_n10720_;
  assign new_n10727_ = ~new_n10724_ & ~new_n10725_;
  assign new_n10728_ = ~new_n10729_ & ~new_n10733_;
  assign new_n10729_ = new_n10721_ & (~new_n10727_ | (~new_n10730_ & ~new_n10715_ & ~new_n10719_));
  assign new_n10730_ = ~new_n10720_ & ~new_n10713_ & (~new_n10711_ | ~new_n10717_ | new_n10731_);
  assign new_n10731_ = new_n10706_ & new_n10708_ & (new_n10732_ | ~\all_features[1477]  | ~\all_features[1478]  | ~\all_features[1479] );
  assign new_n10732_ = ~\all_features[1475]  & ~\all_features[1476]  & (~\all_features[1474]  | new_n10718_);
  assign new_n10733_ = ~new_n10734_ & (\all_features[1475]  | \all_features[1476]  | \all_features[1477]  | \all_features[1478]  | \all_features[1479] );
  assign new_n10734_ = ~new_n10722_ & (new_n10724_ | (~new_n10725_ & (new_n10715_ | (~new_n10719_ & ~new_n10735_))));
  assign new_n10735_ = ~new_n10713_ & (new_n10720_ | (new_n10711_ & (~new_n10717_ | (~new_n10736_ & new_n10706_))));
  assign new_n10736_ = ~\all_features[1477]  & \all_features[1478]  & \all_features[1479]  & (\all_features[1476]  ? new_n10709_ : (new_n10710_ | ~new_n10709_));
  assign new_n10737_ = new_n10738_ & new_n10762_;
  assign new_n10738_ = ~new_n10739_ & ~new_n10761_;
  assign new_n10739_ = new_n10740_ & (~new_n10749_ | (new_n10759_ & new_n10760_ & new_n10756_ & new_n10758_));
  assign new_n10740_ = new_n10741_ & ~new_n10745_ & ~new_n10746_;
  assign new_n10741_ = ~new_n10742_ & (\all_features[1947]  | \all_features[1948]  | \all_features[1949]  | \all_features[1950]  | \all_features[1951] );
  assign new_n10742_ = ~\all_features[1949]  & new_n10744_ & ((~\all_features[1946]  & new_n10743_) | ~\all_features[1948]  | ~\all_features[1947] );
  assign new_n10743_ = ~\all_features[1944]  & ~\all_features[1945] ;
  assign new_n10744_ = ~\all_features[1950]  & ~\all_features[1951] ;
  assign new_n10745_ = new_n10744_ & (~\all_features[1949]  | (~\all_features[1948]  & (~\all_features[1947]  | (~\all_features[1946]  & ~\all_features[1945] ))));
  assign new_n10746_ = new_n10744_ & (~\all_features[1947]  | ~new_n10747_ | (~\all_features[1946]  & ~new_n10748_));
  assign new_n10747_ = \all_features[1948]  & \all_features[1949] ;
  assign new_n10748_ = \all_features[1944]  & \all_features[1945] ;
  assign new_n10749_ = ~new_n10755_ & ~new_n10754_ & ~new_n10750_ & ~new_n10752_;
  assign new_n10750_ = ~\all_features[1951]  & (~\all_features[1950]  | (~\all_features[1949]  & (new_n10743_ | ~new_n10751_ | ~\all_features[1948] )));
  assign new_n10751_ = \all_features[1946]  & \all_features[1947] ;
  assign new_n10752_ = ~new_n10753_ & ~\all_features[1951] ;
  assign new_n10753_ = \all_features[1949]  & \all_features[1950]  & (\all_features[1948]  | (\all_features[1946]  & \all_features[1947]  & \all_features[1945] ));
  assign new_n10754_ = ~\all_features[1951]  & (~\all_features[1950]  | ~new_n10747_ | ~new_n10748_ | ~new_n10751_);
  assign new_n10755_ = ~\all_features[1951]  & (~\all_features[1950]  | (~\all_features[1948]  & ~\all_features[1949]  & ~new_n10751_));
  assign new_n10756_ = \all_features[1951]  & (\all_features[1950]  | (\all_features[1949]  & (\all_features[1948]  | ~new_n10743_ | ~new_n10757_)));
  assign new_n10757_ = ~\all_features[1946]  & ~\all_features[1947] ;
  assign new_n10758_ = \all_features[1951]  & (\all_features[1950]  | (new_n10747_ & (\all_features[1946]  | \all_features[1947]  | \all_features[1945] )));
  assign new_n10759_ = \all_features[1950]  & \all_features[1951]  & (\all_features[1948]  | \all_features[1949]  | new_n10748_ | ~new_n10757_);
  assign new_n10760_ = \all_features[1951]  & (\all_features[1949]  | \all_features[1950]  | \all_features[1948] );
  assign new_n10761_ = new_n10740_ & new_n10749_;
  assign new_n10762_ = ~new_n10763_ & ~new_n10767_;
  assign new_n10763_ = ~new_n10764_ & (\all_features[1947]  | \all_features[1948]  | \all_features[1949]  | \all_features[1950]  | \all_features[1951] );
  assign new_n10764_ = ~new_n10742_ & (new_n10745_ | (~new_n10746_ & (new_n10755_ | (~new_n10750_ & ~new_n10765_))));
  assign new_n10765_ = ~new_n10752_ & (new_n10754_ | (new_n10760_ & (~new_n10756_ | (~new_n10766_ & new_n10758_))));
  assign new_n10766_ = ~\all_features[1949]  & \all_features[1950]  & \all_features[1951]  & (\all_features[1948]  ? new_n10757_ : (new_n10748_ | ~new_n10757_));
  assign new_n10767_ = new_n10741_ & (new_n10746_ | new_n10745_ | (~new_n10750_ & ~new_n10755_ & ~new_n10768_));
  assign new_n10768_ = ~new_n10754_ & ~new_n10752_ & (~new_n10760_ | ~new_n10756_ | new_n10769_);
  assign new_n10769_ = new_n10758_ & new_n10759_ & (new_n10770_ | ~\all_features[1949]  | ~\all_features[1950]  | ~\all_features[1951] );
  assign new_n10770_ = ~\all_features[1947]  & ~\all_features[1948]  & (~\all_features[1946]  | new_n10743_);
  assign new_n10771_ = new_n8739_ & (new_n8736_ | new_n8725_);
  assign new_n10772_ = (~new_n10777_ | new_n10737_ | ~new_n10643_) & (new_n10682_ | ~new_n10681_ | ~new_n10773_ | new_n10643_);
  assign new_n10773_ = ~new_n10775_ & (~new_n10776_ | ~new_n10774_);
  assign new_n10774_ = new_n8299_ & new_n8320_;
  assign new_n10775_ = new_n8344_ & new_n8346_;
  assign new_n10776_ = ~new_n8346_ & new_n8344_;
  assign new_n10777_ = new_n10805_ & new_n10830_ & new_n10833_ & new_n10834_ & (new_n10801_ | new_n10778_);
  assign new_n10778_ = new_n10798_ & ~new_n10779_ & new_n10793_;
  assign new_n10779_ = ~new_n10787_ & ~new_n10789_ & ~new_n10791_ & ~new_n10792_ & (~new_n10783_ | ~new_n10780_);
  assign new_n10780_ = \all_features[4391]  & (\all_features[4390]  | (~new_n10781_ & \all_features[4389] ));
  assign new_n10781_ = new_n10782_ & ~\all_features[4388]  & ~\all_features[4386]  & ~\all_features[4387] ;
  assign new_n10782_ = ~\all_features[4384]  & ~\all_features[4385] ;
  assign new_n10783_ = \all_features[4391]  & \all_features[4390]  & ~new_n10786_ & new_n10784_;
  assign new_n10784_ = \all_features[4391]  & (\all_features[4390]  | (new_n10785_ & (\all_features[4386]  | \all_features[4387]  | \all_features[4385] )));
  assign new_n10785_ = \all_features[4388]  & \all_features[4389] ;
  assign new_n10786_ = ~\all_features[4386]  & ~\all_features[4387]  & ~\all_features[4388]  & ~\all_features[4389]  & (~\all_features[4385]  | ~\all_features[4384] );
  assign new_n10787_ = ~\all_features[4391]  & (~\all_features[4390]  | (~\all_features[4389]  & (new_n10782_ | ~new_n10788_ | ~\all_features[4388] )));
  assign new_n10788_ = \all_features[4386]  & \all_features[4387] ;
  assign new_n10789_ = ~new_n10790_ & ~\all_features[4391] ;
  assign new_n10790_ = \all_features[4389]  & \all_features[4390]  & (\all_features[4388]  | (\all_features[4386]  & \all_features[4387]  & \all_features[4385] ));
  assign new_n10791_ = ~\all_features[4391]  & (~\all_features[4390]  | (~\all_features[4388]  & ~\all_features[4389]  & ~new_n10788_));
  assign new_n10792_ = ~\all_features[4391]  & (~new_n10788_ | ~\all_features[4384]  | ~\all_features[4385]  | ~\all_features[4390]  | ~new_n10785_);
  assign new_n10793_ = ~new_n10794_ & ~new_n10797_;
  assign new_n10794_ = new_n10795_ & ~\all_features[4387]  & ~\all_features[4388] ;
  assign new_n10795_ = ~\all_features[4389]  & new_n10796_;
  assign new_n10796_ = ~\all_features[4390]  & ~\all_features[4391] ;
  assign new_n10797_ = new_n10795_ & ((~\all_features[4386]  & new_n10782_) | ~\all_features[4388]  | ~\all_features[4387] );
  assign new_n10798_ = ~new_n10799_ & ~new_n10800_;
  assign new_n10799_ = new_n10796_ & (~new_n10785_ | ~\all_features[4387]  | (~\all_features[4386]  & (~\all_features[4384]  | ~\all_features[4385] )));
  assign new_n10800_ = new_n10796_ & (~\all_features[4389]  | (~\all_features[4388]  & (~\all_features[4387]  | (~\all_features[4386]  & ~\all_features[4385] ))));
  assign new_n10801_ = new_n10793_ & (~new_n10798_ | (new_n10804_ & (new_n10802_ | new_n10789_ | new_n10792_)));
  assign new_n10802_ = new_n10780_ & (~new_n10783_ | (~new_n10803_ & \all_features[4389]  & \all_features[4390]  & \all_features[4391] ));
  assign new_n10803_ = ~\all_features[4387]  & ~\all_features[4388]  & (~\all_features[4386]  | new_n10782_);
  assign new_n10804_ = ~new_n10787_ & ~new_n10791_;
  assign new_n10805_ = new_n10828_ & (~new_n10816_ | (new_n10820_ & (~new_n10824_ | new_n10806_)));
  assign new_n10806_ = new_n10807_ & (~new_n10810_ | (~new_n10815_ & \all_features[1661]  & \all_features[1662]  & \all_features[1663] ));
  assign new_n10807_ = \all_features[1663]  & (\all_features[1662]  | (~new_n10808_ & \all_features[1661] ));
  assign new_n10808_ = new_n10809_ & ~\all_features[1660]  & ~\all_features[1658]  & ~\all_features[1659] ;
  assign new_n10809_ = ~\all_features[1656]  & ~\all_features[1657] ;
  assign new_n10810_ = \all_features[1663]  & \all_features[1662]  & ~new_n10813_ & new_n10811_;
  assign new_n10811_ = \all_features[1663]  & (\all_features[1662]  | (new_n10812_ & (\all_features[1658]  | \all_features[1659]  | \all_features[1657] )));
  assign new_n10812_ = \all_features[1660]  & \all_features[1661] ;
  assign new_n10813_ = ~\all_features[1661]  & ~\all_features[1660]  & ~\all_features[1659]  & ~new_n10814_ & ~\all_features[1658] ;
  assign new_n10814_ = \all_features[1656]  & \all_features[1657] ;
  assign new_n10815_ = ~\all_features[1659]  & ~\all_features[1660]  & (~\all_features[1658]  | new_n10809_);
  assign new_n10816_ = ~new_n10817_ & ~new_n10818_;
  assign new_n10817_ = ~\all_features[1662]  & ~\all_features[1663]  & (~\all_features[1659]  | ~new_n10812_ | (~\all_features[1658]  & ~new_n10814_));
  assign new_n10818_ = ~\all_features[1663]  & ~new_n10819_ & ~\all_features[1662] ;
  assign new_n10819_ = \all_features[1661]  & (\all_features[1660]  | (\all_features[1659]  & (\all_features[1658]  | \all_features[1657] )));
  assign new_n10820_ = ~new_n10821_ & ~new_n10823_;
  assign new_n10821_ = ~\all_features[1663]  & (~\all_features[1662]  | (~\all_features[1660]  & ~\all_features[1661]  & ~new_n10822_));
  assign new_n10822_ = \all_features[1658]  & \all_features[1659] ;
  assign new_n10823_ = ~\all_features[1663]  & (~\all_features[1662]  | (~\all_features[1661]  & (new_n10809_ | ~new_n10822_ | ~\all_features[1660] )));
  assign new_n10824_ = ~new_n10825_ & ~new_n10826_;
  assign new_n10825_ = ~\all_features[1663]  & (~\all_features[1662]  | ~new_n10814_ | ~new_n10812_ | ~new_n10822_);
  assign new_n10826_ = ~new_n10827_ & ~\all_features[1663] ;
  assign new_n10827_ = \all_features[1661]  & \all_features[1662]  & (\all_features[1660]  | (\all_features[1658]  & \all_features[1659]  & \all_features[1657] ));
  assign new_n10828_ = ~new_n10829_ | (\all_features[1659]  & \all_features[1660]  & (\all_features[1658]  | ~new_n10809_));
  assign new_n10829_ = ~\all_features[1663]  & ~\all_features[1661]  & ~\all_features[1662] ;
  assign new_n10830_ = new_n10831_ & (new_n10823_ | new_n10826_ | ~new_n10832_ | (new_n10810_ & new_n10807_));
  assign new_n10831_ = new_n10816_ & new_n10828_;
  assign new_n10832_ = ~new_n10821_ & ~new_n10825_;
  assign new_n10833_ = new_n10824_ & new_n10831_ & new_n10820_;
  assign new_n10834_ = new_n10804_ & new_n10798_ & ~new_n10792_ & ~new_n10789_ & ~new_n10794_ & ~new_n10797_;
  assign new_n10835_ = new_n10836_ & (new_n10910_ | ((new_n10976_ | ~new_n11095_ | ~new_n10837_) & (new_n11024_ | new_n10837_)));
  assign new_n10836_ = (~new_n10910_ | (new_n10947_ ? new_n11023_ : new_n10872_)) & (~new_n10975_ | ~new_n10837_ | new_n10910_);
  assign new_n10837_ = ~new_n10838_ & ~new_n10871_;
  assign new_n10838_ = ~new_n10839_ & new_n10868_;
  assign new_n10839_ = ~new_n10840_ & ~new_n10861_;
  assign new_n10840_ = ~new_n10841_ & (\all_features[2763]  | \all_features[2764]  | \all_features[2765]  | \all_features[2766]  | \all_features[2767] );
  assign new_n10841_ = ~new_n10857_ & (new_n10855_ | (~new_n10859_ & (new_n10860_ | (~new_n10858_ & ~new_n10842_))));
  assign new_n10842_ = ~new_n10843_ & (new_n10845_ | (new_n10854_ & (~new_n10849_ | (~new_n10853_ & new_n10852_))));
  assign new_n10843_ = ~new_n10844_ & ~\all_features[2767] ;
  assign new_n10844_ = \all_features[2765]  & \all_features[2766]  & (\all_features[2764]  | (\all_features[2762]  & \all_features[2763]  & \all_features[2761] ));
  assign new_n10845_ = ~\all_features[2767]  & (~\all_features[2766]  | ~new_n10846_ | ~new_n10847_ | ~new_n10848_);
  assign new_n10846_ = \all_features[2762]  & \all_features[2763] ;
  assign new_n10847_ = \all_features[2760]  & \all_features[2761] ;
  assign new_n10848_ = \all_features[2764]  & \all_features[2765] ;
  assign new_n10849_ = \all_features[2767]  & (\all_features[2766]  | (\all_features[2765]  & (\all_features[2764]  | ~new_n10851_ | ~new_n10850_)));
  assign new_n10850_ = ~\all_features[2760]  & ~\all_features[2761] ;
  assign new_n10851_ = ~\all_features[2762]  & ~\all_features[2763] ;
  assign new_n10852_ = \all_features[2767]  & (\all_features[2766]  | (new_n10848_ & (\all_features[2762]  | \all_features[2763]  | \all_features[2761] )));
  assign new_n10853_ = ~\all_features[2765]  & \all_features[2766]  & \all_features[2767]  & (\all_features[2764]  ? new_n10851_ : (new_n10847_ | ~new_n10851_));
  assign new_n10854_ = \all_features[2767]  & (\all_features[2765]  | \all_features[2766]  | \all_features[2764] );
  assign new_n10855_ = new_n10856_ & (~\all_features[2765]  | (~\all_features[2764]  & (~\all_features[2763]  | (~\all_features[2762]  & ~\all_features[2761] ))));
  assign new_n10856_ = ~\all_features[2766]  & ~\all_features[2767] ;
  assign new_n10857_ = ~\all_features[2765]  & new_n10856_ & ((~\all_features[2762]  & new_n10850_) | ~\all_features[2764]  | ~\all_features[2763] );
  assign new_n10858_ = ~\all_features[2767]  & (~\all_features[2766]  | (~\all_features[2765]  & (new_n10850_ | ~new_n10846_ | ~\all_features[2764] )));
  assign new_n10859_ = new_n10856_ & (~\all_features[2763]  | ~new_n10848_ | (~\all_features[2762]  & ~new_n10847_));
  assign new_n10860_ = ~\all_features[2767]  & (~\all_features[2766]  | (~\all_features[2764]  & ~\all_features[2765]  & ~new_n10846_));
  assign new_n10861_ = new_n10866_ & (~new_n10867_ | (~new_n10862_ & ~new_n10858_ & ~new_n10860_));
  assign new_n10862_ = ~new_n10843_ & ~new_n10845_ & (~new_n10854_ | ~new_n10849_ | new_n10863_);
  assign new_n10863_ = new_n10852_ & new_n10864_ & (new_n10865_ | ~\all_features[2765]  | ~\all_features[2766]  | ~\all_features[2767] );
  assign new_n10864_ = \all_features[2766]  & \all_features[2767]  & (\all_features[2764]  | \all_features[2765]  | new_n10847_ | ~new_n10851_);
  assign new_n10865_ = ~\all_features[2763]  & ~\all_features[2764]  & (~\all_features[2762]  | new_n10850_);
  assign new_n10866_ = ~new_n10857_ & (\all_features[2763]  | \all_features[2764]  | \all_features[2765]  | \all_features[2766]  | \all_features[2767] );
  assign new_n10867_ = ~new_n10855_ & ~new_n10859_;
  assign new_n10868_ = new_n10866_ & new_n10867_ & (new_n10870_ | new_n10843_ | new_n10858_ | ~new_n10869_);
  assign new_n10869_ = ~new_n10845_ & ~new_n10860_;
  assign new_n10870_ = new_n10854_ & new_n10864_ & new_n10849_ & new_n10852_;
  assign new_n10871_ = new_n10869_ & new_n10866_ & ~new_n10859_ & ~new_n10858_ & ~new_n10843_ & ~new_n10855_;
  assign new_n10872_ = (~new_n10906_ & new_n10873_ & (~new_n10908_ | new_n10877_)) | (~new_n10876_ & new_n8662_ & ~new_n10873_);
  assign new_n10873_ = ~new_n10874_ & new_n10875_;
  assign new_n10874_ = ~new_n8357_ & ~new_n8381_;
  assign new_n10875_ = new_n8385_ & new_n8388_;
  assign new_n10876_ = ~new_n8632_ & ~new_n8652_;
  assign new_n10877_ = ~new_n10878_ & ~new_n10899_;
  assign new_n10878_ = ~new_n10879_ & (\all_features[2611]  | \all_features[2612]  | \all_features[2613]  | \all_features[2614]  | \all_features[2615] );
  assign new_n10879_ = ~new_n10895_ & (new_n10893_ | (~new_n10897_ & (new_n10898_ | (~new_n10896_ & ~new_n10880_))));
  assign new_n10880_ = ~new_n10881_ & (new_n10883_ | (new_n10892_ & (~new_n10887_ | (~new_n10891_ & new_n10890_))));
  assign new_n10881_ = ~new_n10882_ & ~\all_features[2615] ;
  assign new_n10882_ = \all_features[2613]  & \all_features[2614]  & (\all_features[2612]  | (\all_features[2610]  & \all_features[2611]  & \all_features[2609] ));
  assign new_n10883_ = ~\all_features[2615]  & (~\all_features[2614]  | ~new_n10884_ | ~new_n10885_ | ~new_n10886_);
  assign new_n10884_ = \all_features[2610]  & \all_features[2611] ;
  assign new_n10885_ = \all_features[2608]  & \all_features[2609] ;
  assign new_n10886_ = \all_features[2612]  & \all_features[2613] ;
  assign new_n10887_ = \all_features[2615]  & (\all_features[2614]  | (\all_features[2613]  & (\all_features[2612]  | ~new_n10889_ | ~new_n10888_)));
  assign new_n10888_ = ~\all_features[2608]  & ~\all_features[2609] ;
  assign new_n10889_ = ~\all_features[2610]  & ~\all_features[2611] ;
  assign new_n10890_ = \all_features[2615]  & (\all_features[2614]  | (new_n10886_ & (\all_features[2610]  | \all_features[2611]  | \all_features[2609] )));
  assign new_n10891_ = ~\all_features[2613]  & \all_features[2614]  & \all_features[2615]  & (\all_features[2612]  ? new_n10889_ : (new_n10885_ | ~new_n10889_));
  assign new_n10892_ = \all_features[2615]  & (\all_features[2613]  | \all_features[2614]  | \all_features[2612] );
  assign new_n10893_ = new_n10894_ & (~\all_features[2613]  | (~\all_features[2612]  & (~\all_features[2611]  | (~\all_features[2610]  & ~\all_features[2609] ))));
  assign new_n10894_ = ~\all_features[2614]  & ~\all_features[2615] ;
  assign new_n10895_ = ~\all_features[2613]  & new_n10894_ & ((~\all_features[2610]  & new_n10888_) | ~\all_features[2612]  | ~\all_features[2611] );
  assign new_n10896_ = ~\all_features[2615]  & (~\all_features[2614]  | (~\all_features[2613]  & (new_n10888_ | ~new_n10884_ | ~\all_features[2612] )));
  assign new_n10897_ = new_n10894_ & (~\all_features[2611]  | ~new_n10886_ | (~\all_features[2610]  & ~new_n10885_));
  assign new_n10898_ = ~\all_features[2615]  & (~\all_features[2614]  | (~\all_features[2612]  & ~\all_features[2613]  & ~new_n10884_));
  assign new_n10899_ = new_n10904_ & (~new_n10905_ | (~new_n10900_ & ~new_n10896_ & ~new_n10898_));
  assign new_n10900_ = ~new_n10881_ & ~new_n10883_ & (~new_n10892_ | ~new_n10887_ | new_n10901_);
  assign new_n10901_ = new_n10890_ & new_n10902_ & (new_n10903_ | ~\all_features[2613]  | ~\all_features[2614]  | ~\all_features[2615] );
  assign new_n10902_ = \all_features[2614]  & \all_features[2615]  & (\all_features[2612]  | \all_features[2613]  | new_n10885_ | ~new_n10889_);
  assign new_n10903_ = ~\all_features[2611]  & ~\all_features[2612]  & (~\all_features[2610]  | new_n10888_);
  assign new_n10904_ = ~new_n10895_ & (\all_features[2611]  | \all_features[2612]  | \all_features[2613]  | \all_features[2614]  | \all_features[2615] );
  assign new_n10905_ = ~new_n10893_ & ~new_n10897_;
  assign new_n10906_ = new_n10907_ & new_n10904_ & ~new_n10897_ & ~new_n10896_ & ~new_n10881_ & ~new_n10893_;
  assign new_n10907_ = ~new_n10883_ & ~new_n10898_;
  assign new_n10908_ = new_n10904_ & new_n10905_ & (new_n10909_ | new_n10881_ | new_n10896_ | ~new_n10907_);
  assign new_n10909_ = new_n10892_ & new_n10902_ & new_n10887_ & new_n10890_;
  assign new_n10910_ = new_n10911_ & new_n10938_;
  assign new_n10911_ = ~new_n10912_ & ~new_n10936_;
  assign new_n10912_ = new_n10930_ & ~new_n10935_ & ~new_n10913_ & ~new_n10934_;
  assign new_n10913_ = new_n10914_ & new_n10921_ & (~new_n10928_ | ~new_n10929_ | ~new_n10925_ | ~new_n10927_);
  assign new_n10914_ = ~new_n10915_ & ~new_n10919_;
  assign new_n10915_ = ~\all_features[4567]  & (~\all_features[4566]  | ~new_n10916_ | ~new_n10917_ | ~new_n10918_);
  assign new_n10916_ = \all_features[4564]  & \all_features[4565] ;
  assign new_n10917_ = \all_features[4560]  & \all_features[4561] ;
  assign new_n10918_ = \all_features[4562]  & \all_features[4563] ;
  assign new_n10919_ = ~new_n10920_ & ~\all_features[4567] ;
  assign new_n10920_ = \all_features[4565]  & \all_features[4566]  & (\all_features[4564]  | (\all_features[4562]  & \all_features[4563]  & \all_features[4561] ));
  assign new_n10921_ = ~new_n10922_ & ~new_n10924_;
  assign new_n10922_ = ~\all_features[4567]  & (~\all_features[4566]  | (~\all_features[4565]  & (new_n10923_ | ~new_n10918_ | ~\all_features[4564] )));
  assign new_n10923_ = ~\all_features[4560]  & ~\all_features[4561] ;
  assign new_n10924_ = ~\all_features[4567]  & (~\all_features[4566]  | (~\all_features[4564]  & ~\all_features[4565]  & ~new_n10918_));
  assign new_n10925_ = \all_features[4567]  & (\all_features[4566]  | (\all_features[4565]  & (\all_features[4564]  | ~new_n10923_ | ~new_n10926_)));
  assign new_n10926_ = ~\all_features[4562]  & ~\all_features[4563] ;
  assign new_n10927_ = \all_features[4567]  & (\all_features[4566]  | (new_n10916_ & (\all_features[4562]  | \all_features[4563]  | \all_features[4561] )));
  assign new_n10928_ = \all_features[4566]  & \all_features[4567]  & (\all_features[4564]  | \all_features[4565]  | new_n10917_ | ~new_n10926_);
  assign new_n10929_ = \all_features[4567]  & (\all_features[4565]  | \all_features[4566]  | \all_features[4564] );
  assign new_n10930_ = ~new_n10931_ & ~new_n10933_;
  assign new_n10931_ = ~\all_features[4565]  & new_n10932_ & ((~\all_features[4562]  & new_n10923_) | ~\all_features[4564]  | ~\all_features[4563] );
  assign new_n10932_ = ~\all_features[4566]  & ~\all_features[4567] ;
  assign new_n10933_ = ~\all_features[4567]  & ~\all_features[4566]  & ~\all_features[4565]  & ~\all_features[4563]  & ~\all_features[4564] ;
  assign new_n10934_ = new_n10932_ & (~\all_features[4565]  | (~\all_features[4564]  & (~\all_features[4563]  | (~\all_features[4562]  & ~\all_features[4561] ))));
  assign new_n10935_ = new_n10932_ & (~\all_features[4563]  | ~new_n10916_ | (~\all_features[4562]  & ~new_n10917_));
  assign new_n10936_ = new_n10937_ & new_n10930_ & new_n10914_ & new_n10921_;
  assign new_n10937_ = ~new_n10934_ & ~new_n10935_;
  assign new_n10938_ = ~new_n10939_ & ~new_n10943_;
  assign new_n10939_ = new_n10930_ & (~new_n10937_ | (~new_n10940_ & new_n10921_));
  assign new_n10940_ = new_n10914_ & ((~new_n10941_ & new_n10927_ & new_n10928_) | ~new_n10929_ | ~new_n10925_);
  assign new_n10941_ = \all_features[4567]  & \all_features[4566]  & ~new_n10942_ & \all_features[4565] ;
  assign new_n10942_ = ~\all_features[4563]  & ~\all_features[4564]  & (~\all_features[4562]  | new_n10923_);
  assign new_n10943_ = ~new_n10933_ & (new_n10931_ | new_n10944_);
  assign new_n10944_ = ~new_n10934_ & (new_n10935_ | (~new_n10924_ & (new_n10922_ | (~new_n10919_ & ~new_n10945_))));
  assign new_n10945_ = ~new_n10915_ & (~new_n10929_ | (new_n10925_ & (~new_n10927_ | (~new_n10946_ & new_n10928_))));
  assign new_n10946_ = \all_features[4566]  & \all_features[4567]  & (\all_features[4565]  | (~new_n10926_ & \all_features[4564] ));
  assign new_n10947_ = new_n10948_ & new_n10972_;
  assign new_n10948_ = new_n10949_ & new_n10970_;
  assign new_n10949_ = new_n10967_ & ~new_n10950_ & new_n10964_;
  assign new_n10950_ = ~new_n10958_ & ~new_n10960_ & ~new_n10962_ & ~new_n10963_ & (~new_n10954_ | ~new_n10951_);
  assign new_n10951_ = \all_features[1903]  & (\all_features[1902]  | (~new_n10952_ & \all_features[1901] ));
  assign new_n10952_ = new_n10953_ & ~\all_features[1900]  & ~\all_features[1898]  & ~\all_features[1899] ;
  assign new_n10953_ = ~\all_features[1896]  & ~\all_features[1897] ;
  assign new_n10954_ = \all_features[1903]  & \all_features[1902]  & ~new_n10957_ & new_n10955_;
  assign new_n10955_ = \all_features[1903]  & (\all_features[1902]  | (new_n10956_ & (\all_features[1898]  | \all_features[1899]  | \all_features[1897] )));
  assign new_n10956_ = \all_features[1900]  & \all_features[1901] ;
  assign new_n10957_ = ~\all_features[1898]  & ~\all_features[1899]  & ~\all_features[1900]  & ~\all_features[1901]  & (~\all_features[1897]  | ~\all_features[1896] );
  assign new_n10958_ = ~\all_features[1903]  & (~\all_features[1902]  | (~\all_features[1901]  & (new_n10953_ | ~new_n10959_ | ~\all_features[1900] )));
  assign new_n10959_ = \all_features[1898]  & \all_features[1899] ;
  assign new_n10960_ = ~new_n10961_ & ~\all_features[1903] ;
  assign new_n10961_ = \all_features[1901]  & \all_features[1902]  & (\all_features[1900]  | (\all_features[1898]  & \all_features[1899]  & \all_features[1897] ));
  assign new_n10962_ = ~\all_features[1903]  & (~new_n10959_ | ~\all_features[1896]  | ~\all_features[1897]  | ~\all_features[1902]  | ~new_n10956_);
  assign new_n10963_ = ~\all_features[1903]  & (~\all_features[1902]  | (~\all_features[1900]  & ~\all_features[1901]  & ~new_n10959_));
  assign new_n10964_ = ~new_n10965_ | (\all_features[1899]  & \all_features[1900]  & (\all_features[1898]  | ~new_n10953_));
  assign new_n10965_ = ~\all_features[1901]  & new_n10966_;
  assign new_n10966_ = ~\all_features[1902]  & ~\all_features[1903] ;
  assign new_n10967_ = ~new_n10968_ & ~new_n10969_;
  assign new_n10968_ = new_n10966_ & (~new_n10956_ | ~\all_features[1899]  | (~\all_features[1898]  & (~\all_features[1896]  | ~\all_features[1897] )));
  assign new_n10969_ = new_n10966_ & (~\all_features[1901]  | (~\all_features[1900]  & (~\all_features[1899]  | (~\all_features[1898]  & ~\all_features[1897] ))));
  assign new_n10970_ = new_n10967_ & new_n10964_ & new_n10971_ & ~new_n10960_ & ~new_n10962_;
  assign new_n10971_ = ~new_n10958_ & ~new_n10963_;
  assign new_n10972_ = new_n10964_ & (~new_n10967_ | (new_n10971_ & (new_n10973_ | new_n10960_ | new_n10962_)));
  assign new_n10973_ = new_n10951_ & (~new_n10954_ | (~new_n10974_ & \all_features[1901]  & \all_features[1902]  & \all_features[1903] ));
  assign new_n10974_ = ~\all_features[1899]  & ~\all_features[1900]  & (~\all_features[1898]  | new_n10953_);
  assign new_n10975_ = new_n10976_ & (~new_n11016_ | ~new_n11000_);
  assign new_n10976_ = ~new_n10977_ & ~new_n10999_;
  assign new_n10977_ = new_n10978_ & (~new_n10987_ | (new_n10997_ & new_n10998_ & new_n10994_ & new_n10996_));
  assign new_n10978_ = new_n10979_ & ~new_n10983_ & ~new_n10984_;
  assign new_n10979_ = ~new_n10980_ & (\all_features[3451]  | \all_features[3452]  | \all_features[3453]  | \all_features[3454]  | \all_features[3455] );
  assign new_n10980_ = ~\all_features[3453]  & new_n10982_ & ((~\all_features[3450]  & new_n10981_) | ~\all_features[3452]  | ~\all_features[3451] );
  assign new_n10981_ = ~\all_features[3448]  & ~\all_features[3449] ;
  assign new_n10982_ = ~\all_features[3454]  & ~\all_features[3455] ;
  assign new_n10983_ = new_n10982_ & (~\all_features[3453]  | (~\all_features[3452]  & (~\all_features[3451]  | (~\all_features[3450]  & ~\all_features[3449] ))));
  assign new_n10984_ = new_n10982_ & (~\all_features[3451]  | ~new_n10985_ | (~\all_features[3450]  & ~new_n10986_));
  assign new_n10985_ = \all_features[3452]  & \all_features[3453] ;
  assign new_n10986_ = \all_features[3448]  & \all_features[3449] ;
  assign new_n10987_ = ~new_n10993_ & ~new_n10992_ & ~new_n10988_ & ~new_n10990_;
  assign new_n10988_ = ~\all_features[3455]  & (~\all_features[3454]  | (~\all_features[3453]  & (new_n10981_ | ~new_n10989_ | ~\all_features[3452] )));
  assign new_n10989_ = \all_features[3450]  & \all_features[3451] ;
  assign new_n10990_ = ~new_n10991_ & ~\all_features[3455] ;
  assign new_n10991_ = \all_features[3453]  & \all_features[3454]  & (\all_features[3452]  | (\all_features[3450]  & \all_features[3451]  & \all_features[3449] ));
  assign new_n10992_ = ~\all_features[3455]  & (~\all_features[3454]  | ~new_n10985_ | ~new_n10986_ | ~new_n10989_);
  assign new_n10993_ = ~\all_features[3455]  & (~\all_features[3454]  | (~\all_features[3452]  & ~\all_features[3453]  & ~new_n10989_));
  assign new_n10994_ = \all_features[3455]  & (\all_features[3454]  | (\all_features[3453]  & (\all_features[3452]  | ~new_n10981_ | ~new_n10995_)));
  assign new_n10995_ = ~\all_features[3450]  & ~\all_features[3451] ;
  assign new_n10996_ = \all_features[3455]  & (\all_features[3454]  | (new_n10985_ & (\all_features[3450]  | \all_features[3451]  | \all_features[3449] )));
  assign new_n10997_ = \all_features[3454]  & \all_features[3455]  & (\all_features[3452]  | \all_features[3453]  | new_n10986_ | ~new_n10995_);
  assign new_n10998_ = \all_features[3455]  & (\all_features[3453]  | \all_features[3454]  | \all_features[3452] );
  assign new_n10999_ = new_n10978_ & new_n10987_;
  assign new_n11000_ = new_n11001_ & new_n11010_;
  assign new_n11001_ = ~new_n11009_ & ~new_n11007_ & ~new_n11002_ & ~new_n11005_;
  assign new_n11002_ = ~\all_features[2743]  & (~\all_features[2742]  | (~\all_features[2741]  & (new_n11004_ | ~\all_features[2740]  | ~new_n11003_)));
  assign new_n11003_ = \all_features[2738]  & \all_features[2739] ;
  assign new_n11004_ = ~\all_features[2736]  & ~\all_features[2737] ;
  assign new_n11005_ = ~new_n11006_ & ~\all_features[2743] ;
  assign new_n11006_ = \all_features[2741]  & \all_features[2742]  & (\all_features[2740]  | (\all_features[2738]  & \all_features[2739]  & \all_features[2737] ));
  assign new_n11007_ = ~\all_features[2743]  & (~new_n11008_ | ~\all_features[2736]  | ~\all_features[2737]  | ~\all_features[2742]  | ~new_n11003_);
  assign new_n11008_ = \all_features[2740]  & \all_features[2741] ;
  assign new_n11009_ = ~\all_features[2743]  & (~\all_features[2742]  | (~\all_features[2740]  & ~\all_features[2741]  & ~new_n11003_));
  assign new_n11010_ = ~new_n11015_ & ~new_n11014_ & ~new_n11011_ & ~new_n11013_;
  assign new_n11011_ = new_n11012_ & (~\all_features[2741]  | (~\all_features[2740]  & (~\all_features[2739]  | (~\all_features[2738]  & ~\all_features[2737] ))));
  assign new_n11012_ = ~\all_features[2742]  & ~\all_features[2743] ;
  assign new_n11013_ = new_n11012_ & (~new_n11008_ | ~\all_features[2739]  | (~\all_features[2738]  & (~\all_features[2736]  | ~\all_features[2737] )));
  assign new_n11014_ = ~\all_features[2741]  & new_n11012_ & ((~\all_features[2738]  & new_n11004_) | ~\all_features[2740]  | ~\all_features[2739] );
  assign new_n11015_ = ~\all_features[2743]  & ~\all_features[2742]  & ~\all_features[2741]  & ~\all_features[2739]  & ~\all_features[2740] ;
  assign new_n11016_ = new_n11010_ & (~new_n11001_ | (new_n11020_ & new_n11022_ & new_n11017_ & new_n11019_));
  assign new_n11017_ = \all_features[2743]  & (\all_features[2742]  | (\all_features[2741]  & (\all_features[2740]  | ~new_n11018_ | ~new_n11004_)));
  assign new_n11018_ = ~\all_features[2738]  & ~\all_features[2739] ;
  assign new_n11019_ = \all_features[2743]  & (\all_features[2742]  | (new_n11008_ & (\all_features[2738]  | \all_features[2739]  | \all_features[2737] )));
  assign new_n11020_ = new_n11021_ & (\all_features[2740]  | \all_features[2741]  | ~new_n11018_ | (\all_features[2737]  & \all_features[2736] ));
  assign new_n11021_ = \all_features[2742]  & \all_features[2743] ;
  assign new_n11022_ = \all_features[2743]  & (\all_features[2741]  | \all_features[2742]  | \all_features[2740] );
  assign new_n11023_ = ~new_n8701_ & (~new_n8698_ | new_n8668_);
  assign new_n11024_ = (new_n11060_ | ~new_n11025_) & (~new_n11062_ | ~new_n11094_ | new_n11025_);
  assign new_n11025_ = new_n11059_ & (new_n11055_ | ~new_n11026_);
  assign new_n11026_ = ~new_n11027_ & ~new_n11051_;
  assign new_n11027_ = ~new_n11049_ & ~new_n11048_ & (~new_n11042_ | (~new_n11028_ & ~new_n11046_ & ~new_n11050_));
  assign new_n11028_ = ~new_n11037_ & ~new_n11038_ & (~new_n11041_ | ~new_n11040_ | new_n11029_);
  assign new_n11029_ = new_n11030_ & new_n11032_ & (new_n11035_ | ~\all_features[5461]  | ~\all_features[5462]  | ~\all_features[5463] );
  assign new_n11030_ = \all_features[5463]  & (\all_features[5462]  | (new_n11031_ & (\all_features[5458]  | \all_features[5459]  | \all_features[5457] )));
  assign new_n11031_ = \all_features[5460]  & \all_features[5461] ;
  assign new_n11032_ = \all_features[5462]  & \all_features[5463]  & (\all_features[5460]  | \all_features[5461]  | new_n11033_ | ~new_n11034_);
  assign new_n11033_ = \all_features[5456]  & \all_features[5457] ;
  assign new_n11034_ = ~\all_features[5458]  & ~\all_features[5459] ;
  assign new_n11035_ = ~\all_features[5459]  & ~\all_features[5460]  & (~\all_features[5458]  | new_n11036_);
  assign new_n11036_ = ~\all_features[5456]  & ~\all_features[5457] ;
  assign new_n11037_ = ~\all_features[5463]  & (~new_n11031_ | ~\all_features[5458]  | ~\all_features[5459]  | ~\all_features[5462]  | ~new_n11033_);
  assign new_n11038_ = ~new_n11039_ & ~\all_features[5463] ;
  assign new_n11039_ = \all_features[5461]  & \all_features[5462]  & (\all_features[5460]  | (\all_features[5458]  & \all_features[5459]  & \all_features[5457] ));
  assign new_n11040_ = \all_features[5463]  & (\all_features[5462]  | (\all_features[5461]  & (\all_features[5460]  | ~new_n11034_ | ~new_n11036_)));
  assign new_n11041_ = \all_features[5463]  & (\all_features[5461]  | \all_features[5462]  | \all_features[5460] );
  assign new_n11042_ = ~new_n11043_ & ~new_n11045_;
  assign new_n11043_ = new_n11044_ & (~\all_features[5459]  | ~new_n11031_ | (~\all_features[5458]  & ~new_n11033_));
  assign new_n11044_ = ~\all_features[5462]  & ~\all_features[5463] ;
  assign new_n11045_ = new_n11044_ & (~\all_features[5461]  | (~\all_features[5460]  & (~\all_features[5459]  | (~\all_features[5458]  & ~\all_features[5457] ))));
  assign new_n11046_ = ~\all_features[5463]  & (~\all_features[5462]  | new_n11047_);
  assign new_n11047_ = ~\all_features[5461]  & (new_n11036_ | ~\all_features[5459]  | ~\all_features[5460]  | ~\all_features[5458] );
  assign new_n11048_ = ~\all_features[5461]  & new_n11044_ & ((~\all_features[5458]  & new_n11036_) | ~\all_features[5460]  | ~\all_features[5459] );
  assign new_n11049_ = ~\all_features[5463]  & ~\all_features[5462]  & ~\all_features[5461]  & ~\all_features[5459]  & ~\all_features[5460] ;
  assign new_n11050_ = ~\all_features[5463]  & (~\all_features[5462]  | (~\all_features[5461]  & ~\all_features[5460]  & (~\all_features[5459]  | ~\all_features[5458] )));
  assign new_n11051_ = ~new_n11052_ & ~new_n11049_;
  assign new_n11052_ = ~new_n11048_ & (new_n11045_ | (~new_n11043_ & (new_n11050_ | (~new_n11046_ & ~new_n11053_))));
  assign new_n11053_ = ~new_n11038_ & (new_n11037_ | (new_n11041_ & (~new_n11040_ | (~new_n11054_ & new_n11030_))));
  assign new_n11054_ = ~\all_features[5461]  & \all_features[5462]  & \all_features[5463]  & (\all_features[5460]  ? new_n11034_ : (new_n11033_ | ~new_n11034_));
  assign new_n11055_ = ~new_n11049_ & ~new_n11048_ & ~new_n11045_ & ~new_n11056_ & ~new_n11043_;
  assign new_n11056_ = ~new_n11046_ & ~new_n11037_ & new_n11057_ & (~new_n11040_ | ~new_n11058_);
  assign new_n11057_ = ~new_n11038_ & ~new_n11050_;
  assign new_n11058_ = new_n11041_ & new_n11030_ & new_n11032_;
  assign new_n11059_ = new_n11042_ & new_n11057_ & ~new_n11049_ & ~new_n11037_ & ~new_n11046_ & ~new_n11048_;
  assign new_n11060_ = ~new_n11061_ & new_n6568_;
  assign new_n11061_ = ~new_n6593_ & ~new_n6597_;
  assign new_n11062_ = new_n11092_ & (new_n11083_ | new_n11063_);
  assign new_n11063_ = ~new_n11082_ & (new_n11081_ | (~new_n11080_ & (new_n11078_ | (~new_n11077_ & ~new_n11064_))));
  assign new_n11064_ = ~new_n11071_ & (new_n11073_ | (~new_n11075_ & (~new_n11076_ | new_n11065_)));
  assign new_n11065_ = \all_features[1207]  & ((~new_n11070_ & ~\all_features[1205]  & \all_features[1206] ) | (~new_n11068_ & (\all_features[1206]  | (~new_n11066_ & \all_features[1205] ))));
  assign new_n11066_ = new_n11067_ & ~\all_features[1204]  & ~\all_features[1202]  & ~\all_features[1203] ;
  assign new_n11067_ = ~\all_features[1200]  & ~\all_features[1201] ;
  assign new_n11068_ = \all_features[1207]  & (\all_features[1206]  | (new_n11069_ & (\all_features[1202]  | \all_features[1203]  | \all_features[1201] )));
  assign new_n11069_ = \all_features[1204]  & \all_features[1205] ;
  assign new_n11070_ = (~\all_features[1202]  & ~\all_features[1203]  & ~\all_features[1204]  & (~\all_features[1201]  | ~\all_features[1200] )) | (\all_features[1204]  & (\all_features[1202]  | \all_features[1203] ));
  assign new_n11071_ = ~\all_features[1207]  & (~\all_features[1206]  | (~\all_features[1205]  & (new_n11067_ | ~\all_features[1204]  | ~new_n11072_)));
  assign new_n11072_ = \all_features[1202]  & \all_features[1203] ;
  assign new_n11073_ = ~new_n11074_ & ~\all_features[1207] ;
  assign new_n11074_ = \all_features[1205]  & \all_features[1206]  & (\all_features[1204]  | (\all_features[1202]  & \all_features[1203]  & \all_features[1201] ));
  assign new_n11075_ = ~\all_features[1207]  & (~new_n11069_ | ~\all_features[1200]  | ~\all_features[1201]  | ~\all_features[1206]  | ~new_n11072_);
  assign new_n11076_ = \all_features[1207]  & (\all_features[1205]  | \all_features[1206]  | \all_features[1204] );
  assign new_n11077_ = ~\all_features[1207]  & (~\all_features[1206]  | (~\all_features[1204]  & ~\all_features[1205]  & ~new_n11072_));
  assign new_n11078_ = new_n11079_ & (~new_n11069_ | ~\all_features[1203]  | (~\all_features[1202]  & (~\all_features[1200]  | ~\all_features[1201] )));
  assign new_n11079_ = ~\all_features[1206]  & ~\all_features[1207] ;
  assign new_n11080_ = new_n11079_ & (~\all_features[1205]  | (~\all_features[1204]  & (~\all_features[1203]  | (~\all_features[1202]  & ~\all_features[1201] ))));
  assign new_n11081_ = ~\all_features[1205]  & new_n11079_ & ((~\all_features[1202]  & new_n11067_) | ~\all_features[1204]  | ~\all_features[1203] );
  assign new_n11082_ = ~\all_features[1207]  & ~\all_features[1206]  & ~\all_features[1205]  & ~\all_features[1203]  & ~\all_features[1204] ;
  assign new_n11083_ = new_n11091_ & (~new_n11090_ | (new_n11089_ & (new_n11084_ | new_n11073_ | new_n11075_)));
  assign new_n11084_ = new_n11085_ & (~new_n11086_ | (~new_n11088_ & \all_features[1205]  & \all_features[1206]  & \all_features[1207] ));
  assign new_n11085_ = \all_features[1207]  & (\all_features[1206]  | (~new_n11066_ & \all_features[1205] ));
  assign new_n11086_ = \all_features[1207]  & \all_features[1206]  & ~new_n11087_ & new_n11068_;
  assign new_n11087_ = ~\all_features[1202]  & ~\all_features[1203]  & ~\all_features[1204]  & ~\all_features[1205]  & (~\all_features[1201]  | ~\all_features[1200] );
  assign new_n11088_ = ~\all_features[1203]  & ~\all_features[1204]  & (~\all_features[1202]  | new_n11067_);
  assign new_n11089_ = ~new_n11071_ & ~new_n11077_;
  assign new_n11090_ = ~new_n11078_ & ~new_n11080_;
  assign new_n11091_ = ~new_n11081_ & ~new_n11082_;
  assign new_n11092_ = new_n11091_ & ~new_n11093_ & new_n11090_;
  assign new_n11093_ = ~new_n11071_ & ~new_n11077_ & ~new_n11073_ & ~new_n11075_ & (~new_n11086_ | ~new_n11085_);
  assign new_n11094_ = new_n11090_ & new_n11089_ & new_n11091_ & ~new_n11073_ & ~new_n11075_;
  assign new_n11095_ = ~new_n11123_ & new_n11096_;
  assign new_n11096_ = ~new_n11097_ & ~new_n11120_;
  assign new_n11097_ = new_n11098_ & (new_n11117_ | new_n11118_ | ~new_n11113_ | (new_n11110_ & new_n11108_));
  assign new_n11098_ = new_n11099_ & new_n11105_;
  assign new_n11099_ = ~new_n11100_ & ~new_n11103_;
  assign new_n11100_ = ~\all_features[3726]  & ~\all_features[3727]  & (~\all_features[3723]  | ~new_n11102_ | (~\all_features[3722]  & ~new_n11101_));
  assign new_n11101_ = \all_features[3720]  & \all_features[3721] ;
  assign new_n11102_ = \all_features[3724]  & \all_features[3725] ;
  assign new_n11103_ = ~\all_features[3727]  & ~new_n11104_ & ~\all_features[3726] ;
  assign new_n11104_ = \all_features[3725]  & (\all_features[3724]  | (\all_features[3723]  & (\all_features[3722]  | \all_features[3721] )));
  assign new_n11105_ = ~new_n11107_ | (\all_features[3723]  & \all_features[3724]  & (\all_features[3722]  | ~new_n11106_));
  assign new_n11106_ = ~\all_features[3720]  & ~\all_features[3721] ;
  assign new_n11107_ = ~\all_features[3727]  & ~\all_features[3725]  & ~\all_features[3726] ;
  assign new_n11108_ = \all_features[3727]  & (\all_features[3726]  | (~new_n11109_ & \all_features[3725] ));
  assign new_n11109_ = new_n11106_ & ~\all_features[3724]  & ~\all_features[3722]  & ~\all_features[3723] ;
  assign new_n11110_ = \all_features[3727]  & \all_features[3726]  & ~new_n11112_ & new_n11111_;
  assign new_n11111_ = \all_features[3727]  & (\all_features[3726]  | (new_n11102_ & (\all_features[3722]  | \all_features[3723]  | \all_features[3721] )));
  assign new_n11112_ = ~\all_features[3725]  & ~\all_features[3724]  & ~\all_features[3723]  & ~new_n11101_ & ~\all_features[3722] ;
  assign new_n11113_ = ~new_n11114_ & ~new_n11116_;
  assign new_n11114_ = ~\all_features[3727]  & (~\all_features[3726]  | (~\all_features[3724]  & ~\all_features[3725]  & ~new_n11115_));
  assign new_n11115_ = \all_features[3722]  & \all_features[3723] ;
  assign new_n11116_ = ~\all_features[3727]  & (~\all_features[3726]  | ~new_n11101_ | ~new_n11102_ | ~new_n11115_);
  assign new_n11117_ = ~\all_features[3727]  & (~\all_features[3726]  | (~\all_features[3725]  & (new_n11106_ | ~new_n11115_ | ~\all_features[3724] )));
  assign new_n11118_ = ~new_n11119_ & ~\all_features[3727] ;
  assign new_n11119_ = \all_features[3725]  & \all_features[3726]  & (\all_features[3724]  | (\all_features[3722]  & \all_features[3723]  & \all_features[3721] ));
  assign new_n11120_ = new_n11122_ & new_n11098_ & new_n11121_;
  assign new_n11121_ = ~new_n11114_ & ~new_n11117_;
  assign new_n11122_ = ~new_n11116_ & ~new_n11118_;
  assign new_n11123_ = new_n11105_ & (~new_n11099_ | (new_n11121_ & (~new_n11122_ | new_n11124_)));
  assign new_n11124_ = new_n11108_ & (~new_n11110_ | (~new_n11125_ & \all_features[3725]  & \all_features[3726]  & \all_features[3727] ));
  assign new_n11125_ = ~\all_features[3723]  & ~\all_features[3724]  & (~\all_features[3722]  | new_n11106_);
  assign new_n11126_ = new_n11127_ ? (new_n11374_ ^ new_n11574_) : (~new_n11374_ ^ new_n11574_);
  assign new_n11127_ = new_n11128_ & (new_n11168_ ? (~new_n7636_ | new_n11302_) : new_n11271_);
  assign new_n11128_ = new_n11129_ & (new_n11202_ | new_n11168_ | new_n11170_ | new_n11238_);
  assign new_n11129_ = ~new_n11165_ & (~new_n11130_ | ~new_n11168_ | new_n11171_ | new_n7636_);
  assign new_n11130_ = new_n11131_ & new_n11160_;
  assign new_n11131_ = ~new_n11132_ & ~new_n11154_;
  assign new_n11132_ = ~new_n11133_ & (\all_features[1515]  | \all_features[1516]  | \all_features[1517]  | \all_features[1518]  | \all_features[1519] );
  assign new_n11133_ = ~new_n11151_ & (new_n11149_ | (~new_n11152_ & (new_n11153_ | (~new_n11134_ & ~new_n11147_))));
  assign new_n11134_ = ~new_n11144_ & (new_n11146_ | new_n11135_);
  assign new_n11135_ = \all_features[1519]  & ((new_n11136_ & (\all_features[1518]  | \all_features[1517] )) | (~\all_features[1518]  & (\all_features[1517]  ? new_n11142_ : \all_features[1516] )));
  assign new_n11136_ = new_n11137_ & (\all_features[1517]  | ~new_n11140_ | (~new_n11141_ & ~\all_features[1516]  & new_n11139_) | (\all_features[1516]  & ~new_n11139_));
  assign new_n11137_ = \all_features[1519]  & (\all_features[1518]  | (new_n11138_ & (\all_features[1514]  | \all_features[1515]  | \all_features[1513] )));
  assign new_n11138_ = \all_features[1516]  & \all_features[1517] ;
  assign new_n11139_ = ~\all_features[1514]  & ~\all_features[1515] ;
  assign new_n11140_ = \all_features[1518]  & \all_features[1519] ;
  assign new_n11141_ = \all_features[1512]  & \all_features[1513] ;
  assign new_n11142_ = new_n11139_ & ~\all_features[1516]  & new_n11143_;
  assign new_n11143_ = ~\all_features[1512]  & ~\all_features[1513] ;
  assign new_n11144_ = ~new_n11145_ & ~\all_features[1519] ;
  assign new_n11145_ = \all_features[1517]  & \all_features[1518]  & (\all_features[1516]  | (\all_features[1514]  & \all_features[1515]  & \all_features[1513] ));
  assign new_n11146_ = ~\all_features[1519]  & (~new_n11138_ | ~\all_features[1514]  | ~\all_features[1515]  | ~\all_features[1518]  | ~new_n11141_);
  assign new_n11147_ = ~\all_features[1519]  & (~\all_features[1518]  | new_n11148_);
  assign new_n11148_ = ~\all_features[1517]  & (new_n11143_ | ~\all_features[1515]  | ~\all_features[1516]  | ~\all_features[1514] );
  assign new_n11149_ = new_n11150_ & (~\all_features[1517]  | (~\all_features[1516]  & (~\all_features[1515]  | (~\all_features[1514]  & ~\all_features[1513] ))));
  assign new_n11150_ = ~\all_features[1518]  & ~\all_features[1519] ;
  assign new_n11151_ = ~\all_features[1517]  & new_n11150_ & ((~\all_features[1514]  & new_n11143_) | ~\all_features[1516]  | ~\all_features[1515] );
  assign new_n11152_ = new_n11150_ & (~\all_features[1515]  | ~new_n11138_ | (~\all_features[1514]  & ~new_n11141_));
  assign new_n11153_ = ~\all_features[1519]  & (~\all_features[1518]  | (~\all_features[1517]  & ~\all_features[1516]  & (~\all_features[1515]  | ~\all_features[1514] )));
  assign new_n11154_ = new_n11159_ & (new_n11152_ | new_n11149_ | (~new_n11155_ & ~new_n11147_ & ~new_n11153_));
  assign new_n11155_ = ~new_n11146_ & ~new_n11144_ & (~new_n11156_ | (~new_n11158_ & new_n11137_ & new_n11157_));
  assign new_n11156_ = \all_features[1519]  & (\all_features[1518]  | (~new_n11142_ & \all_features[1517] ));
  assign new_n11157_ = new_n11140_ & (new_n11141_ | \all_features[1516]  | \all_features[1517]  | ~new_n11139_);
  assign new_n11158_ = new_n11140_ & \all_features[1517]  & ((~new_n11143_ & \all_features[1514] ) | \all_features[1516]  | \all_features[1515] );
  assign new_n11159_ = ~new_n11151_ & (\all_features[1515]  | \all_features[1516]  | \all_features[1517]  | \all_features[1518]  | \all_features[1519] );
  assign new_n11160_ = ~new_n11161_ & ~new_n11164_;
  assign new_n11161_ = new_n11159_ & ~new_n11152_ & ~new_n11162_ & ~new_n11149_;
  assign new_n11162_ = ~new_n11147_ & ~new_n11146_ & new_n11163_ & (~new_n11137_ | ~new_n11157_ | ~new_n11156_);
  assign new_n11163_ = ~new_n11144_ & ~new_n11153_;
  assign new_n11164_ = new_n11163_ & new_n11159_ & ~new_n11152_ & ~new_n11149_ & ~new_n11147_ & ~new_n11146_;
  assign new_n11165_ = new_n11170_ & new_n9652_ & ~new_n11166_ & ~new_n11168_;
  assign new_n11166_ = ~new_n11167_ & new_n8666_;
  assign new_n11167_ = ~new_n8652_ & ~new_n8663_;
  assign new_n11168_ = ~new_n7995_ & new_n11169_;
  assign new_n11169_ = ~new_n8028_ & ~new_n8026_;
  assign new_n11170_ = ~new_n10936_ & (~new_n10939_ | ~new_n10912_);
  assign new_n11171_ = ~new_n11201_ & new_n11172_;
  assign new_n11172_ = ~new_n11173_ & ~new_n11199_;
  assign new_n11173_ = new_n11193_ & (~new_n11189_ | (new_n11185_ & (new_n11174_ | new_n11196_ | new_n11198_)));
  assign new_n11174_ = new_n11175_ & (~new_n11179_ | (~new_n11184_ & \all_features[3437]  & \all_features[3438]  & \all_features[3439] ));
  assign new_n11175_ = \all_features[3439]  & (\all_features[3438]  | (~new_n11176_ & \all_features[3437] ));
  assign new_n11176_ = new_n11177_ & ~\all_features[3436]  & new_n11178_;
  assign new_n11177_ = ~\all_features[3432]  & ~\all_features[3433] ;
  assign new_n11178_ = ~\all_features[3434]  & ~\all_features[3435] ;
  assign new_n11179_ = \all_features[3439]  & \all_features[3438]  & ~new_n11182_ & new_n11180_;
  assign new_n11180_ = \all_features[3439]  & (\all_features[3438]  | (new_n11181_ & (\all_features[3434]  | \all_features[3435]  | \all_features[3433] )));
  assign new_n11181_ = \all_features[3436]  & \all_features[3437] ;
  assign new_n11182_ = new_n11178_ & ~\all_features[3437]  & ~new_n11183_ & ~\all_features[3436] ;
  assign new_n11183_ = \all_features[3432]  & \all_features[3433] ;
  assign new_n11184_ = ~\all_features[3435]  & ~\all_features[3436]  & (~\all_features[3434]  | new_n11177_);
  assign new_n11185_ = ~new_n11186_ & ~new_n11188_;
  assign new_n11186_ = ~\all_features[3439]  & (~\all_features[3438]  | (~\all_features[3436]  & ~\all_features[3437]  & ~new_n11187_));
  assign new_n11187_ = \all_features[3434]  & \all_features[3435] ;
  assign new_n11188_ = ~\all_features[3439]  & (~\all_features[3438]  | (~\all_features[3437]  & (new_n11177_ | ~\all_features[3436]  | ~new_n11187_)));
  assign new_n11189_ = ~new_n11190_ & ~new_n11192_;
  assign new_n11190_ = new_n11191_ & (~\all_features[3435]  | ~new_n11181_ | (~\all_features[3434]  & ~new_n11183_));
  assign new_n11191_ = ~\all_features[3438]  & ~\all_features[3439] ;
  assign new_n11192_ = new_n11191_ & (~\all_features[3437]  | (~\all_features[3436]  & (~\all_features[3435]  | (~\all_features[3434]  & ~\all_features[3433] ))));
  assign new_n11193_ = ~new_n11194_ & ~new_n11195_;
  assign new_n11194_ = ~\all_features[3437]  & new_n11191_ & ((~\all_features[3434]  & new_n11177_) | ~\all_features[3436]  | ~\all_features[3435] );
  assign new_n11195_ = ~\all_features[3439]  & ~\all_features[3438]  & ~\all_features[3437]  & ~\all_features[3435]  & ~\all_features[3436] ;
  assign new_n11196_ = ~new_n11197_ & ~\all_features[3439] ;
  assign new_n11197_ = \all_features[3437]  & \all_features[3438]  & (\all_features[3436]  | (\all_features[3434]  & \all_features[3435]  & \all_features[3433] ));
  assign new_n11198_ = ~\all_features[3439]  & (~\all_features[3438]  | ~new_n11187_ | ~new_n11183_ | ~new_n11181_);
  assign new_n11199_ = new_n11193_ & ~new_n11200_ & new_n11189_;
  assign new_n11200_ = ~new_n11186_ & ~new_n11188_ & ~new_n11196_ & ~new_n11198_ & (~new_n11179_ | ~new_n11175_);
  assign new_n11201_ = new_n11189_ & new_n11185_ & new_n11193_ & ~new_n11196_ & ~new_n11198_;
  assign new_n11202_ = new_n11203_ & new_n11232_;
  assign new_n11203_ = ~new_n11204_ & ~new_n11228_;
  assign new_n11204_ = new_n11219_ & (~new_n11224_ | (~new_n11222_ & ~new_n11205_ & ~new_n11227_));
  assign new_n11205_ = ~new_n11217_ & ~new_n11215_ & (~new_n11218_ | ~new_n11214_ | new_n11206_);
  assign new_n11206_ = new_n11207_ & new_n11209_ & (new_n11212_ | ~\all_features[2813]  | ~\all_features[2814]  | ~\all_features[2815] );
  assign new_n11207_ = \all_features[2815]  & (\all_features[2814]  | (new_n11208_ & (\all_features[2810]  | \all_features[2811]  | \all_features[2809] )));
  assign new_n11208_ = \all_features[2812]  & \all_features[2813] ;
  assign new_n11209_ = \all_features[2814]  & \all_features[2815]  & (\all_features[2812]  | \all_features[2813]  | new_n11211_ | ~new_n11210_);
  assign new_n11210_ = ~\all_features[2810]  & ~\all_features[2811] ;
  assign new_n11211_ = \all_features[2808]  & \all_features[2809] ;
  assign new_n11212_ = ~\all_features[2811]  & ~\all_features[2812]  & (~\all_features[2810]  | new_n11213_);
  assign new_n11213_ = ~\all_features[2808]  & ~\all_features[2809] ;
  assign new_n11214_ = \all_features[2815]  & (\all_features[2814]  | (\all_features[2813]  & (\all_features[2812]  | ~new_n11210_ | ~new_n11213_)));
  assign new_n11215_ = ~new_n11216_ & ~\all_features[2815] ;
  assign new_n11216_ = \all_features[2813]  & \all_features[2814]  & (\all_features[2812]  | (\all_features[2810]  & \all_features[2811]  & \all_features[2809] ));
  assign new_n11217_ = ~\all_features[2815]  & (~new_n11211_ | ~\all_features[2810]  | ~\all_features[2811]  | ~\all_features[2814]  | ~new_n11208_);
  assign new_n11218_ = \all_features[2815]  & (\all_features[2813]  | \all_features[2814]  | \all_features[2812] );
  assign new_n11219_ = ~new_n11220_ & (\all_features[2811]  | \all_features[2812]  | \all_features[2813]  | \all_features[2814]  | \all_features[2815] );
  assign new_n11220_ = ~\all_features[2813]  & new_n11221_ & ((~\all_features[2810]  & new_n11213_) | ~\all_features[2812]  | ~\all_features[2811] );
  assign new_n11221_ = ~\all_features[2814]  & ~\all_features[2815] ;
  assign new_n11222_ = ~\all_features[2815]  & (~\all_features[2814]  | new_n11223_);
  assign new_n11223_ = ~\all_features[2813]  & (new_n11213_ | ~\all_features[2811]  | ~\all_features[2812]  | ~\all_features[2810] );
  assign new_n11224_ = ~new_n11225_ & ~new_n11226_;
  assign new_n11225_ = new_n11221_ & (~\all_features[2813]  | (~\all_features[2812]  & (~\all_features[2811]  | (~\all_features[2810]  & ~\all_features[2809] ))));
  assign new_n11226_ = new_n11221_ & (~\all_features[2811]  | ~new_n11208_ | (~new_n11211_ & ~\all_features[2810] ));
  assign new_n11227_ = ~\all_features[2815]  & (~\all_features[2814]  | (~\all_features[2813]  & ~\all_features[2812]  & (~\all_features[2811]  | ~\all_features[2810] )));
  assign new_n11228_ = ~new_n11229_ & (\all_features[2811]  | \all_features[2812]  | \all_features[2813]  | \all_features[2814]  | \all_features[2815] );
  assign new_n11229_ = ~new_n11220_ & (new_n11225_ | (~new_n11226_ & (new_n11227_ | (~new_n11222_ & ~new_n11230_))));
  assign new_n11230_ = ~new_n11215_ & (new_n11217_ | (new_n11218_ & (~new_n11214_ | (~new_n11231_ & new_n11207_))));
  assign new_n11231_ = ~\all_features[2813]  & \all_features[2814]  & \all_features[2815]  & (\all_features[2812]  ? new_n11210_ : (new_n11211_ | ~new_n11210_));
  assign new_n11232_ = ~new_n11233_ & ~new_n11236_;
  assign new_n11233_ = new_n11224_ & ~new_n11234_ & new_n11219_;
  assign new_n11234_ = ~new_n11227_ & ~new_n11217_ & ~new_n11215_ & ~new_n11222_ & ~new_n11235_;
  assign new_n11235_ = new_n11218_ & new_n11214_ & new_n11207_ & new_n11209_;
  assign new_n11236_ = new_n11219_ & new_n11237_ & ~new_n11215_ & ~new_n11225_;
  assign new_n11237_ = ~new_n11227_ & ~new_n11226_ & ~new_n11222_ & ~new_n11217_;
  assign new_n11238_ = ~new_n11267_ & (~new_n11260_ | ~new_n11239_ | ~new_n11269_);
  assign new_n11239_ = ~new_n11240_ & (\all_features[1011]  | \all_features[1012]  | \all_features[1013]  | \all_features[1014]  | \all_features[1015] );
  assign new_n11240_ = ~new_n11256_ & (new_n11254_ | (~new_n11258_ & (new_n11259_ | (~new_n11257_ & ~new_n11241_))));
  assign new_n11241_ = ~new_n11242_ & (new_n11244_ | (new_n11253_ & (~new_n11248_ | (~new_n11252_ & new_n11251_))));
  assign new_n11242_ = ~new_n11243_ & ~\all_features[1015] ;
  assign new_n11243_ = \all_features[1013]  & \all_features[1014]  & (\all_features[1012]  | (\all_features[1010]  & \all_features[1011]  & \all_features[1009] ));
  assign new_n11244_ = ~\all_features[1015]  & (~\all_features[1014]  | ~new_n11245_ | ~new_n11246_ | ~new_n11247_);
  assign new_n11245_ = \all_features[1010]  & \all_features[1011] ;
  assign new_n11246_ = \all_features[1008]  & \all_features[1009] ;
  assign new_n11247_ = \all_features[1012]  & \all_features[1013] ;
  assign new_n11248_ = \all_features[1015]  & (\all_features[1014]  | (\all_features[1013]  & (\all_features[1012]  | ~new_n11250_ | ~new_n11249_)));
  assign new_n11249_ = ~\all_features[1008]  & ~\all_features[1009] ;
  assign new_n11250_ = ~\all_features[1010]  & ~\all_features[1011] ;
  assign new_n11251_ = \all_features[1015]  & (\all_features[1014]  | (new_n11247_ & (\all_features[1010]  | \all_features[1011]  | \all_features[1009] )));
  assign new_n11252_ = ~\all_features[1013]  & \all_features[1014]  & \all_features[1015]  & (\all_features[1012]  ? new_n11250_ : (new_n11246_ | ~new_n11250_));
  assign new_n11253_ = \all_features[1015]  & (\all_features[1013]  | \all_features[1014]  | \all_features[1012] );
  assign new_n11254_ = new_n11255_ & (~\all_features[1013]  | (~\all_features[1012]  & (~\all_features[1011]  | (~\all_features[1010]  & ~\all_features[1009] ))));
  assign new_n11255_ = ~\all_features[1014]  & ~\all_features[1015] ;
  assign new_n11256_ = ~\all_features[1013]  & new_n11255_ & ((~\all_features[1010]  & new_n11249_) | ~\all_features[1012]  | ~\all_features[1011] );
  assign new_n11257_ = ~\all_features[1015]  & (~\all_features[1014]  | (~\all_features[1013]  & (new_n11249_ | ~new_n11245_ | ~\all_features[1012] )));
  assign new_n11258_ = new_n11255_ & (~\all_features[1011]  | ~new_n11247_ | (~\all_features[1010]  & ~new_n11246_));
  assign new_n11259_ = ~\all_features[1015]  & (~\all_features[1014]  | (~\all_features[1012]  & ~\all_features[1013]  & ~new_n11245_));
  assign new_n11260_ = new_n11265_ & (~new_n11266_ | (~new_n11261_ & ~new_n11257_ & ~new_n11259_));
  assign new_n11261_ = ~new_n11242_ & ~new_n11244_ & (~new_n11253_ | ~new_n11248_ | new_n11262_);
  assign new_n11262_ = new_n11251_ & new_n11263_ & (new_n11264_ | ~\all_features[1013]  | ~\all_features[1014]  | ~\all_features[1015] );
  assign new_n11263_ = \all_features[1014]  & \all_features[1015]  & (\all_features[1012]  | \all_features[1013]  | new_n11246_ | ~new_n11250_);
  assign new_n11264_ = ~\all_features[1011]  & ~\all_features[1012]  & (~\all_features[1010]  | new_n11249_);
  assign new_n11265_ = ~new_n11256_ & (\all_features[1011]  | \all_features[1012]  | \all_features[1013]  | \all_features[1014]  | \all_features[1015] );
  assign new_n11266_ = ~new_n11254_ & ~new_n11258_;
  assign new_n11267_ = new_n11268_ & new_n11265_ & ~new_n11258_ & ~new_n11257_ & ~new_n11242_ & ~new_n11254_;
  assign new_n11268_ = ~new_n11244_ & ~new_n11259_;
  assign new_n11269_ = new_n11265_ & new_n11266_ & (new_n11270_ | new_n11242_ | new_n11257_ | ~new_n11268_);
  assign new_n11270_ = new_n11253_ & new_n11263_ & new_n11248_ & new_n11251_;
  assign new_n11271_ = (new_n11272_ | ~new_n11166_ | ~new_n11170_) & (~new_n11202_ | ~new_n11273_ | new_n11170_);
  assign new_n11272_ = new_n11026_ & ~new_n11055_ & ~new_n11059_;
  assign new_n11273_ = new_n11301_ & (new_n11297_ | new_n11274_);
  assign new_n11274_ = new_n11294_ & ~new_n11275_ & new_n11289_;
  assign new_n11275_ = ~new_n11283_ & ~new_n11285_ & ~new_n11286_ & ~new_n11288_ & (~new_n11279_ | ~new_n11276_);
  assign new_n11276_ = \all_features[3911]  & (\all_features[3910]  | (~new_n11277_ & \all_features[3909] ));
  assign new_n11277_ = new_n11278_ & ~\all_features[3908]  & ~\all_features[3906]  & ~\all_features[3907] ;
  assign new_n11278_ = ~\all_features[3904]  & ~\all_features[3905] ;
  assign new_n11279_ = \all_features[3911]  & \all_features[3910]  & ~new_n11282_ & new_n11280_;
  assign new_n11280_ = \all_features[3911]  & (\all_features[3910]  | (new_n11281_ & (\all_features[3906]  | \all_features[3907]  | \all_features[3905] )));
  assign new_n11281_ = \all_features[3908]  & \all_features[3909] ;
  assign new_n11282_ = ~\all_features[3906]  & ~\all_features[3907]  & ~\all_features[3908]  & ~\all_features[3909]  & (~\all_features[3905]  | ~\all_features[3904] );
  assign new_n11283_ = ~\all_features[3911]  & (~\all_features[3910]  | (~\all_features[3908]  & ~\all_features[3909]  & ~new_n11284_));
  assign new_n11284_ = \all_features[3906]  & \all_features[3907] ;
  assign new_n11285_ = ~\all_features[3911]  & (~\all_features[3910]  | (~\all_features[3909]  & (new_n11278_ | ~\all_features[3908]  | ~new_n11284_)));
  assign new_n11286_ = ~new_n11287_ & ~\all_features[3911] ;
  assign new_n11287_ = \all_features[3909]  & \all_features[3910]  & (\all_features[3908]  | (\all_features[3906]  & \all_features[3907]  & \all_features[3905] ));
  assign new_n11288_ = ~\all_features[3911]  & (~new_n11281_ | ~\all_features[3904]  | ~\all_features[3905]  | ~\all_features[3910]  | ~new_n11284_);
  assign new_n11289_ = ~new_n11290_ & ~new_n11293_;
  assign new_n11290_ = new_n11291_ & ((~\all_features[3906]  & new_n11278_) | ~\all_features[3908]  | ~\all_features[3907] );
  assign new_n11291_ = ~\all_features[3909]  & new_n11292_;
  assign new_n11292_ = ~\all_features[3910]  & ~\all_features[3911] ;
  assign new_n11293_ = new_n11291_ & ~\all_features[3907]  & ~\all_features[3908] ;
  assign new_n11294_ = ~new_n11295_ & ~new_n11296_;
  assign new_n11295_ = new_n11292_ & (~new_n11281_ | ~\all_features[3907]  | (~\all_features[3906]  & (~\all_features[3904]  | ~\all_features[3905] )));
  assign new_n11296_ = new_n11292_ & (~\all_features[3909]  | (~\all_features[3908]  & (~\all_features[3907]  | (~\all_features[3906]  & ~\all_features[3905] ))));
  assign new_n11297_ = new_n11289_ & (~new_n11294_ | (new_n11300_ & (new_n11298_ | new_n11286_ | new_n11288_)));
  assign new_n11298_ = new_n11276_ & (~new_n11279_ | (~new_n11299_ & \all_features[3909]  & \all_features[3910]  & \all_features[3911] ));
  assign new_n11299_ = ~\all_features[3907]  & ~\all_features[3908]  & (~\all_features[3906]  | new_n11278_);
  assign new_n11300_ = ~new_n11283_ & ~new_n11285_;
  assign new_n11301_ = new_n11294_ & new_n11300_ & ~new_n11288_ & ~new_n11286_ & ~new_n11290_ & ~new_n11293_;
  assign new_n11302_ = new_n11303_ ? new_n11373_ : ~new_n11337_;
  assign new_n11303_ = new_n11335_ & ~new_n11304_ & new_n11333_;
  assign new_n11304_ = ~new_n11305_ & ~new_n11329_;
  assign new_n11305_ = new_n11321_ & (~new_n11324_ | (~new_n11306_ & ~new_n11327_ & ~new_n11328_));
  assign new_n11306_ = ~new_n11318_ & ~new_n11316_ & (~new_n11320_ | ~new_n11315_ | new_n11307_);
  assign new_n11307_ = new_n11308_ & new_n11310_ & (new_n11313_ | ~\all_features[3069]  | ~\all_features[3070]  | ~\all_features[3071] );
  assign new_n11308_ = \all_features[3071]  & (\all_features[3070]  | (new_n11309_ & (\all_features[3066]  | \all_features[3067]  | \all_features[3065] )));
  assign new_n11309_ = \all_features[3068]  & \all_features[3069] ;
  assign new_n11310_ = \all_features[3070]  & \all_features[3071]  & (\all_features[3068]  | \all_features[3069]  | new_n11312_ | ~new_n11311_);
  assign new_n11311_ = ~\all_features[3066]  & ~\all_features[3067] ;
  assign new_n11312_ = \all_features[3064]  & \all_features[3065] ;
  assign new_n11313_ = ~\all_features[3067]  & ~\all_features[3068]  & (~\all_features[3066]  | new_n11314_);
  assign new_n11314_ = ~\all_features[3064]  & ~\all_features[3065] ;
  assign new_n11315_ = \all_features[3071]  & (\all_features[3070]  | (\all_features[3069]  & (\all_features[3068]  | ~new_n11311_ | ~new_n11314_)));
  assign new_n11316_ = ~\all_features[3071]  & (~\all_features[3070]  | ~new_n11309_ | ~new_n11312_ | ~new_n11317_);
  assign new_n11317_ = \all_features[3066]  & \all_features[3067] ;
  assign new_n11318_ = ~new_n11319_ & ~\all_features[3071] ;
  assign new_n11319_ = \all_features[3069]  & \all_features[3070]  & (\all_features[3068]  | (\all_features[3066]  & \all_features[3067]  & \all_features[3065] ));
  assign new_n11320_ = \all_features[3071]  & (\all_features[3069]  | \all_features[3070]  | \all_features[3068] );
  assign new_n11321_ = ~new_n11322_ & (\all_features[3067]  | \all_features[3068]  | \all_features[3069]  | \all_features[3070]  | \all_features[3071] );
  assign new_n11322_ = ~\all_features[3069]  & new_n11323_ & ((~\all_features[3066]  & new_n11314_) | ~\all_features[3068]  | ~\all_features[3067] );
  assign new_n11323_ = ~\all_features[3070]  & ~\all_features[3071] ;
  assign new_n11324_ = ~new_n11325_ & ~new_n11326_;
  assign new_n11325_ = new_n11323_ & (~\all_features[3069]  | (~\all_features[3068]  & (~\all_features[3067]  | (~\all_features[3066]  & ~\all_features[3065] ))));
  assign new_n11326_ = new_n11323_ & (~\all_features[3067]  | ~new_n11309_ | (~new_n11312_ & ~\all_features[3066] ));
  assign new_n11327_ = ~\all_features[3071]  & (~\all_features[3070]  | (~\all_features[3069]  & (new_n11314_ | ~new_n11317_ | ~\all_features[3068] )));
  assign new_n11328_ = ~\all_features[3071]  & (~\all_features[3070]  | (~\all_features[3068]  & ~\all_features[3069]  & ~new_n11317_));
  assign new_n11329_ = ~new_n11330_ & (\all_features[3067]  | \all_features[3068]  | \all_features[3069]  | \all_features[3070]  | \all_features[3071] );
  assign new_n11330_ = ~new_n11322_ & (new_n11325_ | (~new_n11326_ & (new_n11328_ | (~new_n11327_ & ~new_n11331_))));
  assign new_n11331_ = ~new_n11318_ & (new_n11316_ | (new_n11320_ & (~new_n11315_ | (~new_n11332_ & new_n11308_))));
  assign new_n11332_ = ~\all_features[3069]  & \all_features[3070]  & \all_features[3071]  & (\all_features[3068]  ? new_n11311_ : (new_n11312_ | ~new_n11311_));
  assign new_n11333_ = new_n11334_ & new_n11321_ & ~new_n11326_ & ~new_n11325_ & ~new_n11318_ & ~new_n11327_;
  assign new_n11334_ = ~new_n11316_ & ~new_n11328_;
  assign new_n11335_ = new_n11321_ & new_n11324_ & (new_n11336_ | new_n11318_ | new_n11327_ | ~new_n11334_);
  assign new_n11336_ = new_n11320_ & new_n11315_ & new_n11308_ & new_n11310_;
  assign new_n11337_ = new_n11338_ & new_n11364_;
  assign new_n11338_ = ~new_n11339_ & ~new_n11361_;
  assign new_n11339_ = ~new_n11360_ & ~new_n11359_ & ~new_n11358_ & ~new_n11340_ & ~new_n11356_;
  assign new_n11340_ = new_n11341_ & (~new_n11354_ | ~new_n11355_ | ~new_n11351_ | ~new_n11353_);
  assign new_n11341_ = ~new_n11348_ & ~new_n11347_ & ~new_n11342_ & ~new_n11345_;
  assign new_n11342_ = ~\all_features[2407]  & (~\all_features[2406]  | (~\all_features[2405]  & (new_n11343_ | ~new_n11344_ | ~\all_features[2404] )));
  assign new_n11343_ = ~\all_features[2400]  & ~\all_features[2401] ;
  assign new_n11344_ = \all_features[2402]  & \all_features[2403] ;
  assign new_n11345_ = ~new_n11346_ & ~\all_features[2407] ;
  assign new_n11346_ = \all_features[2405]  & \all_features[2406]  & (\all_features[2404]  | (\all_features[2402]  & \all_features[2403]  & \all_features[2401] ));
  assign new_n11347_ = ~\all_features[2407]  & (~\all_features[2406]  | (~\all_features[2404]  & ~\all_features[2405]  & ~new_n11344_));
  assign new_n11348_ = ~\all_features[2407]  & (~\all_features[2406]  | ~new_n11349_ | ~new_n11350_ | ~new_n11344_);
  assign new_n11349_ = \all_features[2404]  & \all_features[2405] ;
  assign new_n11350_ = \all_features[2400]  & \all_features[2401] ;
  assign new_n11351_ = \all_features[2407]  & (\all_features[2406]  | (\all_features[2405]  & (\all_features[2404]  | ~new_n11343_ | ~new_n11352_)));
  assign new_n11352_ = ~\all_features[2402]  & ~\all_features[2403] ;
  assign new_n11353_ = \all_features[2407]  & (\all_features[2406]  | (new_n11349_ & (\all_features[2402]  | \all_features[2403]  | \all_features[2401] )));
  assign new_n11354_ = \all_features[2406]  & \all_features[2407]  & (\all_features[2404]  | \all_features[2405]  | new_n11350_ | ~new_n11352_);
  assign new_n11355_ = \all_features[2407]  & (\all_features[2405]  | \all_features[2406]  | \all_features[2404] );
  assign new_n11356_ = new_n11357_ & (~\all_features[2405]  | (~\all_features[2404]  & (~\all_features[2403]  | (~\all_features[2402]  & ~\all_features[2401] ))));
  assign new_n11357_ = ~\all_features[2406]  & ~\all_features[2407] ;
  assign new_n11358_ = ~\all_features[2405]  & new_n11357_ & ((~\all_features[2402]  & new_n11343_) | ~\all_features[2404]  | ~\all_features[2403] );
  assign new_n11359_ = new_n11357_ & (~\all_features[2403]  | ~new_n11349_ | (~\all_features[2402]  & ~new_n11350_));
  assign new_n11360_ = ~\all_features[2407]  & ~\all_features[2406]  & ~\all_features[2405]  & ~\all_features[2403]  & ~\all_features[2404] ;
  assign new_n11361_ = new_n11363_ & new_n11362_ & ~new_n11358_ & ~new_n11348_ & ~new_n11342_ & ~new_n11345_;
  assign new_n11362_ = ~new_n11347_ & ~new_n11360_;
  assign new_n11363_ = ~new_n11356_ & ~new_n11359_;
  assign new_n11364_ = ~new_n11365_ & ~new_n11369_;
  assign new_n11365_ = ~new_n11358_ & ~new_n11360_ & (~new_n11363_ | (~new_n11366_ & ~new_n11342_ & ~new_n11347_));
  assign new_n11366_ = ~new_n11348_ & ~new_n11345_ & (~new_n11355_ | ~new_n11351_ | new_n11367_);
  assign new_n11367_ = new_n11353_ & new_n11354_ & (new_n11368_ | ~\all_features[2405]  | ~\all_features[2406]  | ~\all_features[2407] );
  assign new_n11368_ = ~\all_features[2403]  & ~\all_features[2404]  & (~\all_features[2402]  | new_n11343_);
  assign new_n11369_ = ~new_n11370_ & ~new_n11360_;
  assign new_n11370_ = ~new_n11358_ & (new_n11356_ | (~new_n11359_ & (new_n11347_ | (~new_n11342_ & ~new_n11371_))));
  assign new_n11371_ = ~new_n11345_ & (new_n11348_ | (new_n11355_ & (~new_n11351_ | (~new_n11372_ & new_n11353_))));
  assign new_n11372_ = ~\all_features[2405]  & \all_features[2406]  & \all_features[2407]  & (\all_features[2404]  ? new_n11352_ : (new_n11350_ | ~new_n11352_));
  assign new_n11373_ = ~new_n7041_ & ~new_n7063_;
  assign new_n11374_ = (new_n11550_ | ~new_n11549_ | new_n11515_) & (~new_n11515_ | (~new_n11375_ & (new_n11471_ | new_n11376_)));
  assign new_n11375_ = (new_n11471_ & (new_n11377_ ? new_n11498_ : ~new_n11411_)) | (new_n11445_ & new_n11376_ & ~new_n11471_);
  assign new_n11376_ = new_n8594_ & (new_n8591_ | new_n8558_);
  assign new_n11377_ = ~new_n11407_ & (~new_n11409_ | ~new_n11378_);
  assign new_n11378_ = new_n11379_ & new_n11403_;
  assign new_n11379_ = new_n11395_ & (~new_n11398_ | (~new_n11380_ & ~new_n11401_ & ~new_n11402_));
  assign new_n11380_ = ~new_n11389_ & ~new_n11391_ & (~new_n11394_ | ~new_n11393_ | new_n11381_);
  assign new_n11381_ = new_n11382_ & new_n11384_ & (new_n11387_ | ~\all_features[2085]  | ~\all_features[2086]  | ~\all_features[2087] );
  assign new_n11382_ = \all_features[2087]  & (\all_features[2086]  | (new_n11383_ & (\all_features[2082]  | \all_features[2083]  | \all_features[2081] )));
  assign new_n11383_ = \all_features[2084]  & \all_features[2085] ;
  assign new_n11384_ = \all_features[2086]  & \all_features[2087]  & (\all_features[2084]  | \all_features[2085]  | new_n11385_ | ~new_n11386_);
  assign new_n11385_ = \all_features[2080]  & \all_features[2081] ;
  assign new_n11386_ = ~\all_features[2082]  & ~\all_features[2083] ;
  assign new_n11387_ = ~\all_features[2083]  & ~\all_features[2084]  & (~\all_features[2082]  | new_n11388_);
  assign new_n11388_ = ~\all_features[2080]  & ~\all_features[2081] ;
  assign new_n11389_ = ~new_n11390_ & ~\all_features[2087] ;
  assign new_n11390_ = \all_features[2085]  & \all_features[2086]  & (\all_features[2084]  | (\all_features[2082]  & \all_features[2083]  & \all_features[2081] ));
  assign new_n11391_ = ~\all_features[2087]  & (~\all_features[2086]  | ~new_n11392_ | ~new_n11385_ | ~new_n11383_);
  assign new_n11392_ = \all_features[2082]  & \all_features[2083] ;
  assign new_n11393_ = \all_features[2087]  & (\all_features[2086]  | (\all_features[2085]  & (\all_features[2084]  | ~new_n11386_ | ~new_n11388_)));
  assign new_n11394_ = \all_features[2087]  & (\all_features[2085]  | \all_features[2086]  | \all_features[2084] );
  assign new_n11395_ = ~new_n11396_ & (\all_features[2083]  | \all_features[2084]  | \all_features[2085]  | \all_features[2086]  | \all_features[2087] );
  assign new_n11396_ = ~\all_features[2085]  & new_n11397_ & ((~\all_features[2082]  & new_n11388_) | ~\all_features[2084]  | ~\all_features[2083] );
  assign new_n11397_ = ~\all_features[2086]  & ~\all_features[2087] ;
  assign new_n11398_ = ~new_n11399_ & ~new_n11400_;
  assign new_n11399_ = new_n11397_ & (~\all_features[2085]  | (~\all_features[2084]  & (~\all_features[2083]  | (~\all_features[2082]  & ~\all_features[2081] ))));
  assign new_n11400_ = new_n11397_ & (~\all_features[2083]  | ~new_n11383_ | (~\all_features[2082]  & ~new_n11385_));
  assign new_n11401_ = ~\all_features[2087]  & (~\all_features[2086]  | (~\all_features[2085]  & (new_n11388_ | ~new_n11392_ | ~\all_features[2084] )));
  assign new_n11402_ = ~\all_features[2087]  & (~\all_features[2086]  | (~\all_features[2084]  & ~\all_features[2085]  & ~new_n11392_));
  assign new_n11403_ = ~new_n11404_ & (\all_features[2083]  | \all_features[2084]  | \all_features[2085]  | \all_features[2086]  | \all_features[2087] );
  assign new_n11404_ = ~new_n11396_ & (new_n11399_ | (~new_n11400_ & (new_n11402_ | (~new_n11401_ & ~new_n11405_))));
  assign new_n11405_ = ~new_n11389_ & (new_n11391_ | (new_n11394_ & (~new_n11393_ | (~new_n11406_ & new_n11382_))));
  assign new_n11406_ = ~\all_features[2085]  & \all_features[2086]  & \all_features[2087]  & (\all_features[2084]  ? new_n11386_ : (new_n11385_ | ~new_n11386_));
  assign new_n11407_ = new_n11408_ & new_n11395_ & ~new_n11400_ & ~new_n11401_ & ~new_n11389_ & ~new_n11399_;
  assign new_n11408_ = ~new_n11391_ & ~new_n11402_;
  assign new_n11409_ = new_n11395_ & new_n11398_ & (new_n11410_ | new_n11389_ | new_n11401_ | ~new_n11408_);
  assign new_n11410_ = new_n11394_ & new_n11384_ & new_n11393_ & new_n11382_;
  assign new_n11411_ = new_n11444_ & (new_n11442_ | new_n11412_);
  assign new_n11412_ = new_n11413_ & new_n11433_;
  assign new_n11413_ = ~new_n11432_ & (new_n11431_ | (~new_n11430_ & (new_n11428_ | (~new_n11427_ & ~new_n11414_))));
  assign new_n11414_ = ~new_n11421_ & (new_n11423_ | (~new_n11425_ & (~new_n11426_ | new_n11415_)));
  assign new_n11415_ = \all_features[4855]  & ((~new_n11420_ & ~\all_features[4853]  & \all_features[4854] ) | (~new_n11418_ & (\all_features[4854]  | (~new_n11416_ & \all_features[4853] ))));
  assign new_n11416_ = new_n11417_ & ~\all_features[4852]  & ~\all_features[4850]  & ~\all_features[4851] ;
  assign new_n11417_ = ~\all_features[4848]  & ~\all_features[4849] ;
  assign new_n11418_ = \all_features[4855]  & (\all_features[4854]  | (new_n11419_ & (\all_features[4850]  | \all_features[4851]  | \all_features[4849] )));
  assign new_n11419_ = \all_features[4852]  & \all_features[4853] ;
  assign new_n11420_ = (~\all_features[4850]  & ~\all_features[4851]  & ~\all_features[4852]  & (~\all_features[4849]  | ~\all_features[4848] )) | (\all_features[4852]  & (\all_features[4850]  | \all_features[4851] ));
  assign new_n11421_ = ~\all_features[4855]  & (~\all_features[4854]  | (~\all_features[4853]  & (new_n11417_ | ~\all_features[4852]  | ~new_n11422_)));
  assign new_n11422_ = \all_features[4850]  & \all_features[4851] ;
  assign new_n11423_ = ~new_n11424_ & ~\all_features[4855] ;
  assign new_n11424_ = \all_features[4853]  & \all_features[4854]  & (\all_features[4852]  | (\all_features[4850]  & \all_features[4851]  & \all_features[4849] ));
  assign new_n11425_ = ~\all_features[4855]  & (~new_n11419_ | ~\all_features[4848]  | ~\all_features[4849]  | ~\all_features[4854]  | ~new_n11422_);
  assign new_n11426_ = \all_features[4855]  & (\all_features[4853]  | \all_features[4854]  | \all_features[4852] );
  assign new_n11427_ = ~\all_features[4855]  & (~\all_features[4854]  | (~\all_features[4852]  & ~\all_features[4853]  & ~new_n11422_));
  assign new_n11428_ = new_n11429_ & (~new_n11419_ | ~\all_features[4851]  | (~\all_features[4850]  & (~\all_features[4848]  | ~\all_features[4849] )));
  assign new_n11429_ = ~\all_features[4854]  & ~\all_features[4855] ;
  assign new_n11430_ = new_n11429_ & (~\all_features[4853]  | (~\all_features[4852]  & (~\all_features[4851]  | (~\all_features[4850]  & ~\all_features[4849] ))));
  assign new_n11431_ = ~\all_features[4853]  & new_n11429_ & ((~\all_features[4850]  & new_n11417_) | ~\all_features[4852]  | ~\all_features[4851] );
  assign new_n11432_ = ~\all_features[4855]  & ~\all_features[4854]  & ~\all_features[4853]  & ~\all_features[4851]  & ~\all_features[4852] ;
  assign new_n11433_ = new_n11441_ & (~new_n11440_ | (new_n11439_ & (new_n11434_ | new_n11423_ | new_n11425_)));
  assign new_n11434_ = new_n11435_ & (~new_n11436_ | (~new_n11438_ & \all_features[4853]  & \all_features[4854]  & \all_features[4855] ));
  assign new_n11435_ = \all_features[4855]  & (\all_features[4854]  | (~new_n11416_ & \all_features[4853] ));
  assign new_n11436_ = \all_features[4855]  & \all_features[4854]  & ~new_n11437_ & new_n11418_;
  assign new_n11437_ = ~\all_features[4850]  & ~\all_features[4851]  & ~\all_features[4852]  & ~\all_features[4853]  & (~\all_features[4849]  | ~\all_features[4848] );
  assign new_n11438_ = ~\all_features[4851]  & ~\all_features[4852]  & (~\all_features[4850]  | new_n11417_);
  assign new_n11439_ = ~new_n11421_ & ~new_n11427_;
  assign new_n11440_ = ~new_n11428_ & ~new_n11430_;
  assign new_n11441_ = ~new_n11431_ & ~new_n11432_;
  assign new_n11442_ = new_n11441_ & ~new_n11443_ & new_n11440_;
  assign new_n11443_ = ~new_n11421_ & ~new_n11427_ & ~new_n11423_ & ~new_n11425_ & (~new_n11436_ | ~new_n11435_);
  assign new_n11444_ = new_n11440_ & new_n11439_ & new_n11441_ & ~new_n11423_ & ~new_n11425_;
  assign new_n11445_ = ~new_n11446_ & ~new_n11468_;
  assign new_n11446_ = ~new_n11467_ & ~new_n11466_ & ~new_n11465_ & ~new_n11447_ & ~new_n11463_;
  assign new_n11447_ = new_n11448_ & (~new_n11461_ | ~new_n11462_ | ~new_n11458_ | ~new_n11460_);
  assign new_n11448_ = ~new_n11455_ & ~new_n11454_ & ~new_n11449_ & ~new_n11452_;
  assign new_n11449_ = ~\all_features[5039]  & (~\all_features[5038]  | (~\all_features[5037]  & (new_n11450_ | ~new_n11451_ | ~\all_features[5036] )));
  assign new_n11450_ = ~\all_features[5032]  & ~\all_features[5033] ;
  assign new_n11451_ = \all_features[5034]  & \all_features[5035] ;
  assign new_n11452_ = ~new_n11453_ & ~\all_features[5039] ;
  assign new_n11453_ = \all_features[5037]  & \all_features[5038]  & (\all_features[5036]  | (\all_features[5034]  & \all_features[5035]  & \all_features[5033] ));
  assign new_n11454_ = ~\all_features[5039]  & (~\all_features[5038]  | (~\all_features[5036]  & ~\all_features[5037]  & ~new_n11451_));
  assign new_n11455_ = ~\all_features[5039]  & (~\all_features[5038]  | ~new_n11456_ | ~new_n11457_ | ~new_n11451_);
  assign new_n11456_ = \all_features[5036]  & \all_features[5037] ;
  assign new_n11457_ = \all_features[5032]  & \all_features[5033] ;
  assign new_n11458_ = \all_features[5039]  & (\all_features[5038]  | (\all_features[5037]  & (\all_features[5036]  | ~new_n11450_ | ~new_n11459_)));
  assign new_n11459_ = ~\all_features[5034]  & ~\all_features[5035] ;
  assign new_n11460_ = \all_features[5039]  & (\all_features[5038]  | (new_n11456_ & (\all_features[5034]  | \all_features[5035]  | \all_features[5033] )));
  assign new_n11461_ = \all_features[5038]  & \all_features[5039]  & (\all_features[5036]  | \all_features[5037]  | new_n11457_ | ~new_n11459_);
  assign new_n11462_ = \all_features[5039]  & (\all_features[5037]  | \all_features[5038]  | \all_features[5036] );
  assign new_n11463_ = new_n11464_ & (~\all_features[5037]  | (~\all_features[5036]  & (~\all_features[5035]  | (~\all_features[5034]  & ~\all_features[5033] ))));
  assign new_n11464_ = ~\all_features[5038]  & ~\all_features[5039] ;
  assign new_n11465_ = ~\all_features[5037]  & new_n11464_ & ((~\all_features[5034]  & new_n11450_) | ~\all_features[5036]  | ~\all_features[5035] );
  assign new_n11466_ = new_n11464_ & (~\all_features[5035]  | ~new_n11456_ | (~\all_features[5034]  & ~new_n11457_));
  assign new_n11467_ = ~\all_features[5039]  & ~\all_features[5038]  & ~\all_features[5037]  & ~\all_features[5035]  & ~\all_features[5036] ;
  assign new_n11468_ = new_n11470_ & new_n11469_ & ~new_n11465_ & ~new_n11455_ & ~new_n11449_ & ~new_n11452_;
  assign new_n11469_ = ~new_n11454_ & ~new_n11467_;
  assign new_n11470_ = ~new_n11463_ & ~new_n11466_;
  assign new_n11471_ = new_n11497_ | ((new_n11493_ | (~new_n11472_ & ~new_n11494_ & ~new_n11496_)) & (new_n11493_ | new_n11494_ | new_n11496_));
  assign new_n11472_ = new_n11486_ & (~new_n11481_ | (~new_n11473_ & new_n11489_ & new_n11490_));
  assign new_n11473_ = new_n11474_ & new_n11478_ & (new_n11476_ | ~\all_features[5085]  | ~\all_features[5086]  | ~\all_features[5087] );
  assign new_n11474_ = \all_features[5087]  & (\all_features[5086]  | (new_n11475_ & (\all_features[5082]  | \all_features[5083]  | \all_features[5081] )));
  assign new_n11475_ = \all_features[5084]  & \all_features[5085] ;
  assign new_n11476_ = ~\all_features[5083]  & ~\all_features[5084]  & (~\all_features[5082]  | new_n11477_);
  assign new_n11477_ = ~\all_features[5080]  & ~\all_features[5081] ;
  assign new_n11478_ = \all_features[5086]  & \all_features[5087]  & (\all_features[5084]  | \all_features[5085]  | new_n11480_ | ~new_n11479_);
  assign new_n11479_ = ~\all_features[5082]  & ~\all_features[5083] ;
  assign new_n11480_ = \all_features[5080]  & \all_features[5081] ;
  assign new_n11481_ = ~new_n11482_ & ~new_n11484_;
  assign new_n11482_ = ~new_n11483_ & ~\all_features[5087] ;
  assign new_n11483_ = \all_features[5085]  & \all_features[5086]  & (\all_features[5084]  | (\all_features[5082]  & \all_features[5083]  & \all_features[5081] ));
  assign new_n11484_ = ~\all_features[5087]  & (~\all_features[5086]  | ~new_n11475_ | ~new_n11480_ | ~new_n11485_);
  assign new_n11485_ = \all_features[5082]  & \all_features[5083] ;
  assign new_n11486_ = ~new_n11487_ & ~new_n11488_;
  assign new_n11487_ = ~\all_features[5087]  & (~\all_features[5086]  | (~\all_features[5084]  & ~\all_features[5085]  & ~new_n11485_));
  assign new_n11488_ = ~\all_features[5087]  & (~\all_features[5086]  | (~\all_features[5085]  & (new_n11477_ | ~new_n11485_ | ~\all_features[5084] )));
  assign new_n11489_ = \all_features[5087]  & (\all_features[5086]  | (\all_features[5085]  & (\all_features[5084]  | ~new_n11479_ | ~new_n11477_)));
  assign new_n11490_ = \all_features[5087]  & (\all_features[5085]  | \all_features[5086]  | \all_features[5084] );
  assign new_n11493_ = ~\all_features[5087]  & ~\all_features[5086]  & ~\all_features[5085]  & ~\all_features[5083]  & ~\all_features[5084] ;
  assign new_n11494_ = new_n11495_ & (~\all_features[5085]  | (~\all_features[5084]  & (~\all_features[5083]  | (~\all_features[5082]  & ~\all_features[5081] ))));
  assign new_n11495_ = ~\all_features[5086]  & ~\all_features[5087] ;
  assign new_n11496_ = new_n11495_ & (~\all_features[5083]  | ~new_n11475_ | (~\all_features[5082]  & ~new_n11480_));
  assign new_n11497_ = ~\all_features[5085]  & new_n11495_ & ((~\all_features[5082]  & new_n11477_) | ~\all_features[5084]  | ~\all_features[5083] );
  assign new_n11498_ = new_n11505_ & new_n11499_ & ~new_n11514_ & ~new_n11512_ & ~new_n11509_ & ~new_n11511_;
  assign new_n11499_ = ~new_n11500_ & ~new_n11504_;
  assign new_n11500_ = ~\all_features[799]  & (~\all_features[798]  | ~new_n11501_ | ~new_n11502_ | ~new_n11503_);
  assign new_n11501_ = \all_features[792]  & \all_features[793] ;
  assign new_n11502_ = \all_features[796]  & \all_features[797] ;
  assign new_n11503_ = \all_features[794]  & \all_features[795] ;
  assign new_n11504_ = ~\all_features[799]  & ~\all_features[798]  & ~\all_features[797]  & ~\all_features[795]  & ~\all_features[796] ;
  assign new_n11505_ = ~new_n11506_ & ~new_n11508_;
  assign new_n11506_ = new_n11507_ & (~\all_features[795]  | ~new_n11502_ | (~\all_features[794]  & ~new_n11501_));
  assign new_n11507_ = ~\all_features[798]  & ~\all_features[799] ;
  assign new_n11508_ = new_n11507_ & (~\all_features[797]  | (~\all_features[796]  & (~\all_features[795]  | (~\all_features[794]  & ~\all_features[793] ))));
  assign new_n11509_ = ~new_n11510_ & ~\all_features[799] ;
  assign new_n11510_ = \all_features[797]  & \all_features[798]  & (\all_features[796]  | (\all_features[794]  & \all_features[795]  & \all_features[793] ));
  assign new_n11511_ = ~\all_features[799]  & (~\all_features[798]  | (~\all_features[796]  & ~\all_features[797]  & ~new_n11503_));
  assign new_n11512_ = ~\all_features[797]  & new_n11507_ & ((~\all_features[794]  & new_n11513_) | ~\all_features[796]  | ~\all_features[795] );
  assign new_n11513_ = ~\all_features[792]  & ~\all_features[793] ;
  assign new_n11514_ = ~\all_features[799]  & (~\all_features[798]  | (~\all_features[797]  & (new_n11513_ | ~\all_features[796]  | ~new_n11503_)));
  assign new_n11515_ = ~new_n11545_ & (~new_n11547_ | ~new_n11516_);
  assign new_n11516_ = new_n11517_ & new_n11541_;
  assign new_n11517_ = new_n11533_ & (~new_n11536_ | (~new_n11518_ & ~new_n11539_ & ~new_n11540_));
  assign new_n11518_ = ~new_n11527_ & ~new_n11529_ & (~new_n11532_ | ~new_n11531_ | new_n11519_);
  assign new_n11519_ = new_n11520_ & new_n11522_ & (new_n11525_ | ~\all_features[3557]  | ~\all_features[3558]  | ~\all_features[3559] );
  assign new_n11520_ = \all_features[3559]  & (\all_features[3558]  | (new_n11521_ & (\all_features[3554]  | \all_features[3555]  | \all_features[3553] )));
  assign new_n11521_ = \all_features[3556]  & \all_features[3557] ;
  assign new_n11522_ = \all_features[3558]  & \all_features[3559]  & (\all_features[3556]  | \all_features[3557]  | new_n11523_ | ~new_n11524_);
  assign new_n11523_ = \all_features[3552]  & \all_features[3553] ;
  assign new_n11524_ = ~\all_features[3554]  & ~\all_features[3555] ;
  assign new_n11525_ = ~\all_features[3555]  & ~\all_features[3556]  & (~\all_features[3554]  | new_n11526_);
  assign new_n11526_ = ~\all_features[3552]  & ~\all_features[3553] ;
  assign new_n11527_ = ~new_n11528_ & ~\all_features[3559] ;
  assign new_n11528_ = \all_features[3557]  & \all_features[3558]  & (\all_features[3556]  | (\all_features[3554]  & \all_features[3555]  & \all_features[3553] ));
  assign new_n11529_ = ~\all_features[3559]  & (~\all_features[3558]  | ~new_n11530_ | ~new_n11523_ | ~new_n11521_);
  assign new_n11530_ = \all_features[3554]  & \all_features[3555] ;
  assign new_n11531_ = \all_features[3559]  & (\all_features[3558]  | (\all_features[3557]  & (\all_features[3556]  | ~new_n11524_ | ~new_n11526_)));
  assign new_n11532_ = \all_features[3559]  & (\all_features[3557]  | \all_features[3558]  | \all_features[3556] );
  assign new_n11533_ = ~new_n11534_ & (\all_features[3555]  | \all_features[3556]  | \all_features[3557]  | \all_features[3558]  | \all_features[3559] );
  assign new_n11534_ = ~\all_features[3557]  & new_n11535_ & ((~\all_features[3554]  & new_n11526_) | ~\all_features[3556]  | ~\all_features[3555] );
  assign new_n11535_ = ~\all_features[3558]  & ~\all_features[3559] ;
  assign new_n11536_ = ~new_n11537_ & ~new_n11538_;
  assign new_n11537_ = new_n11535_ & (~\all_features[3557]  | (~\all_features[3556]  & (~\all_features[3555]  | (~\all_features[3554]  & ~\all_features[3553] ))));
  assign new_n11538_ = new_n11535_ & (~\all_features[3555]  | ~new_n11521_ | (~\all_features[3554]  & ~new_n11523_));
  assign new_n11539_ = ~\all_features[3559]  & (~\all_features[3558]  | (~\all_features[3557]  & (new_n11526_ | ~new_n11530_ | ~\all_features[3556] )));
  assign new_n11540_ = ~\all_features[3559]  & (~\all_features[3558]  | (~\all_features[3556]  & ~\all_features[3557]  & ~new_n11530_));
  assign new_n11541_ = ~new_n11542_ & (\all_features[3555]  | \all_features[3556]  | \all_features[3557]  | \all_features[3558]  | \all_features[3559] );
  assign new_n11542_ = ~new_n11534_ & (new_n11537_ | (~new_n11538_ & (new_n11540_ | (~new_n11539_ & ~new_n11543_))));
  assign new_n11543_ = ~new_n11527_ & (new_n11529_ | (new_n11532_ & (~new_n11531_ | (~new_n11544_ & new_n11520_))));
  assign new_n11544_ = ~\all_features[3557]  & \all_features[3558]  & \all_features[3559]  & (\all_features[3556]  ? new_n11524_ : (new_n11523_ | ~new_n11524_));
  assign new_n11545_ = new_n11546_ & new_n11533_ & ~new_n11538_ & ~new_n11539_ & ~new_n11527_ & ~new_n11537_;
  assign new_n11546_ = ~new_n11529_ & ~new_n11540_;
  assign new_n11547_ = new_n11533_ & new_n11536_ & (new_n11548_ | new_n11527_ | new_n11539_ | ~new_n11546_);
  assign new_n11548_ = new_n11532_ & new_n11522_ & new_n11531_ & new_n11520_;
  assign new_n11549_ = new_n10539_ & (~new_n10569_ | ~new_n10565_);
  assign new_n11550_ = new_n11551_ & new_n11573_;
  assign new_n11551_ = new_n11552_ & (~new_n11561_ | (new_n11571_ & new_n11572_ & new_n11568_ & new_n11570_));
  assign new_n11552_ = new_n11553_ & ~new_n11557_ & ~new_n11558_;
  assign new_n11553_ = ~new_n11554_ & (\all_features[2963]  | \all_features[2964]  | \all_features[2965]  | \all_features[2966]  | \all_features[2967] );
  assign new_n11554_ = ~\all_features[2965]  & new_n11556_ & ((~\all_features[2962]  & new_n11555_) | ~\all_features[2964]  | ~\all_features[2963] );
  assign new_n11555_ = ~\all_features[2960]  & ~\all_features[2961] ;
  assign new_n11556_ = ~\all_features[2966]  & ~\all_features[2967] ;
  assign new_n11557_ = new_n11556_ & (~\all_features[2965]  | (~\all_features[2964]  & (~\all_features[2963]  | (~\all_features[2962]  & ~\all_features[2961] ))));
  assign new_n11558_ = new_n11556_ & (~\all_features[2963]  | ~new_n11559_ | (~\all_features[2962]  & ~new_n11560_));
  assign new_n11559_ = \all_features[2964]  & \all_features[2965] ;
  assign new_n11560_ = \all_features[2960]  & \all_features[2961] ;
  assign new_n11561_ = ~new_n11567_ & ~new_n11566_ & ~new_n11562_ & ~new_n11564_;
  assign new_n11562_ = ~\all_features[2967]  & (~\all_features[2966]  | (~\all_features[2965]  & (new_n11555_ | ~new_n11563_ | ~\all_features[2964] )));
  assign new_n11563_ = \all_features[2962]  & \all_features[2963] ;
  assign new_n11564_ = ~new_n11565_ & ~\all_features[2967] ;
  assign new_n11565_ = \all_features[2965]  & \all_features[2966]  & (\all_features[2964]  | (\all_features[2962]  & \all_features[2963]  & \all_features[2961] ));
  assign new_n11566_ = ~\all_features[2967]  & (~\all_features[2966]  | ~new_n11559_ | ~new_n11560_ | ~new_n11563_);
  assign new_n11567_ = ~\all_features[2967]  & (~\all_features[2966]  | (~\all_features[2964]  & ~\all_features[2965]  & ~new_n11563_));
  assign new_n11568_ = \all_features[2967]  & (\all_features[2966]  | (\all_features[2965]  & (\all_features[2964]  | ~new_n11555_ | ~new_n11569_)));
  assign new_n11569_ = ~\all_features[2962]  & ~\all_features[2963] ;
  assign new_n11570_ = \all_features[2967]  & (\all_features[2966]  | (new_n11559_ & (\all_features[2962]  | \all_features[2963]  | \all_features[2961] )));
  assign new_n11571_ = \all_features[2966]  & \all_features[2967]  & (\all_features[2964]  | \all_features[2965]  | new_n11560_ | ~new_n11569_);
  assign new_n11572_ = \all_features[2967]  & (\all_features[2965]  | \all_features[2966]  | \all_features[2964] );
  assign new_n11573_ = new_n11552_ & new_n11561_;
  assign new_n11574_ = new_n11575_ ? new_n11613_ : ((new_n11704_ | ~new_n11635_ | new_n11673_) & (~new_n11633_ | ~new_n11673_));
  assign new_n11575_ = new_n11576_ & new_n11608_;
  assign new_n11576_ = new_n11577_ & new_n11598_;
  assign new_n11577_ = ~new_n11578_ & (\all_features[3731]  | \all_features[3732]  | \all_features[3733]  | \all_features[3734]  | \all_features[3735] );
  assign new_n11578_ = ~new_n11592_ & (new_n11594_ | (~new_n11595_ & (new_n11596_ | (~new_n11579_ & ~new_n11597_))));
  assign new_n11579_ = ~new_n11587_ & (new_n11589_ | (~new_n11580_ & new_n11591_));
  assign new_n11580_ = \all_features[3735]  & ((~new_n11585_ & ~\all_features[3733]  & \all_features[3734] ) | (~new_n11583_ & (\all_features[3734]  | (~new_n11581_ & \all_features[3733] ))));
  assign new_n11581_ = new_n11582_ & ~\all_features[3732]  & ~\all_features[3730]  & ~\all_features[3731] ;
  assign new_n11582_ = ~\all_features[3728]  & ~\all_features[3729] ;
  assign new_n11583_ = \all_features[3735]  & (\all_features[3734]  | (new_n11584_ & (\all_features[3730]  | \all_features[3731]  | \all_features[3729] )));
  assign new_n11584_ = \all_features[3732]  & \all_features[3733] ;
  assign new_n11585_ = (\all_features[3732]  & (\all_features[3730]  | \all_features[3731] )) | (~new_n11586_ & ~\all_features[3730]  & ~\all_features[3731]  & ~\all_features[3732] );
  assign new_n11586_ = \all_features[3728]  & \all_features[3729] ;
  assign new_n11587_ = ~new_n11588_ & ~\all_features[3735] ;
  assign new_n11588_ = \all_features[3733]  & \all_features[3734]  & (\all_features[3732]  | (\all_features[3730]  & \all_features[3731]  & \all_features[3729] ));
  assign new_n11589_ = ~\all_features[3735]  & (~\all_features[3734]  | ~new_n11586_ | ~new_n11584_ | ~new_n11590_);
  assign new_n11590_ = \all_features[3730]  & \all_features[3731] ;
  assign new_n11591_ = \all_features[3735]  & (\all_features[3733]  | \all_features[3734]  | \all_features[3732] );
  assign new_n11592_ = ~\all_features[3733]  & new_n11593_ & ((~\all_features[3730]  & new_n11582_) | ~\all_features[3732]  | ~\all_features[3731] );
  assign new_n11593_ = ~\all_features[3734]  & ~\all_features[3735] ;
  assign new_n11594_ = new_n11593_ & (~\all_features[3733]  | (~\all_features[3732]  & (~\all_features[3731]  | (~\all_features[3730]  & ~\all_features[3729] ))));
  assign new_n11595_ = new_n11593_ & (~\all_features[3731]  | ~new_n11584_ | (~\all_features[3730]  & ~new_n11586_));
  assign new_n11596_ = ~\all_features[3735]  & (~\all_features[3734]  | (~\all_features[3732]  & ~\all_features[3733]  & ~new_n11590_));
  assign new_n11597_ = ~\all_features[3735]  & (~\all_features[3734]  | (~\all_features[3733]  & (new_n11582_ | ~new_n11590_ | ~\all_features[3732] )));
  assign new_n11598_ = new_n11604_ & (~new_n11605_ | (new_n11606_ & (~new_n11607_ | new_n11599_)));
  assign new_n11599_ = new_n11600_ & (~new_n11601_ | (~new_n11603_ & \all_features[3733]  & \all_features[3734]  & \all_features[3735] ));
  assign new_n11600_ = \all_features[3735]  & (\all_features[3734]  | (~new_n11581_ & \all_features[3733] ));
  assign new_n11601_ = \all_features[3735]  & \all_features[3734]  & ~new_n11602_ & new_n11583_;
  assign new_n11602_ = ~\all_features[3733]  & ~\all_features[3732]  & ~\all_features[3731]  & ~new_n11586_ & ~\all_features[3730] ;
  assign new_n11603_ = ~\all_features[3731]  & ~\all_features[3732]  & (~\all_features[3730]  | new_n11582_);
  assign new_n11604_ = ~new_n11592_ & (\all_features[3731]  | \all_features[3732]  | \all_features[3733]  | \all_features[3734]  | \all_features[3735] );
  assign new_n11605_ = ~new_n11594_ & ~new_n11595_;
  assign new_n11606_ = ~new_n11596_ & ~new_n11597_;
  assign new_n11607_ = ~new_n11587_ & ~new_n11589_;
  assign new_n11608_ = new_n11609_ & new_n11612_;
  assign new_n11609_ = new_n11610_ & (new_n11597_ | new_n11587_ | ~new_n11611_ | (new_n11601_ & new_n11600_));
  assign new_n11610_ = new_n11604_ & new_n11605_;
  assign new_n11611_ = ~new_n11596_ & ~new_n11589_;
  assign new_n11612_ = new_n11607_ & new_n11610_ & new_n11606_;
  assign new_n11613_ = (~new_n8388_ & new_n11622_ & ~new_n11621_) | (new_n11621_ & (new_n11614_ | (new_n11629_ & new_n7040_)));
  assign new_n11614_ = new_n11615_ & new_n11616_;
  assign new_n11615_ = ~new_n7164_ & ~new_n7192_;
  assign new_n11616_ = ~new_n7188_ & ~new_n11617_;
  assign new_n11617_ = ~new_n7170_ & (new_n7167_ | (~new_n7171_ & ~new_n11618_));
  assign new_n11618_ = ~new_n7172_ & (new_n7185_ | (~new_n7180_ & (new_n7182_ | (~new_n7184_ & ~new_n11619_))));
  assign new_n11619_ = new_n7178_ & (~new_n7176_ | (new_n7187_ & (new_n11620_ | ~new_n7186_)));
  assign new_n11620_ = \all_features[3646]  & \all_features[3647]  & (\all_features[3645]  | (~new_n7177_ & \all_features[3644] ));
  assign new_n11621_ = ~new_n11172_ & new_n11201_;
  assign new_n11622_ = new_n8962_ & new_n11623_;
  assign new_n11623_ = new_n8987_ & new_n11624_;
  assign new_n11624_ = ~new_n8981_ & (new_n8979_ | (~new_n8984_ & (new_n8983_ | (~new_n11625_ & ~new_n8977_))));
  assign new_n11625_ = ~new_n8972_ & (new_n8974_ | (~new_n8976_ & (~new_n11628_ | new_n11626_)));
  assign new_n11626_ = \all_features[1687]  & ((~new_n11627_ & ~\all_features[1685]  & \all_features[1686] ) | (~new_n8969_ & (\all_features[1686]  | (~new_n8966_ & \all_features[1685] ))));
  assign new_n11627_ = (~\all_features[1682]  & ~\all_features[1683]  & ~\all_features[1684]  & (~\all_features[1681]  | ~\all_features[1680] )) | (\all_features[1684]  & (\all_features[1682]  | \all_features[1683] ));
  assign new_n11628_ = \all_features[1687]  & (\all_features[1685]  | \all_features[1686]  | \all_features[1684] );
  assign new_n11629_ = new_n7043_ & (new_n7048_ | new_n7047_ | (~new_n7052_ & ~new_n7057_ & ~new_n11630_));
  assign new_n11630_ = ~new_n7056_ & ~new_n7054_ & (~new_n7062_ | ~new_n7058_ | new_n11631_);
  assign new_n11631_ = new_n7060_ & new_n7061_ & (new_n11632_ | ~\all_features[3077]  | ~\all_features[3078]  | ~\all_features[3079] );
  assign new_n11632_ = ~\all_features[3075]  & ~\all_features[3076]  & (~\all_features[3074]  | new_n7045_);
  assign new_n11633_ = new_n8854_ & (new_n8851_ | new_n11634_);
  assign new_n11634_ = new_n8820_ & new_n8841_;
  assign new_n11635_ = new_n11636_ & new_n11668_;
  assign new_n11636_ = new_n11637_ & new_n11658_;
  assign new_n11637_ = ~new_n11638_ & (\all_features[4171]  | \all_features[4172]  | \all_features[4173]  | \all_features[4174]  | \all_features[4175] );
  assign new_n11638_ = ~new_n11652_ & (new_n11654_ | (~new_n11655_ & (new_n11656_ | (~new_n11639_ & ~new_n11657_))));
  assign new_n11639_ = ~new_n11647_ & (new_n11649_ | (~new_n11640_ & new_n11651_));
  assign new_n11640_ = \all_features[4175]  & ((~new_n11645_ & ~\all_features[4173]  & \all_features[4174] ) | (~new_n11643_ & (\all_features[4174]  | (~new_n11641_ & \all_features[4173] ))));
  assign new_n11641_ = new_n11642_ & ~\all_features[4172]  & ~\all_features[4170]  & ~\all_features[4171] ;
  assign new_n11642_ = ~\all_features[4168]  & ~\all_features[4169] ;
  assign new_n11643_ = \all_features[4175]  & (\all_features[4174]  | (new_n11644_ & (\all_features[4170]  | \all_features[4171]  | \all_features[4169] )));
  assign new_n11644_ = \all_features[4172]  & \all_features[4173] ;
  assign new_n11645_ = (\all_features[4172]  & (\all_features[4170]  | \all_features[4171] )) | (~new_n11646_ & ~\all_features[4170]  & ~\all_features[4171]  & ~\all_features[4172] );
  assign new_n11646_ = \all_features[4168]  & \all_features[4169] ;
  assign new_n11647_ = ~new_n11648_ & ~\all_features[4175] ;
  assign new_n11648_ = \all_features[4173]  & \all_features[4174]  & (\all_features[4172]  | (\all_features[4170]  & \all_features[4171]  & \all_features[4169] ));
  assign new_n11649_ = ~\all_features[4175]  & (~\all_features[4174]  | ~new_n11646_ | ~new_n11644_ | ~new_n11650_);
  assign new_n11650_ = \all_features[4170]  & \all_features[4171] ;
  assign new_n11651_ = \all_features[4175]  & (\all_features[4173]  | \all_features[4174]  | \all_features[4172] );
  assign new_n11652_ = ~\all_features[4173]  & new_n11653_ & ((~\all_features[4170]  & new_n11642_) | ~\all_features[4172]  | ~\all_features[4171] );
  assign new_n11653_ = ~\all_features[4174]  & ~\all_features[4175] ;
  assign new_n11654_ = new_n11653_ & (~\all_features[4173]  | (~\all_features[4172]  & (~\all_features[4171]  | (~\all_features[4170]  & ~\all_features[4169] ))));
  assign new_n11655_ = new_n11653_ & (~\all_features[4171]  | ~new_n11644_ | (~\all_features[4170]  & ~new_n11646_));
  assign new_n11656_ = ~\all_features[4175]  & (~\all_features[4174]  | (~\all_features[4172]  & ~\all_features[4173]  & ~new_n11650_));
  assign new_n11657_ = ~\all_features[4175]  & (~\all_features[4174]  | (~\all_features[4173]  & (new_n11642_ | ~new_n11650_ | ~\all_features[4172] )));
  assign new_n11658_ = new_n11664_ & (~new_n11665_ | (new_n11666_ & (~new_n11667_ | new_n11659_)));
  assign new_n11659_ = new_n11660_ & (~new_n11661_ | (~new_n11663_ & \all_features[4173]  & \all_features[4174]  & \all_features[4175] ));
  assign new_n11660_ = \all_features[4175]  & (\all_features[4174]  | (~new_n11641_ & \all_features[4173] ));
  assign new_n11661_ = \all_features[4175]  & \all_features[4174]  & ~new_n11662_ & new_n11643_;
  assign new_n11662_ = ~\all_features[4173]  & ~\all_features[4172]  & ~\all_features[4171]  & ~new_n11646_ & ~\all_features[4170] ;
  assign new_n11663_ = ~\all_features[4171]  & ~\all_features[4172]  & (~\all_features[4170]  | new_n11642_);
  assign new_n11664_ = ~new_n11652_ & (\all_features[4171]  | \all_features[4172]  | \all_features[4173]  | \all_features[4174]  | \all_features[4175] );
  assign new_n11665_ = ~new_n11654_ & ~new_n11655_;
  assign new_n11666_ = ~new_n11656_ & ~new_n11657_;
  assign new_n11667_ = ~new_n11647_ & ~new_n11649_;
  assign new_n11668_ = new_n11669_ & new_n11672_;
  assign new_n11669_ = new_n11670_ & (new_n11657_ | new_n11647_ | ~new_n11671_ | (new_n11661_ & new_n11660_));
  assign new_n11670_ = new_n11664_ & new_n11665_;
  assign new_n11671_ = ~new_n11656_ & ~new_n11649_;
  assign new_n11672_ = new_n11667_ & new_n11670_ & new_n11666_;
  assign new_n11673_ = new_n11674_ & new_n11700_;
  assign new_n11674_ = new_n11675_ & new_n11699_;
  assign new_n11675_ = new_n11693_ & ~new_n11698_ & ~new_n11676_ & ~new_n11697_;
  assign new_n11676_ = ~new_n11686_ & ~new_n11692_ & new_n11682_ & (~new_n11690_ | ~new_n11688_ | ~new_n11677_);
  assign new_n11677_ = new_n11678_ & new_n11681_;
  assign new_n11678_ = \all_features[3639]  & (\all_features[3638]  | (\all_features[3637]  & (\all_features[3636]  | ~new_n11680_ | ~new_n11679_)));
  assign new_n11679_ = ~\all_features[3634]  & ~\all_features[3635] ;
  assign new_n11680_ = ~\all_features[3632]  & ~\all_features[3633] ;
  assign new_n11681_ = \all_features[3639]  & (\all_features[3637]  | \all_features[3638]  | \all_features[3636] );
  assign new_n11682_ = ~new_n11683_ & ~new_n11685_;
  assign new_n11683_ = ~new_n11684_ & ~\all_features[3639] ;
  assign new_n11684_ = \all_features[3637]  & \all_features[3638]  & (\all_features[3636]  | (\all_features[3634]  & \all_features[3635]  & \all_features[3633] ));
  assign new_n11685_ = ~\all_features[3639]  & (~\all_features[3638]  | (~\all_features[3637]  & ~\all_features[3636]  & (~\all_features[3635]  | ~\all_features[3634] )));
  assign new_n11686_ = ~\all_features[3639]  & (~\all_features[3638]  | new_n11687_);
  assign new_n11687_ = ~\all_features[3637]  & (new_n11680_ | ~\all_features[3635]  | ~\all_features[3636]  | ~\all_features[3634] );
  assign new_n11688_ = \all_features[3638]  & \all_features[3639]  & (\all_features[3636]  | \all_features[3637]  | new_n11689_ | ~new_n11679_);
  assign new_n11689_ = \all_features[3632]  & \all_features[3633] ;
  assign new_n11690_ = \all_features[3639]  & (\all_features[3638]  | (new_n11691_ & (\all_features[3634]  | \all_features[3635]  | \all_features[3633] )));
  assign new_n11691_ = \all_features[3636]  & \all_features[3637] ;
  assign new_n11692_ = ~\all_features[3639]  & (~new_n11691_ | ~\all_features[3634]  | ~\all_features[3635]  | ~\all_features[3638]  | ~new_n11689_);
  assign new_n11693_ = ~new_n11694_ & ~new_n11696_;
  assign new_n11694_ = ~\all_features[3637]  & new_n11695_ & ((~\all_features[3634]  & new_n11680_) | ~\all_features[3636]  | ~\all_features[3635] );
  assign new_n11695_ = ~\all_features[3638]  & ~\all_features[3639] ;
  assign new_n11696_ = ~\all_features[3639]  & ~\all_features[3638]  & ~\all_features[3637]  & ~\all_features[3635]  & ~\all_features[3636] ;
  assign new_n11697_ = new_n11695_ & (~\all_features[3637]  | (~\all_features[3636]  & (~\all_features[3635]  | (~\all_features[3634]  & ~\all_features[3633] ))));
  assign new_n11698_ = new_n11695_ & (~\all_features[3635]  | ~new_n11691_ | (~\all_features[3634]  & ~new_n11689_));
  assign new_n11699_ = new_n11682_ & new_n11693_ & ~new_n11698_ & ~new_n11697_ & ~new_n11686_ & ~new_n11692_;
  assign new_n11700_ = new_n11693_ & (new_n11698_ | new_n11697_ | (~new_n11701_ & ~new_n11686_ & ~new_n11685_));
  assign new_n11701_ = ~new_n11683_ & ~new_n11692_ & (~new_n11677_ | (~new_n11702_ & new_n11688_ & new_n11690_));
  assign new_n11702_ = \all_features[3639]  & \all_features[3638]  & ~new_n11703_ & \all_features[3637] ;
  assign new_n11703_ = ~\all_features[3635]  & ~\all_features[3636]  & (~\all_features[3634]  | new_n11680_);
  assign new_n11704_ = new_n11710_ & new_n11705_ & ~new_n11720_ & ~new_n11719_ & ~new_n11716_ & ~new_n11718_;
  assign new_n11705_ = ~new_n11706_ & ~new_n11709_;
  assign new_n11706_ = ~\all_features[3541]  & new_n11707_ & ((~\all_features[3538]  & new_n11708_) | ~\all_features[3540]  | ~\all_features[3539] );
  assign new_n11707_ = ~\all_features[3542]  & ~\all_features[3543] ;
  assign new_n11708_ = ~\all_features[3536]  & ~\all_features[3537] ;
  assign new_n11709_ = ~\all_features[3543]  & ~\all_features[3542]  & ~\all_features[3541]  & ~\all_features[3539]  & ~\all_features[3540] ;
  assign new_n11710_ = ~new_n11711_ & ~new_n11715_;
  assign new_n11711_ = ~\all_features[3543]  & (~\all_features[3542]  | ~new_n11712_ | ~new_n11713_ | ~new_n11714_);
  assign new_n11712_ = \all_features[3538]  & \all_features[3539] ;
  assign new_n11713_ = \all_features[3536]  & \all_features[3537] ;
  assign new_n11714_ = \all_features[3540]  & \all_features[3541] ;
  assign new_n11715_ = ~\all_features[3543]  & (~\all_features[3542]  | (~\all_features[3540]  & ~\all_features[3541]  & ~new_n11712_));
  assign new_n11716_ = ~new_n11717_ & ~\all_features[3543] ;
  assign new_n11717_ = \all_features[3541]  & \all_features[3542]  & (\all_features[3540]  | (\all_features[3538]  & \all_features[3539]  & \all_features[3537] ));
  assign new_n11718_ = new_n11707_ & (~\all_features[3541]  | (~\all_features[3540]  & (~\all_features[3539]  | (~\all_features[3538]  & ~\all_features[3537] ))));
  assign new_n11719_ = ~\all_features[3543]  & (~\all_features[3542]  | (~\all_features[3541]  & (new_n11708_ | ~new_n11712_ | ~\all_features[3540] )));
  assign new_n11720_ = new_n11707_ & (~\all_features[3539]  | ~new_n11714_ | (~\all_features[3538]  & ~new_n11713_));
  assign new_n11721_ = ~new_n11722_ & new_n12039_;
  assign new_n11722_ = new_n11723_ & (~new_n11901_ | new_n11941_);
  assign new_n11723_ = new_n11724_ & (new_n11897_ | new_n11901_ | (new_n11902_ ? new_n11905_ : ~new_n11907_));
  assign new_n11724_ = (~new_n11897_ | new_n11755_ | new_n11901_) & (new_n11725_ | ~new_n11895_ | ~new_n11859_ | ~new_n11901_);
  assign new_n11725_ = ~new_n11751_ & new_n11726_;
  assign new_n11726_ = ~new_n11727_ & ~new_n11750_;
  assign new_n11727_ = new_n11728_ & (~new_n11740_ | (new_n11737_ & new_n11748_));
  assign new_n11728_ = new_n11729_ & new_n11733_;
  assign new_n11729_ = ~new_n11730_ & (\all_features[4619]  | \all_features[4620]  | ~new_n11731_);
  assign new_n11730_ = new_n11731_ & ((~\all_features[4617]  & ~\all_features[4618]  & ~\all_features[4616] ) | ~\all_features[4620]  | ~\all_features[4619] );
  assign new_n11731_ = ~\all_features[4621]  & new_n11732_;
  assign new_n11732_ = ~\all_features[4622]  & ~\all_features[4623] ;
  assign new_n11733_ = ~new_n11734_ & ~new_n11736_;
  assign new_n11734_ = new_n11732_ & (~new_n11735_ | ~\all_features[4619]  | (~\all_features[4618]  & (~\all_features[4616]  | ~\all_features[4617] )));
  assign new_n11735_ = \all_features[4620]  & \all_features[4621] ;
  assign new_n11736_ = new_n11732_ & (~\all_features[4621]  | (~\all_features[4620]  & (~\all_features[4619]  | (~\all_features[4618]  & ~\all_features[4617] ))));
  assign new_n11737_ = \all_features[4623]  & \all_features[4622]  & ~new_n11739_ & new_n11738_;
  assign new_n11738_ = \all_features[4623]  & (\all_features[4622]  | (new_n11735_ & (\all_features[4618]  | \all_features[4619]  | \all_features[4617] )));
  assign new_n11739_ = ~\all_features[4618]  & ~\all_features[4619]  & ~\all_features[4620]  & ~\all_features[4621]  & (~\all_features[4617]  | ~\all_features[4616] );
  assign new_n11740_ = ~new_n11747_ & ~new_n11745_ & ~new_n11741_ & ~new_n11743_;
  assign new_n11741_ = ~new_n11742_ & ~\all_features[4623] ;
  assign new_n11742_ = \all_features[4621]  & \all_features[4622]  & (\all_features[4620]  | (\all_features[4618]  & \all_features[4619]  & \all_features[4617] ));
  assign new_n11743_ = ~\all_features[4623]  & (~\all_features[4619]  | ~new_n11735_ | ~new_n11744_ | ~\all_features[4618] );
  assign new_n11744_ = \all_features[4622]  & \all_features[4616]  & \all_features[4617] ;
  assign new_n11745_ = ~\all_features[4623]  & (~\all_features[4622]  | new_n11746_);
  assign new_n11746_ = ~\all_features[4621]  & (~\all_features[4619]  | ~\all_features[4620]  | ~\all_features[4618]  | (~\all_features[4617]  & ~\all_features[4616] ));
  assign new_n11747_ = ~\all_features[4623]  & (~\all_features[4622]  | (~\all_features[4621]  & ~\all_features[4620]  & (~\all_features[4619]  | ~\all_features[4618] )));
  assign new_n11748_ = \all_features[4623]  & (\all_features[4622]  | (~new_n11749_ & \all_features[4621] ));
  assign new_n11749_ = ~\all_features[4620]  & ~\all_features[4619]  & ~\all_features[4618]  & ~\all_features[4616]  & ~\all_features[4617] ;
  assign new_n11750_ = new_n11728_ & new_n11740_;
  assign new_n11751_ = new_n11729_ & (~new_n11733_ | (~new_n11752_ & ~new_n11745_ & ~new_n11747_));
  assign new_n11752_ = ~new_n11741_ & ~new_n11743_ & (~new_n11748_ | (~new_n11753_ & new_n11737_));
  assign new_n11753_ = \all_features[4623]  & \all_features[4622]  & ~new_n11754_ & \all_features[4621] ;
  assign new_n11754_ = ~\all_features[4619]  & ~\all_features[4620]  & (~\all_features[4618]  | (~\all_features[4617]  & ~\all_features[4616] ));
  assign new_n11755_ = new_n11756_ ? ~new_n11824_ : ~new_n11792_;
  assign new_n11756_ = new_n11757_ & new_n11783_;
  assign new_n11757_ = ~new_n11758_ & ~new_n11781_;
  assign new_n11758_ = new_n11776_ & ~new_n11780_ & ~new_n11759_ & ~new_n11779_;
  assign new_n11759_ = ~new_n11774_ & ~new_n11775_ & new_n11767_ & (~new_n11772_ | ~new_n11760_);
  assign new_n11760_ = new_n11766_ & new_n11761_ & new_n11763_;
  assign new_n11761_ = \all_features[5519]  & (\all_features[5518]  | (new_n11762_ & (\all_features[5514]  | \all_features[5515]  | \all_features[5513] )));
  assign new_n11762_ = \all_features[5516]  & \all_features[5517] ;
  assign new_n11763_ = \all_features[5518]  & \all_features[5519]  & (\all_features[5516]  | \all_features[5517]  | new_n11765_ | ~new_n11764_);
  assign new_n11764_ = ~\all_features[5514]  & ~\all_features[5515] ;
  assign new_n11765_ = \all_features[5512]  & \all_features[5513] ;
  assign new_n11766_ = \all_features[5519]  & (\all_features[5517]  | \all_features[5518]  | \all_features[5516] );
  assign new_n11767_ = ~new_n11768_ & ~new_n11770_;
  assign new_n11768_ = ~new_n11769_ & ~\all_features[5519] ;
  assign new_n11769_ = \all_features[5517]  & \all_features[5518]  & (\all_features[5516]  | (\all_features[5514]  & \all_features[5515]  & \all_features[5513] ));
  assign new_n11770_ = ~\all_features[5519]  & (~\all_features[5518]  | (~\all_features[5516]  & ~\all_features[5517]  & ~new_n11771_));
  assign new_n11771_ = \all_features[5514]  & \all_features[5515] ;
  assign new_n11772_ = \all_features[5519]  & (\all_features[5518]  | (\all_features[5517]  & (\all_features[5516]  | ~new_n11773_ | ~new_n11764_)));
  assign new_n11773_ = ~\all_features[5512]  & ~\all_features[5513] ;
  assign new_n11774_ = ~\all_features[5519]  & (~\all_features[5518]  | (~\all_features[5517]  & (new_n11773_ | ~new_n11771_ | ~\all_features[5516] )));
  assign new_n11775_ = ~\all_features[5519]  & (~\all_features[5518]  | ~new_n11762_ | ~new_n11765_ | ~new_n11771_);
  assign new_n11776_ = ~new_n11777_ & (\all_features[5515]  | \all_features[5516]  | \all_features[5517]  | \all_features[5518]  | \all_features[5519] );
  assign new_n11777_ = ~\all_features[5517]  & new_n11778_ & ((~\all_features[5514]  & new_n11773_) | ~\all_features[5516]  | ~\all_features[5515] );
  assign new_n11778_ = ~\all_features[5518]  & ~\all_features[5519] ;
  assign new_n11779_ = new_n11778_ & (~\all_features[5517]  | (~\all_features[5516]  & (~\all_features[5515]  | (~\all_features[5514]  & ~\all_features[5513] ))));
  assign new_n11780_ = new_n11778_ & (~\all_features[5515]  | ~new_n11762_ | (~\all_features[5514]  & ~new_n11765_));
  assign new_n11781_ = new_n11776_ & new_n11767_ & new_n11782_ & ~new_n11774_ & ~new_n11775_;
  assign new_n11782_ = ~new_n11779_ & ~new_n11780_;
  assign new_n11783_ = ~new_n11784_ & ~new_n11788_;
  assign new_n11784_ = new_n11776_ & (~new_n11782_ | (~new_n11785_ & ~new_n11770_ & ~new_n11774_));
  assign new_n11785_ = ~new_n11775_ & ~new_n11768_ & (~new_n11766_ | ~new_n11772_ | new_n11786_);
  assign new_n11786_ = new_n11761_ & new_n11763_ & (new_n11787_ | ~\all_features[5517]  | ~\all_features[5518]  | ~\all_features[5519] );
  assign new_n11787_ = ~\all_features[5515]  & ~\all_features[5516]  & (~\all_features[5514]  | new_n11773_);
  assign new_n11788_ = ~new_n11789_ & (\all_features[5515]  | \all_features[5516]  | \all_features[5517]  | \all_features[5518]  | \all_features[5519] );
  assign new_n11789_ = ~new_n11777_ & (new_n11779_ | (~new_n11780_ & (new_n11770_ | (~new_n11774_ & ~new_n11790_))));
  assign new_n11790_ = ~new_n11768_ & (new_n11775_ | (new_n11766_ & (~new_n11772_ | (~new_n11791_ & new_n11761_))));
  assign new_n11791_ = ~\all_features[5517]  & \all_features[5518]  & \all_features[5519]  & (\all_features[5516]  ? new_n11764_ : (new_n11765_ | ~new_n11764_));
  assign new_n11792_ = ~new_n11793_ & new_n11823_;
  assign new_n11793_ = ~new_n11794_ & ~new_n11820_;
  assign new_n11794_ = new_n11806_ & (~new_n11809_ | (new_n11812_ & (~new_n11816_ | new_n11795_)));
  assign new_n11795_ = new_n11796_ & (~new_n11801_ | (~new_n11805_ & \all_features[1445]  & \all_features[1446]  & \all_features[1447] ));
  assign new_n11796_ = \all_features[1447]  & (\all_features[1446]  | (~new_n11800_ & new_n11797_));
  assign new_n11797_ = \all_features[1445]  & (\all_features[1444]  | ~new_n11799_ | ~new_n11798_);
  assign new_n11798_ = ~\all_features[1440]  & ~\all_features[1441] ;
  assign new_n11799_ = ~\all_features[1442]  & ~\all_features[1443] ;
  assign new_n11800_ = ~\all_features[1444]  & ~\all_features[1445] ;
  assign new_n11801_ = new_n11802_ & \all_features[1446]  & \all_features[1447]  & (~new_n11799_ | ~new_n11800_ | new_n11804_);
  assign new_n11802_ = \all_features[1447]  & (\all_features[1446]  | (new_n11803_ & (\all_features[1442]  | \all_features[1443]  | \all_features[1441] )));
  assign new_n11803_ = \all_features[1444]  & \all_features[1445] ;
  assign new_n11804_ = \all_features[1440]  & \all_features[1441] ;
  assign new_n11805_ = ~\all_features[1443]  & ~\all_features[1444]  & (~\all_features[1442]  | new_n11798_);
  assign new_n11806_ = ~new_n11807_ & (\all_features[1443]  | \all_features[1444]  | \all_features[1445]  | \all_features[1446]  | \all_features[1447] );
  assign new_n11807_ = ~\all_features[1445]  & new_n11808_ & ((~\all_features[1442]  & new_n11798_) | ~\all_features[1444]  | ~\all_features[1443] );
  assign new_n11808_ = ~\all_features[1446]  & ~\all_features[1447] ;
  assign new_n11809_ = ~new_n11810_ & ~new_n11811_;
  assign new_n11810_ = new_n11808_ & (~\all_features[1443]  | ~new_n11803_ | (~\all_features[1442]  & ~new_n11804_));
  assign new_n11811_ = new_n11808_ & (~\all_features[1445]  | (~\all_features[1444]  & (~\all_features[1443]  | (~\all_features[1442]  & ~\all_features[1441] ))));
  assign new_n11812_ = ~new_n11813_ & ~new_n11815_;
  assign new_n11813_ = ~\all_features[1447]  & (~\all_features[1446]  | (~new_n11814_ & new_n11800_));
  assign new_n11814_ = \all_features[1442]  & \all_features[1443] ;
  assign new_n11815_ = ~\all_features[1447]  & (~\all_features[1446]  | (~\all_features[1445]  & (new_n11798_ | ~new_n11814_ | ~\all_features[1444] )));
  assign new_n11816_ = ~new_n11817_ & ~new_n11818_;
  assign new_n11817_ = ~\all_features[1447]  & (~\all_features[1446]  | ~new_n11804_ | ~new_n11803_ | ~new_n11814_);
  assign new_n11818_ = ~new_n11819_ & ~\all_features[1447] ;
  assign new_n11819_ = \all_features[1445]  & \all_features[1446]  & (\all_features[1444]  | (\all_features[1442]  & \all_features[1443]  & \all_features[1441] ));
  assign new_n11820_ = new_n11821_ & (new_n11815_ | new_n11818_ | ~new_n11822_ | (new_n11801_ & new_n11796_));
  assign new_n11821_ = new_n11806_ & new_n11809_;
  assign new_n11822_ = ~new_n11813_ & ~new_n11817_;
  assign new_n11823_ = new_n11816_ & new_n11821_ & new_n11812_;
  assign new_n11824_ = ~new_n11857_ & ~new_n11846_ & ~new_n11854_ & (new_n11852_ | (~new_n11851_ & ~new_n11825_));
  assign new_n11825_ = ~new_n11839_ & (new_n11841_ | (~new_n11842_ & (new_n11843_ | (~new_n11826_ & ~new_n11844_))));
  assign new_n11826_ = ~new_n11833_ & (~new_n11837_ | (new_n11827_ & (~new_n11836_ | (~new_n11838_ & new_n11830_))));
  assign new_n11827_ = \all_features[5711]  & (\all_features[5710]  | new_n11828_);
  assign new_n11828_ = \all_features[5709]  & (\all_features[5706]  | \all_features[5707]  | \all_features[5708]  | ~new_n11829_);
  assign new_n11829_ = ~\all_features[5704]  & ~\all_features[5705] ;
  assign new_n11830_ = \all_features[5711]  & ~new_n11831_ & \all_features[5710] ;
  assign new_n11831_ = ~\all_features[5709]  & ~\all_features[5708]  & ~\all_features[5707]  & ~new_n11832_ & ~\all_features[5706] ;
  assign new_n11832_ = \all_features[5704]  & \all_features[5705] ;
  assign new_n11833_ = ~\all_features[5711]  & (~\all_features[5710]  | ~new_n11832_ | ~new_n11834_ | ~new_n11835_);
  assign new_n11834_ = \all_features[5708]  & \all_features[5709] ;
  assign new_n11835_ = \all_features[5706]  & \all_features[5707] ;
  assign new_n11836_ = \all_features[5711]  & (\all_features[5710]  | (new_n11834_ & (\all_features[5706]  | \all_features[5707]  | \all_features[5705] )));
  assign new_n11837_ = \all_features[5711]  & (\all_features[5709]  | \all_features[5710]  | \all_features[5708] );
  assign new_n11838_ = \all_features[5710]  & \all_features[5711]  & (\all_features[5709]  | (\all_features[5708]  & (\all_features[5707]  | \all_features[5706] )));
  assign new_n11839_ = new_n11840_ & (~\all_features[5709]  | (~\all_features[5708]  & (~\all_features[5707]  | (~\all_features[5706]  & ~\all_features[5705] ))));
  assign new_n11840_ = ~\all_features[5710]  & ~\all_features[5711] ;
  assign new_n11841_ = new_n11840_ & (~\all_features[5707]  | ~new_n11834_ | (~\all_features[5706]  & ~new_n11832_));
  assign new_n11842_ = ~\all_features[5711]  & (~\all_features[5710]  | (~\all_features[5708]  & ~\all_features[5709]  & ~new_n11835_));
  assign new_n11843_ = ~\all_features[5711]  & (~\all_features[5710]  | (~\all_features[5709]  & (new_n11829_ | ~new_n11835_ | ~\all_features[5708] )));
  assign new_n11844_ = ~new_n11845_ & ~\all_features[5711] ;
  assign new_n11845_ = \all_features[5709]  & \all_features[5710]  & (\all_features[5708]  | (\all_features[5706]  & \all_features[5707]  & \all_features[5705] ));
  assign new_n11846_ = new_n11850_ & (~new_n11853_ | (~new_n11847_ & ~new_n11842_ & ~new_n11843_));
  assign new_n11847_ = ~new_n11833_ & ~new_n11844_ & (~new_n11837_ | new_n11848_ | ~new_n11827_);
  assign new_n11848_ = ~new_n11831_ & new_n11836_ & \all_features[5710]  & \all_features[5711]  & (~\all_features[5709]  | new_n11849_);
  assign new_n11849_ = ~\all_features[5707]  & ~\all_features[5708]  & (~\all_features[5706]  | new_n11829_);
  assign new_n11850_ = ~new_n11851_ & ~new_n11852_;
  assign new_n11851_ = ~\all_features[5709]  & new_n11840_ & ((~\all_features[5706]  & new_n11829_) | ~\all_features[5708]  | ~\all_features[5707] );
  assign new_n11852_ = ~\all_features[5711]  & ~\all_features[5710]  & ~\all_features[5709]  & ~\all_features[5707]  & ~\all_features[5708] ;
  assign new_n11853_ = ~new_n11839_ & ~new_n11841_;
  assign new_n11854_ = new_n11853_ & ~new_n11855_ & new_n11850_;
  assign new_n11855_ = new_n11856_ & (~new_n11836_ | ~new_n11837_ | ~new_n11830_ | ~new_n11827_);
  assign new_n11856_ = ~new_n11833_ & ~new_n11844_ & ~new_n11842_ & ~new_n11843_;
  assign new_n11857_ = new_n11858_ & new_n11850_ & ~new_n11839_ & ~new_n11844_;
  assign new_n11858_ = ~new_n11833_ & ~new_n11843_ & ~new_n11841_ & ~new_n11842_;
  assign new_n11859_ = new_n11860_ & new_n11886_;
  assign new_n11860_ = new_n11861_ & new_n11884_;
  assign new_n11861_ = new_n11879_ & ~new_n11883_ & ~new_n11862_ & ~new_n11882_;
  assign new_n11862_ = ~new_n11877_ & ~new_n11878_ & new_n11870_ & (~new_n11875_ | ~new_n11863_);
  assign new_n11863_ = new_n11869_ & new_n11864_ & new_n11866_;
  assign new_n11864_ = \all_features[2799]  & (\all_features[2798]  | (new_n11865_ & (\all_features[2794]  | \all_features[2795]  | \all_features[2793] )));
  assign new_n11865_ = \all_features[2796]  & \all_features[2797] ;
  assign new_n11866_ = \all_features[2798]  & \all_features[2799]  & (\all_features[2796]  | \all_features[2797]  | new_n11868_ | ~new_n11867_);
  assign new_n11867_ = ~\all_features[2794]  & ~\all_features[2795] ;
  assign new_n11868_ = \all_features[2792]  & \all_features[2793] ;
  assign new_n11869_ = \all_features[2799]  & (\all_features[2797]  | \all_features[2798]  | \all_features[2796] );
  assign new_n11870_ = ~new_n11871_ & ~new_n11873_;
  assign new_n11871_ = ~new_n11872_ & ~\all_features[2799] ;
  assign new_n11872_ = \all_features[2797]  & \all_features[2798]  & (\all_features[2796]  | (\all_features[2794]  & \all_features[2795]  & \all_features[2793] ));
  assign new_n11873_ = ~\all_features[2799]  & (~\all_features[2798]  | (~\all_features[2796]  & ~\all_features[2797]  & ~new_n11874_));
  assign new_n11874_ = \all_features[2794]  & \all_features[2795] ;
  assign new_n11875_ = \all_features[2799]  & (\all_features[2798]  | (\all_features[2797]  & (\all_features[2796]  | ~new_n11876_ | ~new_n11867_)));
  assign new_n11876_ = ~\all_features[2792]  & ~\all_features[2793] ;
  assign new_n11877_ = ~\all_features[2799]  & (~\all_features[2798]  | (~\all_features[2797]  & (new_n11876_ | ~new_n11874_ | ~\all_features[2796] )));
  assign new_n11878_ = ~\all_features[2799]  & (~\all_features[2798]  | ~new_n11865_ | ~new_n11868_ | ~new_n11874_);
  assign new_n11879_ = ~new_n11880_ & (\all_features[2795]  | \all_features[2796]  | \all_features[2797]  | \all_features[2798]  | \all_features[2799] );
  assign new_n11880_ = ~\all_features[2797]  & new_n11881_ & ((~\all_features[2794]  & new_n11876_) | ~\all_features[2796]  | ~\all_features[2795] );
  assign new_n11881_ = ~\all_features[2798]  & ~\all_features[2799] ;
  assign new_n11882_ = new_n11881_ & (~\all_features[2797]  | (~\all_features[2796]  & (~\all_features[2795]  | (~\all_features[2794]  & ~\all_features[2793] ))));
  assign new_n11883_ = new_n11881_ & (~\all_features[2795]  | ~new_n11865_ | (~\all_features[2794]  & ~new_n11868_));
  assign new_n11884_ = new_n11879_ & new_n11870_ & new_n11885_ & ~new_n11877_ & ~new_n11878_;
  assign new_n11885_ = ~new_n11882_ & ~new_n11883_;
  assign new_n11886_ = new_n11887_ & new_n11891_;
  assign new_n11887_ = new_n11879_ & (~new_n11885_ | (~new_n11888_ & ~new_n11873_ & ~new_n11877_));
  assign new_n11888_ = ~new_n11878_ & ~new_n11871_ & (~new_n11869_ | ~new_n11875_ | new_n11889_);
  assign new_n11889_ = new_n11864_ & new_n11866_ & (new_n11890_ | ~\all_features[2797]  | ~\all_features[2798]  | ~\all_features[2799] );
  assign new_n11890_ = ~\all_features[2795]  & ~\all_features[2796]  & (~\all_features[2794]  | new_n11876_);
  assign new_n11891_ = ~new_n11892_ & (\all_features[2795]  | \all_features[2796]  | \all_features[2797]  | \all_features[2798]  | \all_features[2799] );
  assign new_n11892_ = ~new_n11880_ & (new_n11882_ | (~new_n11883_ & (new_n11873_ | (~new_n11877_ & ~new_n11893_))));
  assign new_n11893_ = ~new_n11871_ & (new_n11878_ | (new_n11869_ & (~new_n11875_ | (~new_n11894_ & new_n11864_))));
  assign new_n11894_ = ~\all_features[2797]  & \all_features[2798]  & \all_features[2799]  & (\all_features[2796]  ? new_n11867_ : (new_n11868_ | ~new_n11867_));
  assign new_n11895_ = new_n11896_ & new_n8295_;
  assign new_n11896_ = new_n8269_ & new_n8292_;
  assign new_n11897_ = new_n11471_ & (new_n11493_ | (~new_n11497_ & (new_n11494_ | (~new_n11898_ & ~new_n11496_))));
  assign new_n11898_ = ~new_n11487_ & (new_n11488_ | (~new_n11482_ & ~new_n11899_));
  assign new_n11899_ = ~new_n11484_ & (~new_n11490_ | (new_n11489_ & (~new_n11474_ | (~new_n11900_ & new_n11478_))));
  assign new_n11900_ = \all_features[5086]  & \all_features[5087]  & (\all_features[5085]  | (~new_n11479_ & \all_features[5084] ));
  assign new_n11901_ = new_n6563_ & new_n6566_;
  assign new_n11902_ = new_n11903_ & new_n11904_;
  assign new_n11903_ = ~new_n11577_ & ~new_n11598_;
  assign new_n11904_ = ~new_n11609_ & ~new_n11612_;
  assign new_n11905_ = new_n7446_ & new_n11906_;
  assign new_n11906_ = new_n7475_ & new_n7477_;
  assign new_n11907_ = new_n11940_ & (new_n11908_ | (new_n11931_ & new_n11935_));
  assign new_n11908_ = new_n11928_ & ~new_n11909_ & new_n11923_;
  assign new_n11909_ = ~new_n11917_ & ~new_n11919_ & ~new_n11920_ & ~new_n11922_ & (~new_n11914_ | ~new_n11910_);
  assign new_n11910_ = \all_features[999]  & \all_features[998]  & ~new_n11913_ & new_n11911_;
  assign new_n11911_ = \all_features[999]  & (\all_features[998]  | (new_n11912_ & (\all_features[994]  | \all_features[995]  | \all_features[993] )));
  assign new_n11912_ = \all_features[996]  & \all_features[997] ;
  assign new_n11913_ = ~\all_features[994]  & ~\all_features[995]  & ~\all_features[996]  & ~\all_features[997]  & (~\all_features[993]  | ~\all_features[992] );
  assign new_n11914_ = \all_features[999]  & (\all_features[998]  | (~new_n11915_ & \all_features[997] ));
  assign new_n11915_ = new_n11916_ & ~\all_features[996]  & ~\all_features[994]  & ~\all_features[995] ;
  assign new_n11916_ = ~\all_features[992]  & ~\all_features[993] ;
  assign new_n11917_ = ~\all_features[999]  & (~\all_features[998]  | (~\all_features[996]  & ~\all_features[997]  & ~new_n11918_));
  assign new_n11918_ = \all_features[994]  & \all_features[995] ;
  assign new_n11919_ = ~\all_features[999]  & (~\all_features[998]  | (~\all_features[997]  & (new_n11916_ | ~\all_features[996]  | ~new_n11918_)));
  assign new_n11920_ = ~new_n11921_ & ~\all_features[999] ;
  assign new_n11921_ = \all_features[997]  & \all_features[998]  & (\all_features[996]  | (\all_features[994]  & \all_features[995]  & \all_features[993] ));
  assign new_n11922_ = ~\all_features[999]  & (~new_n11912_ | ~\all_features[992]  | ~\all_features[993]  | ~\all_features[998]  | ~new_n11918_);
  assign new_n11923_ = ~new_n11924_ & ~new_n11927_;
  assign new_n11924_ = new_n11925_ & ((~\all_features[994]  & new_n11916_) | ~\all_features[996]  | ~\all_features[995] );
  assign new_n11925_ = ~\all_features[997]  & new_n11926_;
  assign new_n11926_ = ~\all_features[998]  & ~\all_features[999] ;
  assign new_n11927_ = new_n11925_ & ~\all_features[995]  & ~\all_features[996] ;
  assign new_n11928_ = ~new_n11929_ & ~new_n11930_;
  assign new_n11929_ = new_n11926_ & (~new_n11912_ | ~\all_features[995]  | (~\all_features[994]  & (~\all_features[992]  | ~\all_features[993] )));
  assign new_n11930_ = new_n11926_ & (~\all_features[997]  | (~\all_features[996]  & (~\all_features[995]  | (~\all_features[994]  & ~\all_features[993] ))));
  assign new_n11931_ = new_n11923_ & (~new_n11928_ | (new_n11934_ & (new_n11932_ | new_n11920_ | new_n11922_)));
  assign new_n11932_ = new_n11914_ & (~new_n11910_ | (~new_n11933_ & \all_features[997]  & \all_features[998]  & \all_features[999] ));
  assign new_n11933_ = ~\all_features[995]  & ~\all_features[996]  & (~\all_features[994]  | new_n11916_);
  assign new_n11934_ = ~new_n11917_ & ~new_n11919_;
  assign new_n11935_ = ~new_n11927_ & (new_n11924_ | (~new_n11930_ & (new_n11929_ | (~new_n11917_ & ~new_n11936_))));
  assign new_n11936_ = ~new_n11919_ & (new_n11920_ | (~new_n11922_ & (~new_n11939_ | new_n11937_)));
  assign new_n11937_ = \all_features[999]  & ((~new_n11938_ & ~\all_features[997]  & \all_features[998] ) | (~new_n11911_ & (\all_features[998]  | (~new_n11915_ & \all_features[997] ))));
  assign new_n11938_ = (~\all_features[994]  & ~\all_features[995]  & ~\all_features[996]  & (~\all_features[993]  | ~\all_features[992] )) | (\all_features[996]  & (\all_features[994]  | \all_features[995] ));
  assign new_n11939_ = \all_features[999]  & (\all_features[997]  | \all_features[998]  | \all_features[996] );
  assign new_n11940_ = new_n11928_ & new_n11934_ & ~new_n11922_ & ~new_n11920_ & ~new_n11924_ & ~new_n11927_;
  assign new_n11941_ = (~new_n11725_ | ~new_n11859_ | (new_n12030_ & new_n12006_)) & (~new_n11942_ | ~new_n11976_ | new_n11859_);
  assign new_n11942_ = new_n11943_ & new_n11975_;
  assign new_n11943_ = new_n11972_ & new_n11944_ & new_n11965_;
  assign new_n11944_ = ~new_n11945_ & (\all_features[4787]  | \all_features[4788]  | \all_features[4789]  | \all_features[4790]  | \all_features[4791] );
  assign new_n11945_ = ~new_n11961_ & (new_n11959_ | (~new_n11963_ & (new_n11964_ | (~new_n11962_ & ~new_n11946_))));
  assign new_n11946_ = ~new_n11947_ & (new_n11949_ | (new_n11958_ & (~new_n11953_ | (~new_n11957_ & new_n11956_))));
  assign new_n11947_ = ~new_n11948_ & ~\all_features[4791] ;
  assign new_n11948_ = \all_features[4789]  & \all_features[4790]  & (\all_features[4788]  | (\all_features[4786]  & \all_features[4787]  & \all_features[4785] ));
  assign new_n11949_ = ~\all_features[4791]  & (~\all_features[4790]  | ~new_n11950_ | ~new_n11951_ | ~new_n11952_);
  assign new_n11950_ = \all_features[4786]  & \all_features[4787] ;
  assign new_n11951_ = \all_features[4784]  & \all_features[4785] ;
  assign new_n11952_ = \all_features[4788]  & \all_features[4789] ;
  assign new_n11953_ = \all_features[4791]  & (\all_features[4790]  | (\all_features[4789]  & (\all_features[4788]  | ~new_n11955_ | ~new_n11954_)));
  assign new_n11954_ = ~\all_features[4784]  & ~\all_features[4785] ;
  assign new_n11955_ = ~\all_features[4786]  & ~\all_features[4787] ;
  assign new_n11956_ = \all_features[4791]  & (\all_features[4790]  | (new_n11952_ & (\all_features[4786]  | \all_features[4787]  | \all_features[4785] )));
  assign new_n11957_ = ~\all_features[4789]  & \all_features[4790]  & \all_features[4791]  & (\all_features[4788]  ? new_n11955_ : (new_n11951_ | ~new_n11955_));
  assign new_n11958_ = \all_features[4791]  & (\all_features[4789]  | \all_features[4790]  | \all_features[4788] );
  assign new_n11959_ = new_n11960_ & (~\all_features[4789]  | (~\all_features[4788]  & (~\all_features[4787]  | (~\all_features[4786]  & ~\all_features[4785] ))));
  assign new_n11960_ = ~\all_features[4790]  & ~\all_features[4791] ;
  assign new_n11961_ = ~\all_features[4789]  & new_n11960_ & ((~\all_features[4786]  & new_n11954_) | ~\all_features[4788]  | ~\all_features[4787] );
  assign new_n11962_ = ~\all_features[4791]  & (~\all_features[4790]  | (~\all_features[4789]  & (new_n11954_ | ~new_n11950_ | ~\all_features[4788] )));
  assign new_n11963_ = new_n11960_ & (~\all_features[4787]  | ~new_n11952_ | (~\all_features[4786]  & ~new_n11951_));
  assign new_n11964_ = ~\all_features[4791]  & (~\all_features[4790]  | (~\all_features[4788]  & ~\all_features[4789]  & ~new_n11950_));
  assign new_n11965_ = new_n11970_ & (~new_n11971_ | (~new_n11966_ & ~new_n11962_ & ~new_n11964_));
  assign new_n11966_ = ~new_n11947_ & ~new_n11949_ & (~new_n11958_ | ~new_n11953_ | new_n11967_);
  assign new_n11967_ = new_n11956_ & new_n11968_ & (new_n11969_ | ~\all_features[4789]  | ~\all_features[4790]  | ~\all_features[4791] );
  assign new_n11968_ = \all_features[4790]  & \all_features[4791]  & (\all_features[4788]  | \all_features[4789]  | new_n11951_ | ~new_n11955_);
  assign new_n11969_ = ~\all_features[4787]  & ~\all_features[4788]  & (~\all_features[4786]  | new_n11954_);
  assign new_n11970_ = ~new_n11961_ & (\all_features[4787]  | \all_features[4788]  | \all_features[4789]  | \all_features[4790]  | \all_features[4791] );
  assign new_n11971_ = ~new_n11959_ & ~new_n11963_;
  assign new_n11972_ = new_n11970_ & new_n11971_ & (new_n11974_ | new_n11947_ | new_n11962_ | ~new_n11973_);
  assign new_n11973_ = ~new_n11949_ & ~new_n11964_;
  assign new_n11974_ = new_n11958_ & new_n11968_ & new_n11953_ & new_n11956_;
  assign new_n11975_ = new_n11973_ & new_n11970_ & ~new_n11963_ & ~new_n11962_ & ~new_n11947_ & ~new_n11959_;
  assign new_n11976_ = ~new_n12002_ & new_n11977_;
  assign new_n11977_ = ~new_n11978_ & ~new_n12001_;
  assign new_n11978_ = new_n11989_ & (~new_n11979_ | (new_n11999_ & new_n12000_ & new_n11996_ & new_n11997_));
  assign new_n11979_ = ~new_n11988_ & ~new_n11986_ & ~new_n11980_ & ~new_n11983_;
  assign new_n11980_ = ~\all_features[3463]  & (~\all_features[3462]  | new_n11981_);
  assign new_n11981_ = ~\all_features[3461]  & (new_n11982_ | ~\all_features[3459]  | ~\all_features[3460]  | ~\all_features[3458] );
  assign new_n11982_ = ~\all_features[3456]  & ~\all_features[3457] ;
  assign new_n11983_ = ~\all_features[3463]  & (~new_n11985_ | ~\all_features[3458]  | ~\all_features[3459]  | ~\all_features[3462]  | ~new_n11984_);
  assign new_n11984_ = \all_features[3456]  & \all_features[3457] ;
  assign new_n11985_ = \all_features[3460]  & \all_features[3461] ;
  assign new_n11986_ = ~new_n11987_ & ~\all_features[3463] ;
  assign new_n11987_ = \all_features[3461]  & \all_features[3462]  & (\all_features[3460]  | (\all_features[3458]  & \all_features[3459]  & \all_features[3457] ));
  assign new_n11988_ = ~\all_features[3463]  & (~\all_features[3462]  | (~\all_features[3461]  & ~\all_features[3460]  & (~\all_features[3459]  | ~\all_features[3458] )));
  assign new_n11989_ = new_n11990_ & new_n11994_;
  assign new_n11990_ = ~new_n11991_ & ~new_n11993_;
  assign new_n11991_ = new_n11992_ & (~\all_features[3459]  | ~new_n11985_ | (~\all_features[3458]  & ~new_n11984_));
  assign new_n11992_ = ~\all_features[3462]  & ~\all_features[3463] ;
  assign new_n11993_ = new_n11992_ & (~\all_features[3461]  | (~\all_features[3460]  & (~\all_features[3459]  | (~\all_features[3458]  & ~\all_features[3457] ))));
  assign new_n11994_ = ~new_n11995_ & (\all_features[3459]  | \all_features[3460]  | \all_features[3461]  | \all_features[3462]  | \all_features[3463] );
  assign new_n11995_ = ~\all_features[3461]  & new_n11992_ & ((~\all_features[3458]  & new_n11982_) | ~\all_features[3460]  | ~\all_features[3459] );
  assign new_n11996_ = \all_features[3463]  & (\all_features[3462]  | (new_n11985_ & (\all_features[3458]  | \all_features[3459]  | \all_features[3457] )));
  assign new_n11997_ = \all_features[3462]  & \all_features[3463]  & (\all_features[3460]  | \all_features[3461]  | new_n11984_ | ~new_n11998_);
  assign new_n11998_ = ~\all_features[3458]  & ~\all_features[3459] ;
  assign new_n11999_ = \all_features[3463]  & (\all_features[3462]  | (\all_features[3461]  & (\all_features[3460]  | ~new_n11998_ | ~new_n11982_)));
  assign new_n12000_ = \all_features[3463]  & (\all_features[3461]  | \all_features[3462]  | \all_features[3460] );
  assign new_n12001_ = new_n11979_ & new_n11989_;
  assign new_n12002_ = new_n11994_ & (~new_n11990_ | (~new_n12003_ & ~new_n11980_ & ~new_n11988_));
  assign new_n12003_ = ~new_n11986_ & ~new_n11983_ & (~new_n12000_ | ~new_n11999_ | new_n12004_);
  assign new_n12004_ = new_n11996_ & new_n11997_ & (new_n12005_ | ~\all_features[3461]  | ~\all_features[3462]  | ~\all_features[3463] );
  assign new_n12005_ = ~\all_features[3459]  & ~\all_features[3460]  & (~\all_features[3458]  | new_n11982_);
  assign new_n12006_ = new_n12007_ & new_n12029_;
  assign new_n12007_ = new_n12008_ & (~new_n12017_ | (new_n12027_ & new_n12028_ & new_n12024_ & new_n12026_));
  assign new_n12008_ = new_n12009_ & ~new_n12013_ & ~new_n12014_;
  assign new_n12009_ = ~new_n12010_ & (\all_features[3667]  | \all_features[3668]  | \all_features[3669]  | \all_features[3670]  | \all_features[3671] );
  assign new_n12010_ = ~\all_features[3669]  & new_n12012_ & ((~\all_features[3666]  & new_n12011_) | ~\all_features[3668]  | ~\all_features[3667] );
  assign new_n12011_ = ~\all_features[3664]  & ~\all_features[3665] ;
  assign new_n12012_ = ~\all_features[3670]  & ~\all_features[3671] ;
  assign new_n12013_ = new_n12012_ & (~\all_features[3669]  | (~\all_features[3668]  & (~\all_features[3667]  | (~\all_features[3666]  & ~\all_features[3665] ))));
  assign new_n12014_ = new_n12012_ & (~\all_features[3667]  | ~new_n12015_ | (~\all_features[3666]  & ~new_n12016_));
  assign new_n12015_ = \all_features[3668]  & \all_features[3669] ;
  assign new_n12016_ = \all_features[3664]  & \all_features[3665] ;
  assign new_n12017_ = ~new_n12023_ & ~new_n12022_ & ~new_n12018_ & ~new_n12020_;
  assign new_n12018_ = ~\all_features[3671]  & (~\all_features[3670]  | (~\all_features[3669]  & (new_n12011_ | ~new_n12019_ | ~\all_features[3668] )));
  assign new_n12019_ = \all_features[3666]  & \all_features[3667] ;
  assign new_n12020_ = ~new_n12021_ & ~\all_features[3671] ;
  assign new_n12021_ = \all_features[3669]  & \all_features[3670]  & (\all_features[3668]  | (\all_features[3666]  & \all_features[3667]  & \all_features[3665] ));
  assign new_n12022_ = ~\all_features[3671]  & (~\all_features[3670]  | ~new_n12015_ | ~new_n12016_ | ~new_n12019_);
  assign new_n12023_ = ~\all_features[3671]  & (~\all_features[3670]  | (~\all_features[3668]  & ~\all_features[3669]  & ~new_n12019_));
  assign new_n12024_ = \all_features[3671]  & (\all_features[3670]  | (\all_features[3669]  & (\all_features[3668]  | ~new_n12011_ | ~new_n12025_)));
  assign new_n12025_ = ~\all_features[3666]  & ~\all_features[3667] ;
  assign new_n12026_ = \all_features[3671]  & (\all_features[3670]  | (new_n12015_ & (\all_features[3666]  | \all_features[3667]  | \all_features[3665] )));
  assign new_n12027_ = \all_features[3670]  & \all_features[3671]  & (\all_features[3668]  | \all_features[3669]  | new_n12016_ | ~new_n12025_);
  assign new_n12028_ = \all_features[3671]  & (\all_features[3669]  | \all_features[3670]  | \all_features[3668] );
  assign new_n12029_ = new_n12008_ & new_n12017_;
  assign new_n12030_ = new_n12031_ & new_n12035_;
  assign new_n12031_ = new_n12009_ & (new_n12014_ | new_n12013_ | (~new_n12018_ & ~new_n12023_ & ~new_n12032_));
  assign new_n12032_ = ~new_n12022_ & ~new_n12020_ & (~new_n12028_ | ~new_n12024_ | new_n12033_);
  assign new_n12033_ = new_n12026_ & new_n12027_ & (new_n12034_ | ~\all_features[3669]  | ~\all_features[3670]  | ~\all_features[3671] );
  assign new_n12034_ = ~\all_features[3667]  & ~\all_features[3668]  & (~\all_features[3666]  | new_n12011_);
  assign new_n12035_ = ~new_n12036_ & (\all_features[3667]  | \all_features[3668]  | \all_features[3669]  | \all_features[3670]  | \all_features[3671] );
  assign new_n12036_ = ~new_n12010_ & (new_n12013_ | (~new_n12014_ & (new_n12023_ | (~new_n12018_ & ~new_n12037_))));
  assign new_n12037_ = ~new_n12020_ & (new_n12022_ | (new_n12028_ & (~new_n12024_ | (~new_n12038_ & new_n12026_))));
  assign new_n12038_ = ~\all_features[3669]  & \all_features[3670]  & \all_features[3671]  & (\all_features[3668]  ? new_n12025_ : (new_n12016_ | ~new_n12025_));
  assign new_n12039_ = ~new_n12040_ & new_n12041_;
  assign new_n12040_ = new_n11901_ & ((~new_n11725_ & ~new_n11895_ & new_n11859_) | (~new_n11859_ & (~new_n11976_ | ~new_n11942_)));
  assign new_n12041_ = new_n11901_ | (new_n11897_ ? new_n12042_ : (new_n11902_ ? ~new_n11905_ : new_n11907_));
  assign new_n12042_ = new_n11756_ ? new_n11824_ : new_n11792_;
  assign new_n12043_ = ~new_n12258_ & new_n12044_;
  assign new_n12044_ = ~new_n12189_ & new_n12045_;
  assign new_n12045_ = new_n7949_ | (new_n8327_ ? (new_n12151_ ? ~new_n12188_ : new_n12153_) : new_n12046_);
  assign new_n12046_ = new_n12047_ ? new_n12082_ : ~new_n12117_;
  assign new_n12047_ = ~new_n12048_ & ~new_n12081_;
  assign new_n12048_ = new_n12049_ & new_n12077_;
  assign new_n12049_ = new_n12050_ & new_n12074_;
  assign new_n12050_ = new_n12066_ & (~new_n12069_ | (~new_n12051_ & ~new_n12072_ & ~new_n12073_));
  assign new_n12051_ = ~new_n12060_ & ~new_n12062_ & (~new_n12065_ | ~new_n12064_ | new_n12052_);
  assign new_n12052_ = new_n12053_ & new_n12055_ & (new_n12058_ | ~\all_features[3229]  | ~\all_features[3230]  | ~\all_features[3231] );
  assign new_n12053_ = \all_features[3231]  & (\all_features[3230]  | (new_n12054_ & (\all_features[3226]  | \all_features[3227]  | \all_features[3225] )));
  assign new_n12054_ = \all_features[3228]  & \all_features[3229] ;
  assign new_n12055_ = \all_features[3230]  & \all_features[3231]  & (\all_features[3228]  | \all_features[3229]  | new_n12056_ | ~new_n12057_);
  assign new_n12056_ = \all_features[3224]  & \all_features[3225] ;
  assign new_n12057_ = ~\all_features[3226]  & ~\all_features[3227] ;
  assign new_n12058_ = ~\all_features[3227]  & ~\all_features[3228]  & (~\all_features[3226]  | new_n12059_);
  assign new_n12059_ = ~\all_features[3224]  & ~\all_features[3225] ;
  assign new_n12060_ = ~new_n12061_ & ~\all_features[3231] ;
  assign new_n12061_ = \all_features[3229]  & \all_features[3230]  & (\all_features[3228]  | (\all_features[3226]  & \all_features[3227]  & \all_features[3225] ));
  assign new_n12062_ = ~\all_features[3231]  & (~\all_features[3230]  | ~new_n12063_ | ~new_n12056_ | ~new_n12054_);
  assign new_n12063_ = \all_features[3226]  & \all_features[3227] ;
  assign new_n12064_ = \all_features[3231]  & (\all_features[3230]  | (\all_features[3229]  & (\all_features[3228]  | ~new_n12057_ | ~new_n12059_)));
  assign new_n12065_ = \all_features[3231]  & (\all_features[3229]  | \all_features[3230]  | \all_features[3228] );
  assign new_n12066_ = ~new_n12067_ & (\all_features[3227]  | \all_features[3228]  | \all_features[3229]  | \all_features[3230]  | \all_features[3231] );
  assign new_n12067_ = ~\all_features[3229]  & new_n12068_ & ((~\all_features[3226]  & new_n12059_) | ~\all_features[3228]  | ~\all_features[3227] );
  assign new_n12068_ = ~\all_features[3230]  & ~\all_features[3231] ;
  assign new_n12069_ = ~new_n12070_ & ~new_n12071_;
  assign new_n12070_ = new_n12068_ & (~\all_features[3229]  | (~\all_features[3228]  & (~\all_features[3227]  | (~\all_features[3226]  & ~\all_features[3225] ))));
  assign new_n12071_ = new_n12068_ & (~\all_features[3227]  | ~new_n12054_ | (~\all_features[3226]  & ~new_n12056_));
  assign new_n12072_ = ~\all_features[3231]  & (~\all_features[3230]  | (~\all_features[3229]  & (new_n12059_ | ~new_n12063_ | ~\all_features[3228] )));
  assign new_n12073_ = ~\all_features[3231]  & (~\all_features[3230]  | (~\all_features[3228]  & ~\all_features[3229]  & ~new_n12063_));
  assign new_n12074_ = new_n12066_ & new_n12069_ & (new_n12076_ | new_n12060_ | new_n12072_ | ~new_n12075_);
  assign new_n12075_ = ~new_n12062_ & ~new_n12073_;
  assign new_n12076_ = new_n12065_ & new_n12055_ & new_n12064_ & new_n12053_;
  assign new_n12077_ = ~new_n12078_ & (\all_features[3227]  | \all_features[3228]  | \all_features[3229]  | \all_features[3230]  | \all_features[3231] );
  assign new_n12078_ = ~new_n12067_ & (new_n12070_ | (~new_n12071_ & (new_n12073_ | (~new_n12072_ & ~new_n12079_))));
  assign new_n12079_ = ~new_n12060_ & (new_n12062_ | (new_n12065_ & (~new_n12064_ | (~new_n12080_ & new_n12053_))));
  assign new_n12080_ = ~\all_features[3229]  & \all_features[3230]  & \all_features[3231]  & (\all_features[3228]  ? new_n12057_ : (new_n12056_ | ~new_n12057_));
  assign new_n12081_ = new_n12075_ & new_n12066_ & ~new_n12071_ & ~new_n12072_ & ~new_n12060_ & ~new_n12070_;
  assign new_n12082_ = new_n12083_ & ~new_n12112_ & ~new_n12115_;
  assign new_n12083_ = ~new_n12084_ & ~new_n12108_;
  assign new_n12084_ = new_n12099_ & (~new_n12104_ | (~new_n12102_ & ~new_n12085_ & ~new_n12107_));
  assign new_n12085_ = ~new_n12097_ & ~new_n12095_ & (~new_n12098_ | ~new_n12094_ | new_n12086_);
  assign new_n12086_ = new_n12087_ & new_n12089_ & (new_n12092_ | ~\all_features[4141]  | ~\all_features[4142]  | ~\all_features[4143] );
  assign new_n12087_ = \all_features[4143]  & (\all_features[4142]  | (new_n12088_ & (\all_features[4138]  | \all_features[4139]  | \all_features[4137] )));
  assign new_n12088_ = \all_features[4140]  & \all_features[4141] ;
  assign new_n12089_ = \all_features[4142]  & \all_features[4143]  & (\all_features[4140]  | \all_features[4141]  | new_n12091_ | ~new_n12090_);
  assign new_n12090_ = ~\all_features[4138]  & ~\all_features[4139] ;
  assign new_n12091_ = \all_features[4136]  & \all_features[4137] ;
  assign new_n12092_ = ~\all_features[4139]  & ~\all_features[4140]  & (~\all_features[4138]  | new_n12093_);
  assign new_n12093_ = ~\all_features[4136]  & ~\all_features[4137] ;
  assign new_n12094_ = \all_features[4143]  & (\all_features[4142]  | (\all_features[4141]  & (\all_features[4140]  | ~new_n12090_ | ~new_n12093_)));
  assign new_n12095_ = ~new_n12096_ & ~\all_features[4143] ;
  assign new_n12096_ = \all_features[4141]  & \all_features[4142]  & (\all_features[4140]  | (\all_features[4138]  & \all_features[4139]  & \all_features[4137] ));
  assign new_n12097_ = ~\all_features[4143]  & (~new_n12091_ | ~\all_features[4138]  | ~\all_features[4139]  | ~\all_features[4142]  | ~new_n12088_);
  assign new_n12098_ = \all_features[4143]  & (\all_features[4141]  | \all_features[4142]  | \all_features[4140] );
  assign new_n12099_ = ~new_n12100_ & (\all_features[4139]  | \all_features[4140]  | \all_features[4141]  | \all_features[4142]  | \all_features[4143] );
  assign new_n12100_ = ~\all_features[4141]  & new_n12101_ & ((~\all_features[4138]  & new_n12093_) | ~\all_features[4140]  | ~\all_features[4139] );
  assign new_n12101_ = ~\all_features[4142]  & ~\all_features[4143] ;
  assign new_n12102_ = ~\all_features[4143]  & (~\all_features[4142]  | new_n12103_);
  assign new_n12103_ = ~\all_features[4141]  & (new_n12093_ | ~\all_features[4139]  | ~\all_features[4140]  | ~\all_features[4138] );
  assign new_n12104_ = ~new_n12105_ & ~new_n12106_;
  assign new_n12105_ = new_n12101_ & (~\all_features[4139]  | ~new_n12088_ | (~new_n12091_ & ~\all_features[4138] ));
  assign new_n12106_ = new_n12101_ & (~\all_features[4141]  | (~\all_features[4140]  & (~\all_features[4139]  | (~\all_features[4138]  & ~\all_features[4137] ))));
  assign new_n12107_ = ~\all_features[4143]  & (~\all_features[4142]  | (~\all_features[4141]  & ~\all_features[4140]  & (~\all_features[4139]  | ~\all_features[4138] )));
  assign new_n12108_ = ~new_n12109_ & (\all_features[4139]  | \all_features[4140]  | \all_features[4141]  | \all_features[4142]  | \all_features[4143] );
  assign new_n12109_ = ~new_n12100_ & (new_n12106_ | (~new_n12105_ & (new_n12107_ | (~new_n12102_ & ~new_n12110_))));
  assign new_n12110_ = ~new_n12095_ & (new_n12097_ | (new_n12098_ & (~new_n12094_ | (~new_n12111_ & new_n12087_))));
  assign new_n12111_ = ~\all_features[4141]  & \all_features[4142]  & \all_features[4143]  & (\all_features[4140]  ? new_n12090_ : (new_n12091_ | ~new_n12090_));
  assign new_n12112_ = new_n12104_ & ~new_n12113_ & new_n12099_;
  assign new_n12113_ = ~new_n12107_ & ~new_n12097_ & ~new_n12095_ & ~new_n12102_ & ~new_n12114_;
  assign new_n12114_ = new_n12098_ & new_n12094_ & new_n12087_ & new_n12089_;
  assign new_n12115_ = new_n12099_ & new_n12116_ & ~new_n12095_ & ~new_n12106_;
  assign new_n12116_ = ~new_n12107_ & ~new_n12105_ & ~new_n12102_ & ~new_n12097_;
  assign new_n12117_ = new_n12118_ & new_n12142_;
  assign new_n12118_ = ~new_n12119_ & ~new_n12141_;
  assign new_n12119_ = new_n12120_ & (~new_n12129_ | (new_n12139_ & new_n12140_ & new_n12136_ & new_n12138_));
  assign new_n12120_ = new_n12121_ & ~new_n12125_ & ~new_n12126_;
  assign new_n12121_ = ~new_n12122_ & (\all_features[3283]  | \all_features[3284]  | \all_features[3285]  | \all_features[3286]  | \all_features[3287] );
  assign new_n12122_ = ~\all_features[3285]  & new_n12124_ & ((~\all_features[3282]  & new_n12123_) | ~\all_features[3284]  | ~\all_features[3283] );
  assign new_n12123_ = ~\all_features[3280]  & ~\all_features[3281] ;
  assign new_n12124_ = ~\all_features[3286]  & ~\all_features[3287] ;
  assign new_n12125_ = new_n12124_ & (~\all_features[3285]  | (~\all_features[3284]  & (~\all_features[3283]  | (~\all_features[3282]  & ~\all_features[3281] ))));
  assign new_n12126_ = new_n12124_ & (~\all_features[3283]  | ~new_n12127_ | (~\all_features[3282]  & ~new_n12128_));
  assign new_n12127_ = \all_features[3284]  & \all_features[3285] ;
  assign new_n12128_ = \all_features[3280]  & \all_features[3281] ;
  assign new_n12129_ = ~new_n12135_ & ~new_n12134_ & ~new_n12130_ & ~new_n12132_;
  assign new_n12130_ = ~\all_features[3287]  & (~\all_features[3286]  | (~\all_features[3285]  & (new_n12123_ | ~new_n12131_ | ~\all_features[3284] )));
  assign new_n12131_ = \all_features[3282]  & \all_features[3283] ;
  assign new_n12132_ = ~new_n12133_ & ~\all_features[3287] ;
  assign new_n12133_ = \all_features[3285]  & \all_features[3286]  & (\all_features[3284]  | (\all_features[3282]  & \all_features[3283]  & \all_features[3281] ));
  assign new_n12134_ = ~\all_features[3287]  & (~\all_features[3286]  | ~new_n12127_ | ~new_n12128_ | ~new_n12131_);
  assign new_n12135_ = ~\all_features[3287]  & (~\all_features[3286]  | (~\all_features[3284]  & ~\all_features[3285]  & ~new_n12131_));
  assign new_n12136_ = \all_features[3287]  & (\all_features[3286]  | (\all_features[3285]  & (\all_features[3284]  | ~new_n12123_ | ~new_n12137_)));
  assign new_n12137_ = ~\all_features[3282]  & ~\all_features[3283] ;
  assign new_n12138_ = \all_features[3287]  & (\all_features[3286]  | (new_n12127_ & (\all_features[3282]  | \all_features[3283]  | \all_features[3281] )));
  assign new_n12139_ = \all_features[3286]  & \all_features[3287]  & (\all_features[3284]  | \all_features[3285]  | new_n12128_ | ~new_n12137_);
  assign new_n12140_ = \all_features[3287]  & (\all_features[3285]  | \all_features[3286]  | \all_features[3284] );
  assign new_n12141_ = new_n12120_ & new_n12129_;
  assign new_n12142_ = ~new_n12143_ & ~new_n12147_;
  assign new_n12143_ = ~new_n12144_ & (\all_features[3283]  | \all_features[3284]  | \all_features[3285]  | \all_features[3286]  | \all_features[3287] );
  assign new_n12144_ = ~new_n12122_ & (new_n12125_ | (~new_n12126_ & (new_n12135_ | (~new_n12130_ & ~new_n12145_))));
  assign new_n12145_ = ~new_n12132_ & (new_n12134_ | (new_n12140_ & (~new_n12136_ | (~new_n12146_ & new_n12138_))));
  assign new_n12146_ = ~\all_features[3285]  & \all_features[3286]  & \all_features[3287]  & (\all_features[3284]  ? new_n12137_ : (new_n12128_ | ~new_n12137_));
  assign new_n12147_ = new_n12121_ & (new_n12126_ | new_n12125_ | (~new_n12130_ & ~new_n12135_ & ~new_n12148_));
  assign new_n12148_ = ~new_n12134_ & ~new_n12132_ & (~new_n12140_ | ~new_n12136_ | new_n12149_);
  assign new_n12149_ = new_n12138_ & new_n12139_ & (new_n12150_ | ~\all_features[3285]  | ~\all_features[3286]  | ~\all_features[3287] );
  assign new_n12150_ = ~\all_features[3283]  & ~\all_features[3284]  & (~\all_features[3282]  | new_n12123_);
  assign new_n12151_ = ~new_n10574_ & new_n12152_;
  assign new_n12152_ = ~new_n10604_ & ~new_n10607_;
  assign new_n12153_ = ~new_n12154_ & new_n12184_;
  assign new_n12154_ = new_n12155_ & new_n12175_;
  assign new_n12155_ = ~new_n12174_ & (new_n12169_ | (~new_n12171_ & (new_n12172_ | (~new_n12156_ & ~new_n12173_))));
  assign new_n12156_ = ~new_n12163_ & (new_n12166_ | (~new_n12165_ & (~new_n12168_ | new_n12157_)));
  assign new_n12157_ = \all_features[3503]  & ((~new_n12162_ & ~\all_features[3501]  & \all_features[3502] ) | (~new_n12160_ & (\all_features[3502]  | (~new_n12158_ & \all_features[3501] ))));
  assign new_n12158_ = new_n12159_ & ~\all_features[3500]  & ~\all_features[3498]  & ~\all_features[3499] ;
  assign new_n12159_ = ~\all_features[3496]  & ~\all_features[3497] ;
  assign new_n12160_ = \all_features[3503]  & (\all_features[3502]  | (new_n12161_ & (\all_features[3498]  | \all_features[3499]  | \all_features[3497] )));
  assign new_n12161_ = \all_features[3500]  & \all_features[3501] ;
  assign new_n12162_ = (~\all_features[3498]  & ~\all_features[3499]  & ~\all_features[3500]  & (~\all_features[3497]  | ~\all_features[3496] )) | (\all_features[3500]  & (\all_features[3498]  | \all_features[3499] ));
  assign new_n12163_ = ~\all_features[3503]  & (~\all_features[3502]  | (~\all_features[3501]  & (new_n12159_ | ~new_n12164_ | ~\all_features[3500] )));
  assign new_n12164_ = \all_features[3498]  & \all_features[3499] ;
  assign new_n12165_ = ~\all_features[3503]  & (~new_n12164_ | ~\all_features[3496]  | ~\all_features[3497]  | ~\all_features[3502]  | ~new_n12161_);
  assign new_n12166_ = ~new_n12167_ & ~\all_features[3503] ;
  assign new_n12167_ = \all_features[3501]  & \all_features[3502]  & (\all_features[3500]  | (\all_features[3498]  & \all_features[3499]  & \all_features[3497] ));
  assign new_n12168_ = \all_features[3503]  & (\all_features[3501]  | \all_features[3502]  | \all_features[3500] );
  assign new_n12169_ = ~\all_features[3501]  & new_n12170_ & ((~\all_features[3498]  & new_n12159_) | ~\all_features[3500]  | ~\all_features[3499] );
  assign new_n12170_ = ~\all_features[3502]  & ~\all_features[3503] ;
  assign new_n12171_ = new_n12170_ & (~\all_features[3501]  | (~\all_features[3500]  & (~\all_features[3499]  | (~\all_features[3498]  & ~\all_features[3497] ))));
  assign new_n12172_ = new_n12170_ & (~new_n12161_ | ~\all_features[3499]  | (~\all_features[3498]  & (~\all_features[3496]  | ~\all_features[3497] )));
  assign new_n12173_ = ~\all_features[3503]  & (~\all_features[3502]  | (~\all_features[3500]  & ~\all_features[3501]  & ~new_n12164_));
  assign new_n12174_ = ~\all_features[3503]  & ~\all_features[3502]  & ~\all_features[3501]  & ~\all_features[3499]  & ~\all_features[3500] ;
  assign new_n12175_ = new_n12181_ & (~new_n12183_ | (~new_n12173_ & ~new_n12163_ & (~new_n12182_ | new_n12176_)));
  assign new_n12176_ = new_n12177_ & (~new_n12178_ | (~new_n12180_ & \all_features[3501]  & \all_features[3502]  & \all_features[3503] ));
  assign new_n12177_ = \all_features[3503]  & (\all_features[3502]  | (~new_n12158_ & \all_features[3501] ));
  assign new_n12178_ = \all_features[3503]  & \all_features[3502]  & ~new_n12179_ & new_n12160_;
  assign new_n12179_ = ~\all_features[3498]  & ~\all_features[3499]  & ~\all_features[3500]  & ~\all_features[3501]  & (~\all_features[3497]  | ~\all_features[3496] );
  assign new_n12180_ = ~\all_features[3499]  & ~\all_features[3500]  & (~\all_features[3498]  | new_n12159_);
  assign new_n12181_ = ~new_n12169_ & ~new_n12174_;
  assign new_n12182_ = ~new_n12165_ & ~new_n12166_;
  assign new_n12183_ = ~new_n12171_ & ~new_n12172_;
  assign new_n12184_ = ~new_n12185_ & ~new_n12187_;
  assign new_n12185_ = new_n12183_ & ~new_n12186_ & new_n12181_;
  assign new_n12186_ = ~new_n12173_ & ~new_n12163_ & ~new_n12165_ & ~new_n12166_ & (~new_n12178_ | ~new_n12177_);
  assign new_n12187_ = new_n12182_ & new_n12181_ & ~new_n12163_ & ~new_n12173_ & ~new_n12171_ & ~new_n12172_;
  assign new_n12188_ = ~new_n9455_ & (~new_n9445_ | ~new_n9452_ | ~new_n9424_);
  assign new_n12189_ = new_n7949_ & (new_n7407_ ? (new_n12228_ ? new_n12196_ : ~new_n12227_) : ~new_n12190_);
  assign new_n12190_ = new_n8201_ & new_n12191_;
  assign new_n12191_ = ~new_n8227_ & ~new_n12192_;
  assign new_n12192_ = ~new_n12193_ & (\all_features[3027]  | \all_features[3028]  | \all_features[3029]  | \all_features[3030]  | \all_features[3031] );
  assign new_n12193_ = ~new_n8220_ & (new_n8223_ | (~new_n8224_ & (new_n8218_ | (~new_n8204_ & ~new_n12194_))));
  assign new_n12194_ = ~new_n8215_ & (new_n8217_ | (new_n8214_ & (~new_n8213_ | (~new_n12195_ & new_n8208_))));
  assign new_n12195_ = ~\all_features[3029]  & \all_features[3030]  & \all_features[3031]  & (\all_features[3028]  ? new_n8211_ : (new_n8212_ | ~new_n8211_));
  assign new_n12196_ = ~new_n12197_ & ~new_n12226_;
  assign new_n12197_ = new_n12198_ & new_n12220_;
  assign new_n12198_ = new_n12215_ & ~new_n12219_ & ~new_n12199_ & ~new_n12218_;
  assign new_n12199_ = new_n12200_ & ~new_n12213_ & (~new_n12208_ | ~new_n12214_ | ~new_n12211_ | ~new_n12212_);
  assign new_n12200_ = ~new_n12205_ & ~new_n12201_ & ~new_n12203_;
  assign new_n12201_ = ~new_n12202_ & ~\all_features[5263] ;
  assign new_n12202_ = \all_features[5261]  & \all_features[5262]  & (\all_features[5260]  | (\all_features[5258]  & \all_features[5259]  & \all_features[5257] ));
  assign new_n12203_ = ~\all_features[5263]  & (~\all_features[5262]  | (~\all_features[5260]  & ~\all_features[5261]  & ~new_n12204_));
  assign new_n12204_ = \all_features[5258]  & \all_features[5259] ;
  assign new_n12205_ = ~\all_features[5263]  & (~\all_features[5262]  | ~new_n12206_ | ~new_n12207_ | ~new_n12204_);
  assign new_n12206_ = \all_features[5260]  & \all_features[5261] ;
  assign new_n12207_ = \all_features[5256]  & \all_features[5257] ;
  assign new_n12208_ = \all_features[5263]  & (\all_features[5262]  | (\all_features[5261]  & (\all_features[5260]  | ~new_n12210_ | ~new_n12209_)));
  assign new_n12209_ = ~\all_features[5258]  & ~\all_features[5259] ;
  assign new_n12210_ = ~\all_features[5256]  & ~\all_features[5257] ;
  assign new_n12211_ = \all_features[5263]  & (\all_features[5262]  | (new_n12206_ & (\all_features[5258]  | \all_features[5259]  | \all_features[5257] )));
  assign new_n12212_ = \all_features[5262]  & \all_features[5263]  & (\all_features[5260]  | \all_features[5261]  | new_n12207_ | ~new_n12209_);
  assign new_n12213_ = ~\all_features[5263]  & (~\all_features[5262]  | (~\all_features[5261]  & (new_n12210_ | ~new_n12204_ | ~\all_features[5260] )));
  assign new_n12214_ = \all_features[5263]  & (\all_features[5261]  | \all_features[5262]  | \all_features[5260] );
  assign new_n12215_ = ~new_n12216_ & (\all_features[5259]  | \all_features[5260]  | \all_features[5261]  | \all_features[5262]  | \all_features[5263] );
  assign new_n12216_ = new_n12217_ & (~\all_features[5259]  | ~new_n12206_ | (~\all_features[5258]  & ~new_n12207_));
  assign new_n12217_ = ~\all_features[5262]  & ~\all_features[5263] ;
  assign new_n12218_ = new_n12217_ & (~\all_features[5261]  | (~\all_features[5260]  & (~\all_features[5259]  | (~\all_features[5258]  & ~\all_features[5257] ))));
  assign new_n12219_ = ~\all_features[5261]  & new_n12217_ & ((~\all_features[5258]  & new_n12210_) | ~\all_features[5260]  | ~\all_features[5259] );
  assign new_n12220_ = new_n12225_ & (~new_n12224_ | (~new_n12221_ & ~new_n12213_ & ~new_n12203_));
  assign new_n12221_ = ~new_n12205_ & ~new_n12201_ & (~new_n12214_ | ~new_n12208_ | new_n12222_);
  assign new_n12222_ = new_n12211_ & new_n12212_ & (new_n12223_ | ~\all_features[5261]  | ~\all_features[5262]  | ~\all_features[5263] );
  assign new_n12223_ = ~\all_features[5259]  & ~\all_features[5260]  & (~\all_features[5258]  | new_n12210_);
  assign new_n12224_ = ~new_n12218_ & ~new_n12216_;
  assign new_n12225_ = ~new_n12219_ & (\all_features[5259]  | \all_features[5260]  | \all_features[5261]  | \all_features[5262]  | \all_features[5263] );
  assign new_n12226_ = new_n12200_ & new_n12225_ & ~new_n12213_ & new_n12224_;
  assign new_n12227_ = new_n10774_ & new_n10775_;
  assign new_n12228_ = ~new_n12229_ & new_n12253_;
  assign new_n12229_ = new_n12250_ & (~new_n12244_ | (~new_n12230_ & ~new_n12248_ & ~new_n12252_));
  assign new_n12230_ = ~new_n12241_ & ~new_n12240_ & (~new_n12243_ | ~new_n12239_ | new_n12231_);
  assign new_n12231_ = new_n12232_ & new_n12234_ & (new_n12237_ | ~\all_features[3013]  | ~\all_features[3014]  | ~\all_features[3015] );
  assign new_n12232_ = \all_features[3015]  & (\all_features[3014]  | (new_n12233_ & (\all_features[3010]  | \all_features[3011]  | \all_features[3009] )));
  assign new_n12233_ = \all_features[3012]  & \all_features[3013] ;
  assign new_n12234_ = \all_features[3014]  & \all_features[3015]  & (\all_features[3012]  | \all_features[3013]  | new_n12235_ | ~new_n12236_);
  assign new_n12235_ = \all_features[3008]  & \all_features[3009] ;
  assign new_n12236_ = ~\all_features[3010]  & ~\all_features[3011] ;
  assign new_n12237_ = ~\all_features[3011]  & ~\all_features[3012]  & (~\all_features[3010]  | new_n12238_);
  assign new_n12238_ = ~\all_features[3008]  & ~\all_features[3009] ;
  assign new_n12239_ = \all_features[3015]  & (\all_features[3014]  | (\all_features[3013]  & (\all_features[3012]  | ~new_n12238_ | ~new_n12236_)));
  assign new_n12240_ = ~\all_features[3015]  & (~new_n12233_ | ~\all_features[3010]  | ~\all_features[3011]  | ~\all_features[3014]  | ~new_n12235_);
  assign new_n12241_ = ~new_n12242_ & ~\all_features[3015] ;
  assign new_n12242_ = \all_features[3013]  & \all_features[3014]  & (\all_features[3012]  | (\all_features[3010]  & \all_features[3011]  & \all_features[3009] ));
  assign new_n12243_ = \all_features[3015]  & (\all_features[3013]  | \all_features[3014]  | \all_features[3012] );
  assign new_n12244_ = ~new_n12245_ & ~new_n12247_;
  assign new_n12245_ = new_n12246_ & (~\all_features[3011]  | ~new_n12233_ | (~\all_features[3010]  & ~new_n12235_));
  assign new_n12246_ = ~\all_features[3014]  & ~\all_features[3015] ;
  assign new_n12247_ = new_n12246_ & (~\all_features[3013]  | (~\all_features[3012]  & (~\all_features[3011]  | (~\all_features[3010]  & ~\all_features[3009] ))));
  assign new_n12248_ = ~\all_features[3015]  & (~\all_features[3014]  | new_n12249_);
  assign new_n12249_ = ~\all_features[3013]  & (new_n12238_ | ~\all_features[3011]  | ~\all_features[3012]  | ~\all_features[3010] );
  assign new_n12250_ = ~new_n12251_ & (\all_features[3011]  | \all_features[3012]  | \all_features[3013]  | \all_features[3014]  | \all_features[3015] );
  assign new_n12251_ = ~\all_features[3013]  & new_n12246_ & ((~\all_features[3010]  & new_n12238_) | ~\all_features[3012]  | ~\all_features[3011] );
  assign new_n12252_ = ~\all_features[3015]  & (~\all_features[3014]  | (~\all_features[3013]  & ~\all_features[3012]  & (~\all_features[3011]  | ~\all_features[3010] )));
  assign new_n12253_ = ~new_n12254_ & ~new_n12257_;
  assign new_n12254_ = new_n12244_ & new_n12250_ & (new_n12248_ | new_n12255_ | new_n12240_ | ~new_n12256_);
  assign new_n12255_ = new_n12243_ & new_n12239_ & new_n12232_ & new_n12234_;
  assign new_n12256_ = ~new_n12241_ & ~new_n12252_;
  assign new_n12257_ = new_n12244_ & new_n12256_ & new_n12250_ & ~new_n12248_ & ~new_n12240_;
  assign new_n12258_ = new_n7949_ ? new_n12259_ : ((new_n12188_ | ~new_n12151_ | ~new_n8327_) & (~new_n12046_ | new_n8327_));
  assign new_n12259_ = new_n7407_ ? (new_n12228_ ? new_n12196_ : ~new_n12227_) : ~new_n12190_;
  assign new_n12260_ = ~new_n12261_ & new_n12449_;
  assign new_n12261_ = new_n12262_ & (~new_n12338_ | new_n12445_);
  assign new_n12262_ = new_n12263_ & (new_n12338_ | (new_n12371_ & (new_n12408_ ? new_n12374_ : new_n12443_)));
  assign new_n12263_ = ~new_n12338_ | ((new_n12267_ | ~new_n12264_) & (new_n12303_ | new_n12354_ | new_n12264_));
  assign new_n12264_ = ~new_n12265_ & new_n12266_;
  assign new_n12265_ = new_n11305_ & new_n11329_;
  assign new_n12266_ = ~new_n11333_ & ~new_n11335_;
  assign new_n12267_ = ~new_n12301_ & (~new_n12298_ | new_n12268_);
  assign new_n12268_ = ~new_n12269_ & ~new_n12294_;
  assign new_n12269_ = new_n12286_ & (~new_n12290_ | (~new_n12284_ & ~new_n12270_ & ~new_n12293_));
  assign new_n12270_ = ~new_n12279_ & ~new_n12281_ & (~new_n12283_ | ~new_n12282_ | new_n12271_);
  assign new_n12271_ = new_n12272_ & new_n12274_ & (new_n12277_ | ~\all_features[1189]  | ~\all_features[1190]  | ~\all_features[1191] );
  assign new_n12272_ = \all_features[1191]  & (\all_features[1190]  | (new_n12273_ & (\all_features[1186]  | \all_features[1187]  | \all_features[1185] )));
  assign new_n12273_ = \all_features[1188]  & \all_features[1189] ;
  assign new_n12274_ = \all_features[1190]  & \all_features[1191]  & (\all_features[1188]  | \all_features[1189]  | new_n12275_ | ~new_n12276_);
  assign new_n12275_ = \all_features[1184]  & \all_features[1185] ;
  assign new_n12276_ = ~\all_features[1186]  & ~\all_features[1187] ;
  assign new_n12277_ = ~\all_features[1187]  & ~\all_features[1188]  & (~\all_features[1186]  | new_n12278_);
  assign new_n12278_ = ~\all_features[1184]  & ~\all_features[1185] ;
  assign new_n12279_ = ~new_n12280_ & ~\all_features[1191] ;
  assign new_n12280_ = \all_features[1189]  & \all_features[1190]  & (\all_features[1188]  | (\all_features[1186]  & \all_features[1187]  & \all_features[1185] ));
  assign new_n12281_ = ~\all_features[1191]  & (~new_n12273_ | ~\all_features[1186]  | ~\all_features[1187]  | ~\all_features[1190]  | ~new_n12275_);
  assign new_n12282_ = \all_features[1191]  & (\all_features[1190]  | (\all_features[1189]  & (\all_features[1188]  | ~new_n12276_ | ~new_n12278_)));
  assign new_n12283_ = \all_features[1191]  & (\all_features[1189]  | \all_features[1190]  | \all_features[1188] );
  assign new_n12284_ = ~\all_features[1191]  & (~\all_features[1190]  | new_n12285_);
  assign new_n12285_ = ~\all_features[1189]  & (new_n12278_ | ~\all_features[1187]  | ~\all_features[1188]  | ~\all_features[1186] );
  assign new_n12286_ = ~new_n12287_ & ~new_n12289_;
  assign new_n12287_ = ~\all_features[1189]  & new_n12288_ & ((~\all_features[1186]  & new_n12278_) | ~\all_features[1188]  | ~\all_features[1187] );
  assign new_n12288_ = ~\all_features[1190]  & ~\all_features[1191] ;
  assign new_n12289_ = ~\all_features[1191]  & ~\all_features[1190]  & ~\all_features[1189]  & ~\all_features[1187]  & ~\all_features[1188] ;
  assign new_n12290_ = ~new_n12291_ & ~new_n12292_;
  assign new_n12291_ = new_n12288_ & (~\all_features[1189]  | (~\all_features[1188]  & (~\all_features[1187]  | (~\all_features[1186]  & ~\all_features[1185] ))));
  assign new_n12292_ = new_n12288_ & (~\all_features[1187]  | ~new_n12273_ | (~\all_features[1186]  & ~new_n12275_));
  assign new_n12293_ = ~\all_features[1191]  & (~\all_features[1190]  | (~\all_features[1189]  & ~\all_features[1188]  & (~\all_features[1187]  | ~\all_features[1186] )));
  assign new_n12294_ = ~new_n12295_ & ~new_n12289_;
  assign new_n12295_ = ~new_n12287_ & (new_n12291_ | (~new_n12292_ & (new_n12293_ | (~new_n12284_ & ~new_n12296_))));
  assign new_n12296_ = ~new_n12279_ & (new_n12281_ | (new_n12283_ & (~new_n12282_ | (~new_n12297_ & new_n12272_))));
  assign new_n12297_ = ~\all_features[1189]  & \all_features[1190]  & \all_features[1191]  & (\all_features[1188]  ? new_n12276_ : (new_n12275_ | ~new_n12276_));
  assign new_n12298_ = new_n12290_ & ~new_n12299_ & new_n12286_;
  assign new_n12299_ = ~new_n12293_ & ~new_n12281_ & ~new_n12279_ & ~new_n12284_ & ~new_n12300_;
  assign new_n12300_ = new_n12283_ & new_n12274_ & new_n12282_ & new_n12272_;
  assign new_n12301_ = new_n12302_ & ~new_n12293_ & ~new_n12287_ & ~new_n12284_ & ~new_n12292_;
  assign new_n12302_ = ~new_n12289_ & ~new_n12281_ & ~new_n12279_ & ~new_n12291_;
  assign new_n12303_ = ~new_n12337_ & (~new_n12334_ | new_n12304_);
  assign new_n12304_ = ~new_n12305_ & (new_n12324_ | (~new_n12330_ & ~new_n12322_));
  assign new_n12305_ = new_n12321_ & (~new_n12325_ | (~new_n12306_ & ~new_n12328_ & ~new_n12329_));
  assign new_n12306_ = ~new_n12318_ & ~new_n12316_ & (~new_n12320_ | new_n12310_ | ~new_n12307_);
  assign new_n12307_ = \all_features[1751]  & (\all_features[1750]  | new_n12308_);
  assign new_n12308_ = \all_features[1749]  & (\all_features[1746]  | \all_features[1747]  | \all_features[1748]  | ~new_n12309_);
  assign new_n12309_ = ~\all_features[1744]  & ~\all_features[1745] ;
  assign new_n12310_ = ~new_n12313_ & new_n12311_ & \all_features[1750]  & \all_features[1751]  & (~\all_features[1749]  | new_n12315_);
  assign new_n12311_ = \all_features[1751]  & (\all_features[1750]  | (new_n12312_ & (\all_features[1746]  | \all_features[1747]  | \all_features[1745] )));
  assign new_n12312_ = \all_features[1748]  & \all_features[1749] ;
  assign new_n12313_ = ~\all_features[1749]  & ~\all_features[1748]  & ~\all_features[1747]  & ~new_n12314_ & ~\all_features[1746] ;
  assign new_n12314_ = \all_features[1744]  & \all_features[1745] ;
  assign new_n12315_ = ~\all_features[1747]  & ~\all_features[1748]  & (~\all_features[1746]  | new_n12309_);
  assign new_n12316_ = ~new_n12317_ & ~\all_features[1751] ;
  assign new_n12317_ = \all_features[1749]  & \all_features[1750]  & (\all_features[1748]  | (\all_features[1746]  & \all_features[1747]  & \all_features[1745] ));
  assign new_n12318_ = ~\all_features[1751]  & (~\all_features[1750]  | ~new_n12319_ | ~new_n12314_ | ~new_n12312_);
  assign new_n12319_ = \all_features[1746]  & \all_features[1747] ;
  assign new_n12320_ = \all_features[1751]  & (\all_features[1749]  | \all_features[1750]  | \all_features[1748] );
  assign new_n12321_ = ~new_n12322_ & ~new_n12324_;
  assign new_n12322_ = ~\all_features[1749]  & new_n12323_ & ((~\all_features[1746]  & new_n12309_) | ~\all_features[1748]  | ~\all_features[1747] );
  assign new_n12323_ = ~\all_features[1750]  & ~\all_features[1751] ;
  assign new_n12324_ = ~\all_features[1751]  & ~\all_features[1750]  & ~\all_features[1749]  & ~\all_features[1747]  & ~\all_features[1748] ;
  assign new_n12325_ = ~new_n12326_ & ~new_n12327_;
  assign new_n12326_ = new_n12323_ & (~\all_features[1749]  | (~\all_features[1748]  & (~\all_features[1747]  | (~\all_features[1746]  & ~\all_features[1745] ))));
  assign new_n12327_ = new_n12323_ & (~\all_features[1747]  | ~new_n12312_ | (~\all_features[1746]  & ~new_n12314_));
  assign new_n12328_ = ~\all_features[1751]  & (~\all_features[1750]  | (~\all_features[1749]  & (new_n12309_ | ~new_n12319_ | ~\all_features[1748] )));
  assign new_n12329_ = ~\all_features[1751]  & (~\all_features[1750]  | (~\all_features[1748]  & ~\all_features[1749]  & ~new_n12319_));
  assign new_n12330_ = ~new_n12326_ & (new_n12327_ | (~new_n12329_ & (new_n12328_ | (~new_n12316_ & ~new_n12331_))));
  assign new_n12331_ = ~new_n12318_ & (~new_n12320_ | (new_n12307_ & (~new_n12311_ | (~new_n12333_ & new_n12332_))));
  assign new_n12332_ = \all_features[1751]  & ~new_n12313_ & \all_features[1750] ;
  assign new_n12333_ = \all_features[1750]  & \all_features[1751]  & (\all_features[1749]  | (\all_features[1748]  & (\all_features[1747]  | \all_features[1746] )));
  assign new_n12334_ = new_n12321_ & new_n12325_ & (new_n12335_ | new_n12316_ | new_n12328_ | ~new_n12336_);
  assign new_n12335_ = new_n12320_ & new_n12311_ & new_n12307_ & new_n12332_;
  assign new_n12336_ = ~new_n12318_ & ~new_n12329_;
  assign new_n12337_ = new_n12336_ & new_n12321_ & ~new_n12327_ & ~new_n12328_ & ~new_n12316_ & ~new_n12326_;
  assign new_n12338_ = new_n12343_ & new_n12339_ & ~new_n12353_ & ~new_n12352_ & ~new_n12349_ & ~new_n12351_;
  assign new_n12339_ = ~new_n12340_ & (\all_features[3403]  | \all_features[3404]  | \all_features[3405]  | \all_features[3406]  | \all_features[3407] );
  assign new_n12340_ = ~\all_features[3405]  & new_n12341_ & ((~\all_features[3402]  & new_n12342_) | ~\all_features[3404]  | ~\all_features[3403] );
  assign new_n12341_ = ~\all_features[3406]  & ~\all_features[3407] ;
  assign new_n12342_ = ~\all_features[3400]  & ~\all_features[3401] ;
  assign new_n12343_ = ~new_n12344_ & ~new_n12348_;
  assign new_n12344_ = ~\all_features[3407]  & (~\all_features[3406]  | ~new_n12345_ | ~new_n12346_ | ~new_n12347_);
  assign new_n12345_ = \all_features[3402]  & \all_features[3403] ;
  assign new_n12346_ = \all_features[3400]  & \all_features[3401] ;
  assign new_n12347_ = \all_features[3404]  & \all_features[3405] ;
  assign new_n12348_ = ~\all_features[3407]  & (~\all_features[3406]  | (~\all_features[3404]  & ~\all_features[3405]  & ~new_n12345_));
  assign new_n12349_ = ~new_n12350_ & ~\all_features[3407] ;
  assign new_n12350_ = \all_features[3405]  & \all_features[3406]  & (\all_features[3404]  | (\all_features[3402]  & \all_features[3403]  & \all_features[3401] ));
  assign new_n12351_ = new_n12341_ & (~\all_features[3405]  | (~\all_features[3404]  & (~\all_features[3403]  | (~\all_features[3402]  & ~\all_features[3401] ))));
  assign new_n12352_ = ~\all_features[3407]  & (~\all_features[3406]  | (~\all_features[3405]  & (new_n12342_ | ~new_n12345_ | ~\all_features[3404] )));
  assign new_n12353_ = new_n12341_ & (~\all_features[3403]  | ~new_n12347_ | (~\all_features[3402]  & ~new_n12346_));
  assign new_n12354_ = new_n12366_ & new_n12358_ & ~new_n12370_ & ~new_n12369_ & ~new_n12355_ & ~new_n12364_;
  assign new_n12355_ = ~\all_features[2391]  & (~\all_features[2390]  | new_n12356_);
  assign new_n12356_ = ~\all_features[2389]  & (new_n12357_ | ~\all_features[2387]  | ~\all_features[2388]  | ~\all_features[2386] );
  assign new_n12357_ = ~\all_features[2384]  & ~\all_features[2385] ;
  assign new_n12358_ = ~new_n12359_ & ~new_n12363_;
  assign new_n12359_ = new_n12360_ & (~\all_features[2387]  | ~new_n12362_ | (~\all_features[2386]  & ~new_n12361_));
  assign new_n12360_ = ~\all_features[2390]  & ~\all_features[2391] ;
  assign new_n12361_ = \all_features[2384]  & \all_features[2385] ;
  assign new_n12362_ = \all_features[2388]  & \all_features[2389] ;
  assign new_n12363_ = new_n12360_ & (~\all_features[2389]  | (~\all_features[2388]  & (~\all_features[2387]  | (~\all_features[2386]  & ~\all_features[2385] ))));
  assign new_n12364_ = ~new_n12365_ & ~\all_features[2391] ;
  assign new_n12365_ = \all_features[2389]  & \all_features[2390]  & (\all_features[2388]  | (\all_features[2386]  & \all_features[2387]  & \all_features[2385] ));
  assign new_n12366_ = ~new_n12367_ & ~new_n12368_;
  assign new_n12367_ = ~\all_features[2391]  & ~\all_features[2390]  & ~\all_features[2389]  & ~\all_features[2387]  & ~\all_features[2388] ;
  assign new_n12368_ = ~\all_features[2391]  & (~\all_features[2390]  | (~\all_features[2389]  & ~\all_features[2388]  & (~\all_features[2387]  | ~\all_features[2386] )));
  assign new_n12369_ = ~\all_features[2389]  & new_n12360_ & ((~\all_features[2386]  & new_n12357_) | ~\all_features[2388]  | ~\all_features[2387] );
  assign new_n12370_ = ~\all_features[2391]  & (~new_n12362_ | ~\all_features[2386]  | ~\all_features[2387]  | ~\all_features[2390]  | ~new_n12361_);
  assign new_n12371_ = new_n12372_ & new_n12373_;
  assign new_n12372_ = ~new_n9551_ & ~new_n9572_;
  assign new_n12373_ = ~new_n9579_ & ~new_n9581_;
  assign new_n12374_ = new_n12375_ & (~new_n12404_ | ~new_n12400_);
  assign new_n12375_ = ~new_n12376_ & ~new_n12398_;
  assign new_n12376_ = new_n12393_ & ~new_n12397_ & ~new_n12377_ & ~new_n12396_;
  assign new_n12377_ = new_n12378_ & (~new_n12391_ | ~new_n12392_ | ~new_n12388_ | ~new_n12390_);
  assign new_n12378_ = ~new_n12387_ & ~new_n12384_ & ~new_n12379_ & ~new_n12382_;
  assign new_n12379_ = ~\all_features[3423]  & (~\all_features[3422]  | (~\all_features[3421]  & (new_n12380_ | ~new_n12381_ | ~\all_features[3420] )));
  assign new_n12380_ = ~\all_features[3416]  & ~\all_features[3417] ;
  assign new_n12381_ = \all_features[3418]  & \all_features[3419] ;
  assign new_n12382_ = ~new_n12383_ & ~\all_features[3423] ;
  assign new_n12383_ = \all_features[3421]  & \all_features[3422]  & (\all_features[3420]  | (\all_features[3418]  & \all_features[3419]  & \all_features[3417] ));
  assign new_n12384_ = ~\all_features[3423]  & (~\all_features[3422]  | ~new_n12385_ | ~new_n12386_ | ~new_n12381_);
  assign new_n12385_ = \all_features[3420]  & \all_features[3421] ;
  assign new_n12386_ = \all_features[3416]  & \all_features[3417] ;
  assign new_n12387_ = ~\all_features[3423]  & (~\all_features[3422]  | (~\all_features[3420]  & ~\all_features[3421]  & ~new_n12381_));
  assign new_n12388_ = \all_features[3423]  & (\all_features[3422]  | (\all_features[3421]  & (\all_features[3420]  | ~new_n12380_ | ~new_n12389_)));
  assign new_n12389_ = ~\all_features[3418]  & ~\all_features[3419] ;
  assign new_n12390_ = \all_features[3423]  & (\all_features[3422]  | (new_n12385_ & (\all_features[3418]  | \all_features[3419]  | \all_features[3417] )));
  assign new_n12391_ = \all_features[3422]  & \all_features[3423]  & (\all_features[3420]  | \all_features[3421]  | new_n12386_ | ~new_n12389_);
  assign new_n12392_ = \all_features[3423]  & (\all_features[3421]  | \all_features[3422]  | \all_features[3420] );
  assign new_n12393_ = ~new_n12394_ & (\all_features[3419]  | \all_features[3420]  | \all_features[3421]  | \all_features[3422]  | \all_features[3423] );
  assign new_n12394_ = ~\all_features[3421]  & new_n12395_ & ((~\all_features[3418]  & new_n12380_) | ~\all_features[3420]  | ~\all_features[3419] );
  assign new_n12395_ = ~\all_features[3422]  & ~\all_features[3423] ;
  assign new_n12396_ = new_n12395_ & (~\all_features[3421]  | (~\all_features[3420]  & (~\all_features[3419]  | (~\all_features[3418]  & ~\all_features[3417] ))));
  assign new_n12397_ = new_n12395_ & (~\all_features[3419]  | ~new_n12385_ | (~\all_features[3418]  & ~new_n12386_));
  assign new_n12398_ = new_n12399_ & new_n12393_ & ~new_n12382_ & ~new_n12396_;
  assign new_n12399_ = ~new_n12397_ & ~new_n12387_ & ~new_n12379_ & ~new_n12384_;
  assign new_n12400_ = ~new_n12401_ & (\all_features[3419]  | \all_features[3420]  | \all_features[3421]  | \all_features[3422]  | \all_features[3423] );
  assign new_n12401_ = ~new_n12394_ & (new_n12396_ | (~new_n12397_ & (new_n12387_ | (~new_n12379_ & ~new_n12402_))));
  assign new_n12402_ = ~new_n12382_ & (new_n12384_ | (new_n12392_ & (~new_n12388_ | (~new_n12403_ & new_n12390_))));
  assign new_n12403_ = ~\all_features[3421]  & \all_features[3422]  & \all_features[3423]  & (\all_features[3420]  ? new_n12389_ : (new_n12386_ | ~new_n12389_));
  assign new_n12404_ = new_n12393_ & (new_n12397_ | new_n12396_ | (~new_n12379_ & ~new_n12387_ & ~new_n12405_));
  assign new_n12405_ = ~new_n12384_ & ~new_n12382_ & (~new_n12392_ | ~new_n12388_ | new_n12406_);
  assign new_n12406_ = new_n12390_ & new_n12391_ & (new_n12407_ | ~\all_features[3421]  | ~\all_features[3422]  | ~\all_features[3423] );
  assign new_n12407_ = ~\all_features[3419]  & ~\all_features[3420]  & (~\all_features[3418]  | new_n12380_);
  assign new_n12408_ = ~new_n12442_ & (~new_n12439_ | new_n12409_);
  assign new_n12409_ = ~new_n12410_ & (new_n12429_ | (~new_n12435_ & ~new_n12427_));
  assign new_n12410_ = new_n12426_ & (~new_n12430_ | (~new_n12411_ & ~new_n12433_ & ~new_n12434_));
  assign new_n12411_ = ~new_n12423_ & ~new_n12421_ & (~new_n12425_ | new_n12415_ | ~new_n12412_);
  assign new_n12412_ = \all_features[3679]  & (\all_features[3678]  | new_n12413_);
  assign new_n12413_ = \all_features[3677]  & (\all_features[3674]  | \all_features[3675]  | \all_features[3676]  | ~new_n12414_);
  assign new_n12414_ = ~\all_features[3672]  & ~\all_features[3673] ;
  assign new_n12415_ = ~new_n12418_ & new_n12416_ & \all_features[3678]  & \all_features[3679]  & (~\all_features[3677]  | new_n12420_);
  assign new_n12416_ = \all_features[3679]  & (\all_features[3678]  | (new_n12417_ & (\all_features[3674]  | \all_features[3675]  | \all_features[3673] )));
  assign new_n12417_ = \all_features[3676]  & \all_features[3677] ;
  assign new_n12418_ = ~\all_features[3677]  & ~\all_features[3676]  & ~\all_features[3675]  & ~new_n12419_ & ~\all_features[3674] ;
  assign new_n12419_ = \all_features[3672]  & \all_features[3673] ;
  assign new_n12420_ = ~\all_features[3675]  & ~\all_features[3676]  & (~\all_features[3674]  | new_n12414_);
  assign new_n12421_ = ~new_n12422_ & ~\all_features[3679] ;
  assign new_n12422_ = \all_features[3677]  & \all_features[3678]  & (\all_features[3676]  | (\all_features[3674]  & \all_features[3675]  & \all_features[3673] ));
  assign new_n12423_ = ~\all_features[3679]  & (~\all_features[3678]  | ~new_n12424_ | ~new_n12419_ | ~new_n12417_);
  assign new_n12424_ = \all_features[3674]  & \all_features[3675] ;
  assign new_n12425_ = \all_features[3679]  & (\all_features[3677]  | \all_features[3678]  | \all_features[3676] );
  assign new_n12426_ = ~new_n12427_ & ~new_n12429_;
  assign new_n12427_ = ~\all_features[3677]  & new_n12428_ & ((~\all_features[3674]  & new_n12414_) | ~\all_features[3676]  | ~\all_features[3675] );
  assign new_n12428_ = ~\all_features[3678]  & ~\all_features[3679] ;
  assign new_n12429_ = ~\all_features[3679]  & ~\all_features[3678]  & ~\all_features[3677]  & ~\all_features[3675]  & ~\all_features[3676] ;
  assign new_n12430_ = ~new_n12431_ & ~new_n12432_;
  assign new_n12431_ = new_n12428_ & (~\all_features[3677]  | (~\all_features[3676]  & (~\all_features[3675]  | (~\all_features[3674]  & ~\all_features[3673] ))));
  assign new_n12432_ = new_n12428_ & (~\all_features[3675]  | ~new_n12417_ | (~\all_features[3674]  & ~new_n12419_));
  assign new_n12433_ = ~\all_features[3679]  & (~\all_features[3678]  | (~\all_features[3677]  & (new_n12414_ | ~new_n12424_ | ~\all_features[3676] )));
  assign new_n12434_ = ~\all_features[3679]  & (~\all_features[3678]  | (~\all_features[3676]  & ~\all_features[3677]  & ~new_n12424_));
  assign new_n12435_ = ~new_n12431_ & (new_n12432_ | (~new_n12434_ & (new_n12433_ | (~new_n12421_ & ~new_n12436_))));
  assign new_n12436_ = ~new_n12423_ & (~new_n12425_ | (new_n12412_ & (~new_n12416_ | (~new_n12438_ & new_n12437_))));
  assign new_n12437_ = \all_features[3679]  & ~new_n12418_ & \all_features[3678] ;
  assign new_n12438_ = \all_features[3678]  & \all_features[3679]  & (\all_features[3677]  | (\all_features[3676]  & (\all_features[3675]  | \all_features[3674] )));
  assign new_n12439_ = new_n12426_ & new_n12430_ & (new_n12440_ | new_n12421_ | new_n12433_ | ~new_n12441_);
  assign new_n12440_ = new_n12425_ & new_n12416_ & new_n12412_ & new_n12437_;
  assign new_n12441_ = ~new_n12423_ & ~new_n12434_;
  assign new_n12442_ = new_n12441_ & new_n12426_ & ~new_n12432_ & ~new_n12433_ & ~new_n12421_ & ~new_n12431_;
  assign new_n12443_ = ~new_n12444_ & new_n10240_;
  assign new_n12444_ = ~new_n10238_ & ~new_n10229_;
  assign new_n12445_ = (~new_n12354_ | new_n12264_ | (new_n8590_ & ~new_n12446_)) & (new_n12447_ | ~new_n12267_ | ~new_n12264_);
  assign new_n12446_ = ~new_n8559_ & ~new_n8580_;
  assign new_n12447_ = new_n12448_ & new_n10681_;
  assign new_n12448_ = ~new_n9101_ & ~new_n9122_;
  assign new_n12449_ = (~new_n12371_ | ~new_n12450_ | new_n12338_) & (new_n12264_ | new_n12354_ | ~new_n12303_ | ~new_n12338_);
  assign new_n12450_ = new_n12374_ & new_n12408_;
  assign new_n12451_ = new_n12561_ & (new_n6879_ | (new_n12452_ & new_n12686_) | (new_n12527_ & ~new_n12686_));
  assign new_n12452_ = new_n9457_ ? new_n12453_ : (new_n12525_ | (~new_n12491_ & new_n12523_));
  assign new_n12453_ = new_n12454_ & new_n12486_;
  assign new_n12454_ = new_n12455_ & new_n12476_;
  assign new_n12455_ = ~new_n12456_ & (\all_features[4123]  | \all_features[4124]  | \all_features[4125]  | \all_features[4126]  | \all_features[4127] );
  assign new_n12456_ = ~new_n12470_ & (new_n12472_ | (~new_n12473_ & (new_n12474_ | (~new_n12457_ & ~new_n12475_))));
  assign new_n12457_ = ~new_n12465_ & (new_n12467_ | (~new_n12458_ & new_n12469_));
  assign new_n12458_ = \all_features[4127]  & ((~new_n12463_ & ~\all_features[4125]  & \all_features[4126] ) | (~new_n12461_ & (\all_features[4126]  | (~new_n12459_ & \all_features[4125] ))));
  assign new_n12459_ = new_n12460_ & ~\all_features[4124]  & ~\all_features[4122]  & ~\all_features[4123] ;
  assign new_n12460_ = ~\all_features[4120]  & ~\all_features[4121] ;
  assign new_n12461_ = \all_features[4127]  & (\all_features[4126]  | (new_n12462_ & (\all_features[4122]  | \all_features[4123]  | \all_features[4121] )));
  assign new_n12462_ = \all_features[4124]  & \all_features[4125] ;
  assign new_n12463_ = (\all_features[4124]  & (\all_features[4122]  | \all_features[4123] )) | (~new_n12464_ & ~\all_features[4122]  & ~\all_features[4123]  & ~\all_features[4124] );
  assign new_n12464_ = \all_features[4120]  & \all_features[4121] ;
  assign new_n12465_ = ~new_n12466_ & ~\all_features[4127] ;
  assign new_n12466_ = \all_features[4125]  & \all_features[4126]  & (\all_features[4124]  | (\all_features[4122]  & \all_features[4123]  & \all_features[4121] ));
  assign new_n12467_ = ~\all_features[4127]  & (~\all_features[4126]  | ~new_n12464_ | ~new_n12462_ | ~new_n12468_);
  assign new_n12468_ = \all_features[4122]  & \all_features[4123] ;
  assign new_n12469_ = \all_features[4127]  & (\all_features[4125]  | \all_features[4126]  | \all_features[4124] );
  assign new_n12470_ = ~\all_features[4125]  & new_n12471_ & ((~\all_features[4122]  & new_n12460_) | ~\all_features[4124]  | ~\all_features[4123] );
  assign new_n12471_ = ~\all_features[4126]  & ~\all_features[4127] ;
  assign new_n12472_ = new_n12471_ & (~\all_features[4125]  | (~\all_features[4124]  & (~\all_features[4123]  | (~\all_features[4122]  & ~\all_features[4121] ))));
  assign new_n12473_ = new_n12471_ & (~\all_features[4123]  | ~new_n12462_ | (~\all_features[4122]  & ~new_n12464_));
  assign new_n12474_ = ~\all_features[4127]  & (~\all_features[4126]  | (~\all_features[4124]  & ~\all_features[4125]  & ~new_n12468_));
  assign new_n12475_ = ~\all_features[4127]  & (~\all_features[4126]  | (~\all_features[4125]  & (new_n12460_ | ~new_n12468_ | ~\all_features[4124] )));
  assign new_n12476_ = new_n12482_ & (~new_n12483_ | (new_n12484_ & (~new_n12485_ | new_n12477_)));
  assign new_n12477_ = new_n12478_ & (~new_n12479_ | (~new_n12481_ & \all_features[4125]  & \all_features[4126]  & \all_features[4127] ));
  assign new_n12478_ = \all_features[4127]  & (\all_features[4126]  | (~new_n12459_ & \all_features[4125] ));
  assign new_n12479_ = \all_features[4127]  & \all_features[4126]  & ~new_n12480_ & new_n12461_;
  assign new_n12480_ = ~\all_features[4125]  & ~\all_features[4124]  & ~\all_features[4123]  & ~new_n12464_ & ~\all_features[4122] ;
  assign new_n12481_ = ~\all_features[4123]  & ~\all_features[4124]  & (~\all_features[4122]  | new_n12460_);
  assign new_n12482_ = ~new_n12470_ & (\all_features[4123]  | \all_features[4124]  | \all_features[4125]  | \all_features[4126]  | \all_features[4127] );
  assign new_n12483_ = ~new_n12472_ & ~new_n12473_;
  assign new_n12484_ = ~new_n12474_ & ~new_n12475_;
  assign new_n12485_ = ~new_n12465_ & ~new_n12467_;
  assign new_n12486_ = new_n12487_ & new_n12490_;
  assign new_n12487_ = new_n12488_ & (new_n12475_ | new_n12465_ | ~new_n12489_ | (new_n12479_ & new_n12478_));
  assign new_n12488_ = new_n12482_ & new_n12483_;
  assign new_n12489_ = ~new_n12474_ & ~new_n12467_;
  assign new_n12490_ = new_n12485_ & new_n12488_ & new_n12484_;
  assign new_n12491_ = ~new_n12492_ & ~new_n12514_;
  assign new_n12492_ = ~new_n12513_ & (new_n12509_ | (~new_n12511_ & (new_n12512_ | (~new_n12493_ & ~new_n12508_))));
  assign new_n12493_ = ~new_n12502_ & (new_n12505_ | (~new_n12504_ & (~new_n12507_ | (~new_n12494_ & new_n12500_))));
  assign new_n12494_ = new_n12495_ & (\all_features[4549]  | ~new_n12498_ | (~new_n12499_ & ~\all_features[4548]  & new_n12497_) | (\all_features[4548]  & ~new_n12497_));
  assign new_n12495_ = \all_features[4551]  & (\all_features[4550]  | (new_n12496_ & (\all_features[4546]  | \all_features[4547]  | \all_features[4545] )));
  assign new_n12496_ = \all_features[4548]  & \all_features[4549] ;
  assign new_n12497_ = ~\all_features[4546]  & ~\all_features[4547] ;
  assign new_n12498_ = \all_features[4550]  & \all_features[4551] ;
  assign new_n12499_ = \all_features[4544]  & \all_features[4545] ;
  assign new_n12500_ = \all_features[4551]  & (\all_features[4550]  | (\all_features[4549]  & (\all_features[4548]  | ~new_n12501_ | ~new_n12497_)));
  assign new_n12501_ = ~\all_features[4544]  & ~\all_features[4545] ;
  assign new_n12502_ = ~\all_features[4551]  & (~\all_features[4550]  | (~\all_features[4549]  & (new_n12501_ | ~new_n12503_ | ~\all_features[4548] )));
  assign new_n12503_ = \all_features[4546]  & \all_features[4547] ;
  assign new_n12504_ = ~\all_features[4551]  & (~\all_features[4550]  | ~new_n12496_ | ~new_n12499_ | ~new_n12503_);
  assign new_n12505_ = ~new_n12506_ & ~\all_features[4551] ;
  assign new_n12506_ = \all_features[4549]  & \all_features[4550]  & (\all_features[4548]  | (\all_features[4546]  & \all_features[4547]  & \all_features[4545] ));
  assign new_n12507_ = \all_features[4551]  & (\all_features[4549]  | \all_features[4550]  | \all_features[4548] );
  assign new_n12508_ = ~\all_features[4551]  & (~\all_features[4550]  | (~\all_features[4548]  & ~\all_features[4549]  & ~new_n12503_));
  assign new_n12509_ = ~\all_features[4549]  & new_n12510_ & ((~\all_features[4546]  & new_n12501_) | ~\all_features[4548]  | ~\all_features[4547] );
  assign new_n12510_ = ~\all_features[4550]  & ~\all_features[4551] ;
  assign new_n12511_ = new_n12510_ & (~\all_features[4549]  | (~\all_features[4548]  & (~\all_features[4547]  | (~\all_features[4546]  & ~\all_features[4545] ))));
  assign new_n12512_ = new_n12510_ & (~\all_features[4547]  | ~new_n12496_ | (~\all_features[4546]  & ~new_n12499_));
  assign new_n12513_ = ~\all_features[4551]  & ~\all_features[4550]  & ~\all_features[4549]  & ~\all_features[4547]  & ~\all_features[4548] ;
  assign new_n12514_ = new_n12521_ & (~new_n12522_ | (new_n12519_ & (~new_n12520_ | new_n12515_)));
  assign new_n12515_ = new_n12507_ & ~new_n12516_ & new_n12500_;
  assign new_n12516_ = new_n12517_ & new_n12495_ & (~\all_features[4549]  | ~new_n12498_ | new_n12518_);
  assign new_n12517_ = new_n12498_ & (new_n12499_ | \all_features[4548]  | \all_features[4549]  | ~new_n12497_);
  assign new_n12518_ = ~\all_features[4547]  & ~\all_features[4548]  & (~\all_features[4546]  | new_n12501_);
  assign new_n12519_ = ~new_n12502_ & ~new_n12508_;
  assign new_n12520_ = ~new_n12504_ & ~new_n12505_;
  assign new_n12521_ = ~new_n12509_ & ~new_n12513_;
  assign new_n12522_ = ~new_n12511_ & ~new_n12512_;
  assign new_n12523_ = new_n12522_ & new_n12521_ & (~new_n12520_ | ~new_n12519_ | (new_n12524_ & new_n12500_));
  assign new_n12524_ = new_n12507_ & new_n12495_ & new_n12517_;
  assign new_n12525_ = new_n12526_ & ~new_n12513_ & ~new_n12511_ & ~new_n12504_ & ~new_n12505_;
  assign new_n12526_ = ~new_n12512_ & ~new_n12509_ & ~new_n12502_ & ~new_n12508_;
  assign new_n12527_ = new_n12528_ ? ~new_n12537_ : new_n12535_;
  assign new_n12528_ = ~new_n12529_ & new_n12534_;
  assign new_n12529_ = new_n9271_ & new_n12530_;
  assign new_n12530_ = ~new_n12531_ & (\all_features[3003]  | \all_features[3004]  | \all_features[3005]  | \all_features[3006]  | \all_features[3007] );
  assign new_n12531_ = ~new_n9252_ & (new_n9255_ | (~new_n9256_ & (new_n9265_ | (~new_n9260_ & ~new_n12532_))));
  assign new_n12532_ = ~new_n9262_ & (new_n9264_ | (new_n9270_ & (~new_n9266_ | (~new_n12533_ & new_n9268_))));
  assign new_n12533_ = ~\all_features[3005]  & \all_features[3006]  & \all_features[3007]  & (\all_features[3004]  ? new_n9267_ : (new_n9258_ | ~new_n9267_));
  assign new_n12534_ = ~new_n9249_ & ~new_n9275_;
  assign new_n12535_ = new_n12536_ & new_n7665_;
  assign new_n12536_ = new_n7637_ & new_n7659_;
  assign new_n12537_ = ~new_n12538_ & ~new_n12560_;
  assign new_n12538_ = new_n12539_ & (~new_n12548_ | (new_n12558_ & new_n12559_ & new_n12555_ & new_n12557_));
  assign new_n12539_ = new_n12540_ & ~new_n12544_ & ~new_n12545_;
  assign new_n12540_ = ~new_n12541_ & (\all_features[3531]  | \all_features[3532]  | \all_features[3533]  | \all_features[3534]  | \all_features[3535] );
  assign new_n12541_ = ~\all_features[3533]  & new_n12543_ & ((~\all_features[3530]  & new_n12542_) | ~\all_features[3532]  | ~\all_features[3531] );
  assign new_n12542_ = ~\all_features[3528]  & ~\all_features[3529] ;
  assign new_n12543_ = ~\all_features[3534]  & ~\all_features[3535] ;
  assign new_n12544_ = new_n12543_ & (~\all_features[3533]  | (~\all_features[3532]  & (~\all_features[3531]  | (~\all_features[3530]  & ~\all_features[3529] ))));
  assign new_n12545_ = new_n12543_ & (~\all_features[3531]  | ~new_n12546_ | (~\all_features[3530]  & ~new_n12547_));
  assign new_n12546_ = \all_features[3532]  & \all_features[3533] ;
  assign new_n12547_ = \all_features[3528]  & \all_features[3529] ;
  assign new_n12548_ = ~new_n12554_ & ~new_n12553_ & ~new_n12549_ & ~new_n12551_;
  assign new_n12549_ = ~\all_features[3535]  & (~\all_features[3534]  | (~\all_features[3533]  & (new_n12542_ | ~new_n12550_ | ~\all_features[3532] )));
  assign new_n12550_ = \all_features[3530]  & \all_features[3531] ;
  assign new_n12551_ = ~new_n12552_ & ~\all_features[3535] ;
  assign new_n12552_ = \all_features[3533]  & \all_features[3534]  & (\all_features[3532]  | (\all_features[3530]  & \all_features[3531]  & \all_features[3529] ));
  assign new_n12553_ = ~\all_features[3535]  & (~\all_features[3534]  | ~new_n12546_ | ~new_n12547_ | ~new_n12550_);
  assign new_n12554_ = ~\all_features[3535]  & (~\all_features[3534]  | (~\all_features[3532]  & ~\all_features[3533]  & ~new_n12550_));
  assign new_n12555_ = \all_features[3535]  & (\all_features[3534]  | (\all_features[3533]  & (\all_features[3532]  | ~new_n12542_ | ~new_n12556_)));
  assign new_n12556_ = ~\all_features[3530]  & ~\all_features[3531] ;
  assign new_n12557_ = \all_features[3535]  & (\all_features[3534]  | (new_n12546_ & (\all_features[3530]  | \all_features[3531]  | \all_features[3529] )));
  assign new_n12558_ = \all_features[3534]  & \all_features[3535]  & (\all_features[3532]  | \all_features[3533]  | new_n12547_ | ~new_n12556_);
  assign new_n12559_ = \all_features[3535]  & (\all_features[3533]  | \all_features[3534]  | \all_features[3532] );
  assign new_n12560_ = new_n12539_ & new_n12548_;
  assign new_n12561_ = ~new_n12599_ & (new_n12600_ | ~new_n6879_ | (new_n12597_ ? new_n12562_ : ~new_n7671_));
  assign new_n12562_ = new_n12563_ & ~new_n12592_ & ~new_n12595_;
  assign new_n12563_ = ~new_n12564_ & ~new_n12588_;
  assign new_n12564_ = new_n12579_ & (~new_n12584_ | (~new_n12582_ & ~new_n12565_ & ~new_n12587_));
  assign new_n12565_ = ~new_n12577_ & ~new_n12575_ & (~new_n12578_ | ~new_n12574_ | new_n12566_);
  assign new_n12566_ = new_n12567_ & new_n12569_ & (new_n12572_ | ~\all_features[5453]  | ~\all_features[5454]  | ~\all_features[5455] );
  assign new_n12567_ = \all_features[5455]  & (\all_features[5454]  | (new_n12568_ & (\all_features[5450]  | \all_features[5451]  | \all_features[5449] )));
  assign new_n12568_ = \all_features[5452]  & \all_features[5453] ;
  assign new_n12569_ = \all_features[5454]  & \all_features[5455]  & (\all_features[5452]  | \all_features[5453]  | new_n12571_ | ~new_n12570_);
  assign new_n12570_ = ~\all_features[5450]  & ~\all_features[5451] ;
  assign new_n12571_ = \all_features[5448]  & \all_features[5449] ;
  assign new_n12572_ = ~\all_features[5451]  & ~\all_features[5452]  & (~\all_features[5450]  | new_n12573_);
  assign new_n12573_ = ~\all_features[5448]  & ~\all_features[5449] ;
  assign new_n12574_ = \all_features[5455]  & (\all_features[5454]  | (\all_features[5453]  & (\all_features[5452]  | ~new_n12570_ | ~new_n12573_)));
  assign new_n12575_ = ~new_n12576_ & ~\all_features[5455] ;
  assign new_n12576_ = \all_features[5453]  & \all_features[5454]  & (\all_features[5452]  | (\all_features[5450]  & \all_features[5451]  & \all_features[5449] ));
  assign new_n12577_ = ~\all_features[5455]  & (~new_n12571_ | ~\all_features[5450]  | ~\all_features[5451]  | ~\all_features[5454]  | ~new_n12568_);
  assign new_n12578_ = \all_features[5455]  & (\all_features[5453]  | \all_features[5454]  | \all_features[5452] );
  assign new_n12579_ = ~new_n12580_ & (\all_features[5451]  | \all_features[5452]  | \all_features[5453]  | \all_features[5454]  | \all_features[5455] );
  assign new_n12580_ = ~\all_features[5453]  & new_n12581_ & ((~\all_features[5450]  & new_n12573_) | ~\all_features[5452]  | ~\all_features[5451] );
  assign new_n12581_ = ~\all_features[5454]  & ~\all_features[5455] ;
  assign new_n12582_ = ~\all_features[5455]  & (~\all_features[5454]  | new_n12583_);
  assign new_n12583_ = ~\all_features[5453]  & (new_n12573_ | ~\all_features[5451]  | ~\all_features[5452]  | ~\all_features[5450] );
  assign new_n12584_ = ~new_n12585_ & ~new_n12586_;
  assign new_n12585_ = new_n12581_ & (~\all_features[5451]  | ~new_n12568_ | (~new_n12571_ & ~\all_features[5450] ));
  assign new_n12586_ = new_n12581_ & (~\all_features[5453]  | (~\all_features[5452]  & (~\all_features[5451]  | (~\all_features[5450]  & ~\all_features[5449] ))));
  assign new_n12587_ = ~\all_features[5455]  & (~\all_features[5454]  | (~\all_features[5453]  & ~\all_features[5452]  & (~\all_features[5451]  | ~\all_features[5450] )));
  assign new_n12588_ = ~new_n12589_ & (\all_features[5451]  | \all_features[5452]  | \all_features[5453]  | \all_features[5454]  | \all_features[5455] );
  assign new_n12589_ = ~new_n12580_ & (new_n12586_ | (~new_n12585_ & (new_n12587_ | (~new_n12582_ & ~new_n12590_))));
  assign new_n12590_ = ~new_n12575_ & (new_n12577_ | (new_n12578_ & (~new_n12574_ | (~new_n12591_ & new_n12567_))));
  assign new_n12591_ = ~\all_features[5453]  & \all_features[5454]  & \all_features[5455]  & (\all_features[5452]  ? new_n12570_ : (new_n12571_ | ~new_n12570_));
  assign new_n12592_ = new_n12584_ & ~new_n12593_ & new_n12579_;
  assign new_n12593_ = ~new_n12587_ & ~new_n12577_ & ~new_n12575_ & ~new_n12582_ & ~new_n12594_;
  assign new_n12594_ = new_n12578_ & new_n12574_ & new_n12567_ & new_n12569_;
  assign new_n12595_ = new_n12579_ & new_n12596_ & ~new_n12575_ & ~new_n12586_;
  assign new_n12596_ = ~new_n12587_ & ~new_n12585_ & ~new_n12582_ & ~new_n12577_;
  assign new_n12597_ = new_n10874_ & new_n12598_;
  assign new_n12598_ = ~new_n8385_ & ~new_n8388_;
  assign new_n12599_ = ~new_n12655_ & ~new_n12685_ & new_n12600_ & new_n6879_ & (~new_n12682_ | new_n12626_);
  assign new_n12600_ = ~new_n12601_ & ~new_n12624_;
  assign new_n12601_ = new_n12619_ & ~new_n12623_ & ~new_n12602_ & ~new_n12622_;
  assign new_n12602_ = ~new_n12617_ & ~new_n12618_ & new_n12610_ & (~new_n12615_ | ~new_n12603_);
  assign new_n12603_ = new_n12609_ & new_n12604_ & new_n12606_;
  assign new_n12604_ = \all_features[4575]  & (\all_features[4574]  | (new_n12605_ & (\all_features[4570]  | \all_features[4571]  | \all_features[4569] )));
  assign new_n12605_ = \all_features[4572]  & \all_features[4573] ;
  assign new_n12606_ = \all_features[4574]  & \all_features[4575]  & (\all_features[4572]  | \all_features[4573]  | new_n12608_ | ~new_n12607_);
  assign new_n12607_ = ~\all_features[4570]  & ~\all_features[4571] ;
  assign new_n12608_ = \all_features[4568]  & \all_features[4569] ;
  assign new_n12609_ = \all_features[4575]  & (\all_features[4573]  | \all_features[4574]  | \all_features[4572] );
  assign new_n12610_ = ~new_n12611_ & ~new_n12613_;
  assign new_n12611_ = ~new_n12612_ & ~\all_features[4575] ;
  assign new_n12612_ = \all_features[4573]  & \all_features[4574]  & (\all_features[4572]  | (\all_features[4570]  & \all_features[4571]  & \all_features[4569] ));
  assign new_n12613_ = ~\all_features[4575]  & (~\all_features[4574]  | (~\all_features[4572]  & ~\all_features[4573]  & ~new_n12614_));
  assign new_n12614_ = \all_features[4570]  & \all_features[4571] ;
  assign new_n12615_ = \all_features[4575]  & (\all_features[4574]  | (\all_features[4573]  & (\all_features[4572]  | ~new_n12616_ | ~new_n12607_)));
  assign new_n12616_ = ~\all_features[4568]  & ~\all_features[4569] ;
  assign new_n12617_ = ~\all_features[4575]  & (~\all_features[4574]  | (~\all_features[4573]  & (new_n12616_ | ~new_n12614_ | ~\all_features[4572] )));
  assign new_n12618_ = ~\all_features[4575]  & (~\all_features[4574]  | ~new_n12605_ | ~new_n12608_ | ~new_n12614_);
  assign new_n12619_ = ~new_n12620_ & (\all_features[4571]  | \all_features[4572]  | \all_features[4573]  | \all_features[4574]  | \all_features[4575] );
  assign new_n12620_ = ~\all_features[4573]  & new_n12621_ & ((~\all_features[4570]  & new_n12616_) | ~\all_features[4572]  | ~\all_features[4571] );
  assign new_n12621_ = ~\all_features[4574]  & ~\all_features[4575] ;
  assign new_n12622_ = new_n12621_ & (~\all_features[4573]  | (~\all_features[4572]  & (~\all_features[4571]  | (~\all_features[4570]  & ~\all_features[4569] ))));
  assign new_n12623_ = new_n12621_ & (~\all_features[4571]  | ~new_n12605_ | (~\all_features[4570]  & ~new_n12608_));
  assign new_n12624_ = new_n12619_ & new_n12610_ & new_n12625_ & ~new_n12617_ & ~new_n12618_;
  assign new_n12625_ = ~new_n12622_ & ~new_n12623_;
  assign new_n12626_ = ~new_n12627_ & ~new_n12651_;
  assign new_n12627_ = new_n12643_ & (~new_n12646_ | (~new_n12628_ & ~new_n12649_ & ~new_n12650_));
  assign new_n12628_ = ~new_n12640_ & ~new_n12638_ & (~new_n12642_ | ~new_n12637_ | new_n12629_);
  assign new_n12629_ = new_n12630_ & new_n12632_ & (new_n12635_ | ~\all_features[5237]  | ~\all_features[5238]  | ~\all_features[5239] );
  assign new_n12630_ = \all_features[5239]  & (\all_features[5238]  | (new_n12631_ & (\all_features[5234]  | \all_features[5235]  | \all_features[5233] )));
  assign new_n12631_ = \all_features[5236]  & \all_features[5237] ;
  assign new_n12632_ = \all_features[5238]  & \all_features[5239]  & (\all_features[5236]  | \all_features[5237]  | new_n12634_ | ~new_n12633_);
  assign new_n12633_ = ~\all_features[5234]  & ~\all_features[5235] ;
  assign new_n12634_ = \all_features[5232]  & \all_features[5233] ;
  assign new_n12635_ = ~\all_features[5235]  & ~\all_features[5236]  & (~\all_features[5234]  | new_n12636_);
  assign new_n12636_ = ~\all_features[5232]  & ~\all_features[5233] ;
  assign new_n12637_ = \all_features[5239]  & (\all_features[5238]  | (\all_features[5237]  & (\all_features[5236]  | ~new_n12636_ | ~new_n12633_)));
  assign new_n12638_ = ~new_n12639_ & ~\all_features[5239] ;
  assign new_n12639_ = \all_features[5237]  & \all_features[5238]  & (\all_features[5236]  | (\all_features[5234]  & \all_features[5235]  & \all_features[5233] ));
  assign new_n12640_ = ~\all_features[5239]  & (~\all_features[5238]  | ~new_n12631_ | ~new_n12634_ | ~new_n12641_);
  assign new_n12641_ = \all_features[5234]  & \all_features[5235] ;
  assign new_n12642_ = \all_features[5239]  & (\all_features[5237]  | \all_features[5238]  | \all_features[5236] );
  assign new_n12643_ = ~new_n12644_ & (\all_features[5235]  | \all_features[5236]  | \all_features[5237]  | \all_features[5238]  | \all_features[5239] );
  assign new_n12644_ = ~\all_features[5237]  & new_n12645_ & ((~\all_features[5234]  & new_n12636_) | ~\all_features[5236]  | ~\all_features[5235] );
  assign new_n12645_ = ~\all_features[5238]  & ~\all_features[5239] ;
  assign new_n12646_ = ~new_n12647_ & ~new_n12648_;
  assign new_n12647_ = new_n12645_ & (~\all_features[5237]  | (~\all_features[5236]  & (~\all_features[5235]  | (~\all_features[5234]  & ~\all_features[5233] ))));
  assign new_n12648_ = new_n12645_ & (~\all_features[5235]  | ~new_n12631_ | (~\all_features[5234]  & ~new_n12634_));
  assign new_n12649_ = ~\all_features[5239]  & (~\all_features[5238]  | (~\all_features[5237]  & (new_n12636_ | ~new_n12641_ | ~\all_features[5236] )));
  assign new_n12650_ = ~\all_features[5239]  & (~\all_features[5238]  | (~\all_features[5236]  & ~\all_features[5237]  & ~new_n12641_));
  assign new_n12651_ = ~new_n12652_ & (\all_features[5235]  | \all_features[5236]  | \all_features[5237]  | \all_features[5238]  | \all_features[5239] );
  assign new_n12652_ = ~new_n12644_ & (new_n12647_ | (~new_n12648_ & (new_n12650_ | (~new_n12649_ & ~new_n12653_))));
  assign new_n12653_ = ~new_n12638_ & (new_n12640_ | (new_n12642_ & (~new_n12637_ | (~new_n12654_ & new_n12630_))));
  assign new_n12654_ = ~\all_features[5237]  & \all_features[5238]  & \all_features[5239]  & (\all_features[5236]  ? new_n12633_ : (new_n12634_ | ~new_n12633_));
  assign new_n12655_ = new_n12656_ & new_n12680_;
  assign new_n12656_ = new_n12674_ & ~new_n12679_ & ~new_n12657_ & ~new_n12678_;
  assign new_n12657_ = ~new_n12672_ & ~new_n12673_ & new_n12667_ & (~new_n12661_ | ~new_n12658_);
  assign new_n12658_ = \all_features[3783]  & (\all_features[3782]  | new_n12659_);
  assign new_n12659_ = \all_features[3781]  & (\all_features[3778]  | \all_features[3779]  | \all_features[3780]  | ~new_n12660_);
  assign new_n12660_ = ~\all_features[3776]  & ~\all_features[3777] ;
  assign new_n12661_ = new_n12666_ & new_n12662_ & new_n12664_;
  assign new_n12662_ = \all_features[3783]  & (\all_features[3782]  | (new_n12663_ & (\all_features[3778]  | \all_features[3779]  | \all_features[3777] )));
  assign new_n12663_ = \all_features[3780]  & \all_features[3781] ;
  assign new_n12664_ = \all_features[3783]  & ~new_n12665_ & \all_features[3782] ;
  assign new_n12665_ = ~\all_features[3778]  & ~\all_features[3779]  & ~\all_features[3780]  & ~\all_features[3781]  & (~\all_features[3777]  | ~\all_features[3776] );
  assign new_n12666_ = \all_features[3783]  & (\all_features[3781]  | \all_features[3782]  | \all_features[3780] );
  assign new_n12667_ = ~new_n12668_ & ~new_n12670_;
  assign new_n12668_ = ~new_n12669_ & ~\all_features[3783] ;
  assign new_n12669_ = \all_features[3781]  & \all_features[3782]  & (\all_features[3780]  | (\all_features[3778]  & \all_features[3779]  & \all_features[3777] ));
  assign new_n12670_ = ~\all_features[3783]  & (~\all_features[3782]  | (~\all_features[3780]  & ~\all_features[3781]  & ~new_n12671_));
  assign new_n12671_ = \all_features[3778]  & \all_features[3779] ;
  assign new_n12672_ = ~\all_features[3783]  & (~\all_features[3782]  | (~\all_features[3781]  & (new_n12660_ | ~new_n12671_ | ~\all_features[3780] )));
  assign new_n12673_ = ~\all_features[3783]  & (~new_n12671_ | ~\all_features[3776]  | ~\all_features[3777]  | ~\all_features[3782]  | ~new_n12663_);
  assign new_n12674_ = ~new_n12675_ & ~new_n12677_;
  assign new_n12675_ = ~\all_features[3781]  & new_n12676_ & ((~\all_features[3778]  & new_n12660_) | ~\all_features[3780]  | ~\all_features[3779] );
  assign new_n12676_ = ~\all_features[3782]  & ~\all_features[3783] ;
  assign new_n12677_ = ~\all_features[3783]  & ~\all_features[3782]  & ~\all_features[3781]  & ~\all_features[3779]  & ~\all_features[3780] ;
  assign new_n12678_ = new_n12676_ & (~\all_features[3781]  | (~\all_features[3780]  & (~\all_features[3779]  | (~\all_features[3778]  & ~\all_features[3777] ))));
  assign new_n12679_ = new_n12676_ & (~new_n12663_ | ~\all_features[3779]  | (~\all_features[3778]  & (~\all_features[3776]  | ~\all_features[3777] )));
  assign new_n12680_ = new_n12674_ & new_n12667_ & new_n12681_ & ~new_n12672_ & ~new_n12673_;
  assign new_n12681_ = ~new_n12678_ & ~new_n12679_;
  assign new_n12682_ = new_n12643_ & new_n12646_ & (new_n12683_ | new_n12649_ | new_n12638_ | ~new_n12684_);
  assign new_n12683_ = new_n12642_ & new_n12632_ & new_n12637_ & new_n12630_;
  assign new_n12684_ = ~new_n12640_ & ~new_n12650_;
  assign new_n12685_ = new_n12643_ & new_n12684_ & ~new_n12648_ & ~new_n12647_ & ~new_n12649_ & ~new_n12638_;
  assign new_n12686_ = ~new_n12687_ & new_n12717_;
  assign new_n12687_ = ~new_n12688_ & ~new_n12709_;
  assign new_n12688_ = ~new_n12689_ & (\all_features[2139]  | \all_features[2140]  | \all_features[2141]  | \all_features[2142]  | \all_features[2143] );
  assign new_n12689_ = ~new_n12703_ & (new_n12708_ | (~new_n12705_ & (new_n12706_ | (~new_n12707_ & ~new_n12690_))));
  assign new_n12690_ = ~new_n12691_ & (new_n12700_ | (new_n12702_ & (~new_n12693_ | (~new_n12698_ & new_n12696_))));
  assign new_n12691_ = ~new_n12692_ & ~\all_features[2143] ;
  assign new_n12692_ = \all_features[2141]  & \all_features[2142]  & (\all_features[2140]  | (\all_features[2138]  & \all_features[2139]  & \all_features[2137] ));
  assign new_n12693_ = \all_features[2143]  & (\all_features[2142]  | (\all_features[2141]  & (\all_features[2140]  | ~new_n12695_ | ~new_n12694_)));
  assign new_n12694_ = ~\all_features[2136]  & ~\all_features[2137] ;
  assign new_n12695_ = ~\all_features[2138]  & ~\all_features[2139] ;
  assign new_n12696_ = \all_features[2143]  & (\all_features[2142]  | (new_n12697_ & (\all_features[2138]  | \all_features[2139]  | \all_features[2137] )));
  assign new_n12697_ = \all_features[2140]  & \all_features[2141] ;
  assign new_n12698_ = ~\all_features[2141]  & \all_features[2142]  & \all_features[2143]  & (\all_features[2140]  ? new_n12695_ : (new_n12699_ | ~new_n12695_));
  assign new_n12699_ = \all_features[2136]  & \all_features[2137] ;
  assign new_n12700_ = ~\all_features[2143]  & (~\all_features[2142]  | ~new_n12699_ | ~new_n12697_ | ~new_n12701_);
  assign new_n12701_ = \all_features[2138]  & \all_features[2139] ;
  assign new_n12702_ = \all_features[2143]  & (\all_features[2141]  | \all_features[2142]  | \all_features[2140] );
  assign new_n12703_ = ~\all_features[2141]  & new_n12704_ & ((~\all_features[2138]  & new_n12694_) | ~\all_features[2140]  | ~\all_features[2139] );
  assign new_n12704_ = ~\all_features[2142]  & ~\all_features[2143] ;
  assign new_n12705_ = new_n12704_ & (~\all_features[2139]  | ~new_n12697_ | (~\all_features[2138]  & ~new_n12699_));
  assign new_n12706_ = ~\all_features[2143]  & (~\all_features[2142]  | (~\all_features[2140]  & ~\all_features[2141]  & ~new_n12701_));
  assign new_n12707_ = ~\all_features[2143]  & (~\all_features[2142]  | (~\all_features[2141]  & (new_n12694_ | ~new_n12701_ | ~\all_features[2140] )));
  assign new_n12708_ = new_n12704_ & (~\all_features[2141]  | (~\all_features[2140]  & (~\all_features[2139]  | (~\all_features[2138]  & ~\all_features[2137] ))));
  assign new_n12709_ = new_n12715_ & (~new_n12716_ | (~new_n12710_ & ~new_n12706_ & ~new_n12707_));
  assign new_n12710_ = new_n12713_ & ((~new_n12711_ & new_n12696_ & new_n12714_) | ~new_n12702_ | ~new_n12693_);
  assign new_n12711_ = \all_features[2143]  & \all_features[2142]  & ~new_n12712_ & \all_features[2141] ;
  assign new_n12712_ = ~\all_features[2139]  & ~\all_features[2140]  & (~\all_features[2138]  | new_n12694_);
  assign new_n12713_ = ~new_n12691_ & ~new_n12700_;
  assign new_n12714_ = \all_features[2142]  & \all_features[2143]  & (\all_features[2140]  | \all_features[2141]  | new_n12699_ | ~new_n12695_);
  assign new_n12715_ = ~new_n12703_ & (\all_features[2139]  | \all_features[2140]  | \all_features[2141]  | \all_features[2142]  | \all_features[2143] );
  assign new_n12716_ = ~new_n12705_ & ~new_n12708_;
  assign new_n12717_ = new_n12718_ & new_n12721_;
  assign new_n12718_ = new_n12716_ & ~new_n12719_ & new_n12715_;
  assign new_n12719_ = new_n12720_ & (~new_n12714_ | ~new_n12702_ | ~new_n12693_ | ~new_n12696_);
  assign new_n12720_ = ~new_n12700_ & ~new_n12691_ & ~new_n12706_ & ~new_n12707_;
  assign new_n12721_ = new_n12713_ & new_n12715_ & ~new_n12708_ & ~new_n12707_ & ~new_n12705_ & ~new_n12706_;
  assign new_n12722_ = new_n12723_ ? (~new_n12837_ ^ new_n13131_) : (new_n12837_ ^ new_n13131_);
  assign new_n12723_ = ~new_n12724_ & new_n12799_;
  assign new_n12724_ = ~new_n12734_ & new_n12725_ & (~new_n12757_ | (~new_n12760_ & new_n12758_) | (~new_n12792_ & ~new_n12758_));
  assign new_n12725_ = new_n12730_ | ((~new_n12726_ | ~new_n10128_) & (new_n12732_ | new_n10976_ | new_n10128_));
  assign new_n12726_ = (new_n8133_ | ~new_n12727_) & (new_n12729_ | ~new_n12187_ | new_n12727_);
  assign new_n12727_ = ~new_n10038_ & new_n12728_;
  assign new_n12728_ = ~new_n10069_ & ~new_n10060_ & ~new_n10066_;
  assign new_n12729_ = ~new_n12175_ & ~new_n12185_;
  assign new_n12730_ = ~new_n12398_ & (~new_n12376_ | new_n12731_);
  assign new_n12731_ = ~new_n12400_ & ~new_n12404_;
  assign new_n12732_ = ~new_n12733_ & new_n8923_;
  assign new_n12733_ = new_n8894_ & new_n8915_;
  assign new_n12734_ = ~new_n12755_ & new_n12735_;
  assign new_n12735_ = new_n12738_ & new_n12730_ & new_n12736_;
  assign new_n12736_ = ~new_n12030_ & new_n12737_;
  assign new_n12737_ = ~new_n12007_ & ~new_n12029_;
  assign new_n12738_ = ~new_n12338_ & (~new_n12753_ | (~new_n12747_ & ~new_n12739_));
  assign new_n12739_ = ~new_n12740_ & (\all_features[3403]  | \all_features[3404]  | \all_features[3405]  | \all_features[3406]  | \all_features[3407] );
  assign new_n12740_ = ~new_n12340_ & (new_n12351_ | (~new_n12353_ & (new_n12348_ | (~new_n12352_ & ~new_n12741_))));
  assign new_n12741_ = ~new_n12349_ & (new_n12344_ | (new_n12746_ & (~new_n12742_ | (~new_n12745_ & new_n12744_))));
  assign new_n12742_ = \all_features[3407]  & (\all_features[3406]  | (\all_features[3405]  & (\all_features[3404]  | ~new_n12743_ | ~new_n12342_)));
  assign new_n12743_ = ~\all_features[3402]  & ~\all_features[3403] ;
  assign new_n12744_ = \all_features[3407]  & (\all_features[3406]  | (new_n12347_ & (\all_features[3402]  | \all_features[3403]  | \all_features[3401] )));
  assign new_n12745_ = ~\all_features[3405]  & \all_features[3406]  & \all_features[3407]  & (\all_features[3404]  ? new_n12743_ : (new_n12346_ | ~new_n12743_));
  assign new_n12746_ = \all_features[3407]  & (\all_features[3405]  | \all_features[3406]  | \all_features[3404] );
  assign new_n12747_ = new_n12339_ & (~new_n12752_ | (~new_n12748_ & ~new_n12352_ & ~new_n12348_));
  assign new_n12748_ = ~new_n12349_ & ~new_n12344_ & (~new_n12746_ | ~new_n12742_ | new_n12749_);
  assign new_n12749_ = new_n12744_ & new_n12750_ & (new_n12751_ | ~\all_features[3405]  | ~\all_features[3406]  | ~\all_features[3407] );
  assign new_n12750_ = \all_features[3406]  & \all_features[3407]  & (\all_features[3404]  | \all_features[3405]  | new_n12346_ | ~new_n12743_);
  assign new_n12751_ = ~\all_features[3403]  & ~\all_features[3404]  & (~\all_features[3402]  | new_n12342_);
  assign new_n12752_ = ~new_n12351_ & ~new_n12353_;
  assign new_n12753_ = new_n12339_ & new_n12752_ & (new_n12754_ | new_n12349_ | new_n12352_ | ~new_n12343_);
  assign new_n12754_ = new_n12746_ & new_n12750_ & new_n12742_ & new_n12744_;
  assign new_n12755_ = ~new_n7834_ & new_n12756_;
  assign new_n12756_ = ~new_n7866_ & ~new_n7863_;
  assign new_n12757_ = ~new_n12736_ & new_n12730_;
  assign new_n12758_ = new_n7509_ & new_n12759_;
  assign new_n12759_ = ~new_n7480_ & ~new_n7501_;
  assign new_n12760_ = ~new_n12761_ & ~new_n12791_;
  assign new_n12761_ = new_n12762_ & new_n12784_;
  assign new_n12762_ = new_n12779_ & ~new_n12783_ & ~new_n12763_ & ~new_n12782_;
  assign new_n12763_ = new_n12764_ & (~new_n12777_ | ~new_n12778_ | ~new_n12774_ | ~new_n12776_);
  assign new_n12764_ = ~new_n12773_ & ~new_n12770_ & ~new_n12765_ & ~new_n12768_;
  assign new_n12765_ = ~\all_features[4343]  & (~\all_features[4342]  | (~\all_features[4341]  & (new_n12766_ | ~new_n12767_ | ~\all_features[4340] )));
  assign new_n12766_ = ~\all_features[4336]  & ~\all_features[4337] ;
  assign new_n12767_ = \all_features[4338]  & \all_features[4339] ;
  assign new_n12768_ = ~new_n12769_ & ~\all_features[4343] ;
  assign new_n12769_ = \all_features[4341]  & \all_features[4342]  & (\all_features[4340]  | (\all_features[4338]  & \all_features[4339]  & \all_features[4337] ));
  assign new_n12770_ = ~\all_features[4343]  & (~\all_features[4342]  | ~new_n12771_ | ~new_n12772_ | ~new_n12767_);
  assign new_n12771_ = \all_features[4340]  & \all_features[4341] ;
  assign new_n12772_ = \all_features[4336]  & \all_features[4337] ;
  assign new_n12773_ = ~\all_features[4343]  & (~\all_features[4342]  | (~\all_features[4340]  & ~\all_features[4341]  & ~new_n12767_));
  assign new_n12774_ = \all_features[4343]  & (\all_features[4342]  | (\all_features[4341]  & (\all_features[4340]  | ~new_n12766_ | ~new_n12775_)));
  assign new_n12775_ = ~\all_features[4338]  & ~\all_features[4339] ;
  assign new_n12776_ = \all_features[4343]  & (\all_features[4342]  | (new_n12771_ & (\all_features[4338]  | \all_features[4339]  | \all_features[4337] )));
  assign new_n12777_ = \all_features[4342]  & \all_features[4343]  & (\all_features[4340]  | \all_features[4341]  | new_n12772_ | ~new_n12775_);
  assign new_n12778_ = \all_features[4343]  & (\all_features[4341]  | \all_features[4342]  | \all_features[4340] );
  assign new_n12779_ = ~new_n12780_ & (\all_features[4339]  | \all_features[4340]  | \all_features[4341]  | \all_features[4342]  | \all_features[4343] );
  assign new_n12780_ = ~\all_features[4341]  & new_n12781_ & ((~\all_features[4338]  & new_n12766_) | ~\all_features[4340]  | ~\all_features[4339] );
  assign new_n12781_ = ~\all_features[4342]  & ~\all_features[4343] ;
  assign new_n12782_ = new_n12781_ & (~\all_features[4341]  | (~\all_features[4340]  & (~\all_features[4339]  | (~\all_features[4338]  & ~\all_features[4337] ))));
  assign new_n12783_ = new_n12781_ & (~\all_features[4339]  | ~new_n12771_ | (~\all_features[4338]  & ~new_n12772_));
  assign new_n12784_ = new_n12779_ & (~new_n12790_ | (~new_n12785_ & new_n12789_));
  assign new_n12785_ = new_n12788_ & ((~new_n12786_ & new_n12776_ & new_n12777_) | ~new_n12778_ | ~new_n12774_);
  assign new_n12786_ = \all_features[4343]  & \all_features[4342]  & ~new_n12787_ & \all_features[4341] ;
  assign new_n12787_ = ~\all_features[4339]  & ~\all_features[4340]  & (~\all_features[4338]  | new_n12766_);
  assign new_n12788_ = ~new_n12768_ & ~new_n12770_;
  assign new_n12789_ = ~new_n12765_ & ~new_n12773_;
  assign new_n12790_ = ~new_n12782_ & ~new_n12783_;
  assign new_n12791_ = new_n12790_ & new_n12789_ & new_n12779_ & new_n12788_;
  assign new_n12792_ = new_n12793_ & new_n12798_;
  assign new_n12793_ = new_n12229_ & new_n12794_;
  assign new_n12794_ = ~new_n12795_ & (\all_features[3011]  | \all_features[3012]  | \all_features[3013]  | \all_features[3014]  | \all_features[3015] );
  assign new_n12795_ = ~new_n12251_ & (new_n12247_ | (~new_n12245_ & (new_n12252_ | (~new_n12248_ & ~new_n12796_))));
  assign new_n12796_ = ~new_n12241_ & (new_n12240_ | (new_n12243_ & (~new_n12239_ | (~new_n12797_ & new_n12232_))));
  assign new_n12797_ = ~\all_features[3013]  & \all_features[3014]  & \all_features[3015]  & (\all_features[3012]  ? new_n12236_ : (new_n12235_ | ~new_n12236_));
  assign new_n12798_ = new_n12254_ & new_n12257_;
  assign new_n12799_ = new_n12800_ & (~new_n12735_ | ~new_n12755_) & (new_n12758_ | new_n12792_ | ~new_n12757_);
  assign new_n12800_ = (new_n12730_ | (new_n10128_ ? new_n12726_ : ~new_n12801_)) & (~new_n12836_ | ~new_n12736_ | ~new_n12730_);
  assign new_n12801_ = new_n10976_ ? new_n12802_ : new_n12732_;
  assign new_n12802_ = new_n12834_ & (new_n12825_ | new_n12829_ | new_n12803_);
  assign new_n12803_ = ~new_n12804_ & ~new_n12824_;
  assign new_n12804_ = ~new_n12819_ & (new_n12821_ | (~new_n12822_ & (new_n12823_ | (~new_n12805_ & ~new_n12808_))));
  assign new_n12805_ = ~\all_features[4231]  & (~\all_features[4230]  | new_n12806_);
  assign new_n12806_ = ~\all_features[4229]  & (new_n12807_ | ~\all_features[4227]  | ~\all_features[4228]  | ~\all_features[4226] );
  assign new_n12807_ = ~\all_features[4224]  & ~\all_features[4225] ;
  assign new_n12808_ = ~new_n12809_ & (new_n12811_ | (new_n12818_ & (~new_n12814_ | (~new_n12817_ & new_n12816_))));
  assign new_n12809_ = ~new_n12810_ & ~\all_features[4231] ;
  assign new_n12810_ = \all_features[4229]  & \all_features[4230]  & (\all_features[4228]  | (\all_features[4226]  & \all_features[4227]  & \all_features[4225] ));
  assign new_n12811_ = ~\all_features[4231]  & (~new_n12813_ | ~\all_features[4226]  | ~\all_features[4227]  | ~\all_features[4230]  | ~new_n12812_);
  assign new_n12812_ = \all_features[4224]  & \all_features[4225] ;
  assign new_n12813_ = \all_features[4228]  & \all_features[4229] ;
  assign new_n12814_ = \all_features[4231]  & (\all_features[4230]  | (\all_features[4229]  & (\all_features[4228]  | ~new_n12815_ | ~new_n12807_)));
  assign new_n12815_ = ~\all_features[4226]  & ~\all_features[4227] ;
  assign new_n12816_ = \all_features[4231]  & (\all_features[4230]  | (new_n12813_ & (\all_features[4226]  | \all_features[4227]  | \all_features[4225] )));
  assign new_n12817_ = ~\all_features[4229]  & \all_features[4230]  & \all_features[4231]  & (\all_features[4228]  ? new_n12815_ : (new_n12812_ | ~new_n12815_));
  assign new_n12818_ = \all_features[4231]  & (\all_features[4229]  | \all_features[4230]  | \all_features[4228] );
  assign new_n12819_ = ~\all_features[4229]  & new_n12820_ & ((~\all_features[4226]  & new_n12807_) | ~\all_features[4228]  | ~\all_features[4227] );
  assign new_n12820_ = ~\all_features[4230]  & ~\all_features[4231] ;
  assign new_n12821_ = new_n12820_ & (~\all_features[4229]  | (~\all_features[4228]  & (~\all_features[4227]  | (~\all_features[4226]  & ~\all_features[4225] ))));
  assign new_n12822_ = new_n12820_ & (~\all_features[4227]  | ~new_n12813_ | (~\all_features[4226]  & ~new_n12812_));
  assign new_n12823_ = ~\all_features[4231]  & (~\all_features[4230]  | (~\all_features[4229]  & ~\all_features[4228]  & (~\all_features[4227]  | ~\all_features[4226] )));
  assign new_n12824_ = ~\all_features[4231]  & ~\all_features[4230]  & ~\all_features[4229]  & ~\all_features[4227]  & ~\all_features[4228] ;
  assign new_n12825_ = ~new_n12824_ & ~new_n12822_ & ~new_n12821_ & ~new_n12826_ & ~new_n12819_;
  assign new_n12826_ = ~new_n12823_ & ~new_n12811_ & ~new_n12809_ & ~new_n12805_ & ~new_n12827_;
  assign new_n12827_ = new_n12818_ & new_n12828_ & new_n12814_ & new_n12816_;
  assign new_n12828_ = \all_features[4230]  & \all_features[4231]  & (\all_features[4228]  | \all_features[4229]  | new_n12812_ | ~new_n12815_);
  assign new_n12829_ = ~new_n12824_ & ~new_n12819_ & (~new_n12833_ | (~new_n12830_ & ~new_n12805_ & ~new_n12823_));
  assign new_n12830_ = ~new_n12809_ & ~new_n12811_ & (~new_n12818_ | ~new_n12814_ | new_n12831_);
  assign new_n12831_ = new_n12816_ & new_n12828_ & (new_n12832_ | ~\all_features[4229]  | ~\all_features[4230]  | ~\all_features[4231] );
  assign new_n12832_ = ~\all_features[4227]  & ~\all_features[4228]  & (~\all_features[4226]  | new_n12807_);
  assign new_n12833_ = ~new_n12821_ & ~new_n12822_;
  assign new_n12834_ = new_n12833_ & new_n12835_ & ~new_n12823_ & ~new_n12819_ & ~new_n12805_ & ~new_n12809_;
  assign new_n12835_ = ~new_n12811_ & ~new_n12824_;
  assign new_n12836_ = ~new_n11095_ & ~new_n12738_;
  assign new_n12837_ = new_n12838_ ? (new_n12867_ ^ new_n13060_) : (~new_n12867_ ^ new_n13060_);
  assign new_n12838_ = new_n12859_ & (~new_n8484_ | (new_n8356_ & new_n10875_ & ~new_n12866_) | (new_n12839_ & new_n12866_));
  assign new_n12839_ = new_n12840_ ? new_n12849_ : (new_n11573_ | (~new_n12850_ & new_n11551_));
  assign new_n12840_ = new_n12841_ & (new_n9481_ | (~new_n12846_ & ~new_n9479_));
  assign new_n12841_ = ~new_n12842_ & new_n9459_;
  assign new_n12842_ = ~new_n9479_ & ~new_n9481_ & (~new_n9484_ | (~new_n12843_ & ~new_n9466_ & ~new_n9470_));
  assign new_n12843_ = ~new_n9471_ & ~new_n9468_ & (~new_n9476_ | new_n12844_ | ~new_n9462_);
  assign new_n12844_ = ~new_n9475_ & new_n9473_ & \all_features[1214]  & \all_features[1215]  & (~\all_features[1213]  | new_n12845_);
  assign new_n12845_ = ~\all_features[1211]  & ~\all_features[1212]  & (~\all_features[1210]  | new_n9464_);
  assign new_n12846_ = ~new_n9477_ & (new_n9480_ | (~new_n9470_ & (new_n9466_ | (~new_n9468_ & ~new_n12847_))));
  assign new_n12847_ = ~new_n9471_ & (~new_n9476_ | (new_n9462_ & (~new_n9473_ | (~new_n12848_ & new_n9474_))));
  assign new_n12848_ = \all_features[1214]  & \all_features[1215]  & (\all_features[1213]  | (\all_features[1212]  & (\all_features[1211]  | \all_features[1210] )));
  assign new_n12849_ = new_n11304_ & new_n12266_;
  assign new_n12850_ = ~new_n12851_ & ~new_n12855_;
  assign new_n12851_ = new_n11553_ & (new_n11558_ | new_n11557_ | (~new_n11562_ & ~new_n11567_ & ~new_n12852_));
  assign new_n12852_ = ~new_n11566_ & ~new_n11564_ & (~new_n11572_ | ~new_n11568_ | new_n12853_);
  assign new_n12853_ = new_n11570_ & new_n11571_ & (new_n12854_ | ~\all_features[2965]  | ~\all_features[2966]  | ~\all_features[2967] );
  assign new_n12854_ = ~\all_features[2963]  & ~\all_features[2964]  & (~\all_features[2962]  | new_n11555_);
  assign new_n12855_ = ~new_n12856_ & (\all_features[2963]  | \all_features[2964]  | \all_features[2965]  | \all_features[2966]  | \all_features[2967] );
  assign new_n12856_ = ~new_n11554_ & (new_n11557_ | (~new_n11558_ & (new_n11567_ | (~new_n11562_ & ~new_n12857_))));
  assign new_n12857_ = ~new_n11564_ & (new_n11566_ | (new_n11572_ & (~new_n11568_ | (~new_n12858_ & new_n11570_))));
  assign new_n12858_ = ~\all_features[2965]  & \all_features[2966]  & \all_features[2967]  & (\all_features[2964]  ? new_n11569_ : (new_n11560_ | ~new_n11569_));
  assign new_n12859_ = ~new_n12860_ & (new_n8484_ | (~new_n12863_ & new_n12861_) | (~new_n12864_ & ~new_n12375_ & ~new_n12861_));
  assign new_n12860_ = ~new_n8484_ & new_n7227_ & new_n12861_ & (~new_n8854_ | (~new_n8851_ & new_n8819_));
  assign new_n12861_ = ~new_n11407_ & (~new_n11409_ | ~new_n11379_);
  assign new_n12863_ = new_n9058_ & new_n9055_ & ~new_n7227_ & new_n9045_;
  assign new_n12864_ = ~new_n11940_ & new_n12865_;
  assign new_n12865_ = ~new_n11908_ & ~new_n11931_;
  assign new_n12866_ = ~new_n12187_ & (~new_n12185_ | ~new_n12154_);
  assign new_n12867_ = ~new_n12944_ & new_n12981_ & (new_n9129_ ? (new_n13014_ | new_n12945_) : new_n12868_);
  assign new_n12868_ = (new_n12869_ | ~new_n12907_) & (~new_n9547_ | ~new_n12908_ | new_n12907_);
  assign new_n12869_ = (new_n12560_ | ~new_n12870_) & (new_n10646_ | ~new_n12906_ | new_n12870_);
  assign new_n12870_ = ~new_n12871_ & new_n12900_;
  assign new_n12871_ = new_n12872_ & new_n12896_;
  assign new_n12872_ = new_n12887_ & (~new_n12892_ | (~new_n12890_ & ~new_n12873_ & ~new_n12895_));
  assign new_n12873_ = ~new_n12885_ & ~new_n12883_ & (~new_n12886_ | ~new_n12882_ | new_n12874_);
  assign new_n12874_ = new_n12875_ & new_n12877_ & (new_n12880_ | ~\all_features[3517]  | ~\all_features[3518]  | ~\all_features[3519] );
  assign new_n12875_ = \all_features[3519]  & (\all_features[3518]  | (new_n12876_ & (\all_features[3514]  | \all_features[3515]  | \all_features[3513] )));
  assign new_n12876_ = \all_features[3516]  & \all_features[3517] ;
  assign new_n12877_ = \all_features[3518]  & \all_features[3519]  & (\all_features[3516]  | \all_features[3517]  | new_n12879_ | ~new_n12878_);
  assign new_n12878_ = ~\all_features[3514]  & ~\all_features[3515] ;
  assign new_n12879_ = \all_features[3512]  & \all_features[3513] ;
  assign new_n12880_ = ~\all_features[3515]  & ~\all_features[3516]  & (~\all_features[3514]  | new_n12881_);
  assign new_n12881_ = ~\all_features[3512]  & ~\all_features[3513] ;
  assign new_n12882_ = \all_features[3519]  & (\all_features[3518]  | (\all_features[3517]  & (\all_features[3516]  | ~new_n12878_ | ~new_n12881_)));
  assign new_n12883_ = ~new_n12884_ & ~\all_features[3519] ;
  assign new_n12884_ = \all_features[3517]  & \all_features[3518]  & (\all_features[3516]  | (\all_features[3514]  & \all_features[3515]  & \all_features[3513] ));
  assign new_n12885_ = ~\all_features[3519]  & (~new_n12879_ | ~\all_features[3514]  | ~\all_features[3515]  | ~\all_features[3518]  | ~new_n12876_);
  assign new_n12886_ = \all_features[3519]  & (\all_features[3517]  | \all_features[3518]  | \all_features[3516] );
  assign new_n12887_ = ~new_n12888_ & (\all_features[3515]  | \all_features[3516]  | \all_features[3517]  | \all_features[3518]  | \all_features[3519] );
  assign new_n12888_ = ~\all_features[3517]  & new_n12889_ & ((~\all_features[3514]  & new_n12881_) | ~\all_features[3516]  | ~\all_features[3515] );
  assign new_n12889_ = ~\all_features[3518]  & ~\all_features[3519] ;
  assign new_n12890_ = ~\all_features[3519]  & (~\all_features[3518]  | new_n12891_);
  assign new_n12891_ = ~\all_features[3517]  & (new_n12881_ | ~\all_features[3515]  | ~\all_features[3516]  | ~\all_features[3514] );
  assign new_n12892_ = ~new_n12893_ & ~new_n12894_;
  assign new_n12893_ = new_n12889_ & (~\all_features[3517]  | (~\all_features[3516]  & (~\all_features[3515]  | (~\all_features[3514]  & ~\all_features[3513] ))));
  assign new_n12894_ = new_n12889_ & (~\all_features[3515]  | ~new_n12876_ | (~new_n12879_ & ~\all_features[3514] ));
  assign new_n12895_ = ~\all_features[3519]  & (~\all_features[3518]  | (~\all_features[3517]  & ~\all_features[3516]  & (~\all_features[3515]  | ~\all_features[3514] )));
  assign new_n12896_ = ~new_n12897_ & (\all_features[3515]  | \all_features[3516]  | \all_features[3517]  | \all_features[3518]  | \all_features[3519] );
  assign new_n12897_ = ~new_n12888_ & (new_n12893_ | (~new_n12894_ & (new_n12895_ | (~new_n12890_ & ~new_n12898_))));
  assign new_n12898_ = ~new_n12883_ & (new_n12885_ | (new_n12886_ & (~new_n12882_ | (~new_n12899_ & new_n12875_))));
  assign new_n12899_ = ~\all_features[3517]  & \all_features[3518]  & \all_features[3519]  & (\all_features[3516]  ? new_n12878_ : (new_n12879_ | ~new_n12878_));
  assign new_n12900_ = ~new_n12901_ & ~new_n12904_;
  assign new_n12901_ = new_n12892_ & ~new_n12902_ & new_n12887_;
  assign new_n12902_ = ~new_n12895_ & ~new_n12885_ & ~new_n12883_ & ~new_n12890_ & ~new_n12903_;
  assign new_n12903_ = new_n12886_ & new_n12882_ & new_n12875_ & new_n12877_;
  assign new_n12904_ = new_n12887_ & new_n12905_ & ~new_n12883_ & ~new_n12893_;
  assign new_n12905_ = ~new_n12895_ & ~new_n12894_ & ~new_n12890_ & ~new_n12885_;
  assign new_n12906_ = new_n9721_ & new_n9724_;
  assign new_n12907_ = new_n6953_ & (new_n6950_ | ~new_n6920_);
  assign new_n12908_ = new_n12909_ & new_n12935_;
  assign new_n12909_ = ~new_n12910_ & ~new_n12933_;
  assign new_n12910_ = new_n12928_ & ~new_n12932_ & ~new_n12911_ & ~new_n12931_;
  assign new_n12911_ = ~new_n12926_ & ~new_n12927_ & new_n12919_ & (~new_n12924_ | ~new_n12912_);
  assign new_n12912_ = new_n12918_ & new_n12913_ & new_n12915_;
  assign new_n12913_ = \all_features[3255]  & (\all_features[3254]  | (new_n12914_ & (\all_features[3250]  | \all_features[3251]  | \all_features[3249] )));
  assign new_n12914_ = \all_features[3252]  & \all_features[3253] ;
  assign new_n12915_ = \all_features[3254]  & \all_features[3255]  & (\all_features[3252]  | \all_features[3253]  | new_n12917_ | ~new_n12916_);
  assign new_n12916_ = ~\all_features[3250]  & ~\all_features[3251] ;
  assign new_n12917_ = \all_features[3248]  & \all_features[3249] ;
  assign new_n12918_ = \all_features[3255]  & (\all_features[3253]  | \all_features[3254]  | \all_features[3252] );
  assign new_n12919_ = ~new_n12920_ & ~new_n12922_;
  assign new_n12920_ = ~new_n12921_ & ~\all_features[3255] ;
  assign new_n12921_ = \all_features[3253]  & \all_features[3254]  & (\all_features[3252]  | (\all_features[3250]  & \all_features[3251]  & \all_features[3249] ));
  assign new_n12922_ = ~\all_features[3255]  & (~\all_features[3254]  | (~\all_features[3252]  & ~\all_features[3253]  & ~new_n12923_));
  assign new_n12923_ = \all_features[3250]  & \all_features[3251] ;
  assign new_n12924_ = \all_features[3255]  & (\all_features[3254]  | (\all_features[3253]  & (\all_features[3252]  | ~new_n12925_ | ~new_n12916_)));
  assign new_n12925_ = ~\all_features[3248]  & ~\all_features[3249] ;
  assign new_n12926_ = ~\all_features[3255]  & (~\all_features[3254]  | (~\all_features[3253]  & (new_n12925_ | ~new_n12923_ | ~\all_features[3252] )));
  assign new_n12927_ = ~\all_features[3255]  & (~\all_features[3254]  | ~new_n12914_ | ~new_n12917_ | ~new_n12923_);
  assign new_n12928_ = ~new_n12929_ & (\all_features[3251]  | \all_features[3252]  | \all_features[3253]  | \all_features[3254]  | \all_features[3255] );
  assign new_n12929_ = ~\all_features[3253]  & new_n12930_ & ((~\all_features[3250]  & new_n12925_) | ~\all_features[3252]  | ~\all_features[3251] );
  assign new_n12930_ = ~\all_features[3254]  & ~\all_features[3255] ;
  assign new_n12931_ = new_n12930_ & (~\all_features[3253]  | (~\all_features[3252]  & (~\all_features[3251]  | (~\all_features[3250]  & ~\all_features[3249] ))));
  assign new_n12932_ = new_n12930_ & (~\all_features[3251]  | ~new_n12914_ | (~\all_features[3250]  & ~new_n12917_));
  assign new_n12933_ = new_n12928_ & new_n12919_ & new_n12934_ & ~new_n12926_ & ~new_n12927_;
  assign new_n12934_ = ~new_n12931_ & ~new_n12932_;
  assign new_n12935_ = ~new_n12936_ & ~new_n12940_;
  assign new_n12936_ = new_n12928_ & (~new_n12934_ | (~new_n12937_ & ~new_n12922_ & ~new_n12926_));
  assign new_n12937_ = ~new_n12927_ & ~new_n12920_ & (~new_n12918_ | ~new_n12924_ | new_n12938_);
  assign new_n12938_ = new_n12913_ & new_n12915_ & (new_n12939_ | ~\all_features[3253]  | ~\all_features[3254]  | ~\all_features[3255] );
  assign new_n12939_ = ~\all_features[3251]  & ~\all_features[3252]  & (~\all_features[3250]  | new_n12925_);
  assign new_n12940_ = ~new_n12941_ & (\all_features[3251]  | \all_features[3252]  | \all_features[3253]  | \all_features[3254]  | \all_features[3255] );
  assign new_n12941_ = ~new_n12929_ & (new_n12931_ | (~new_n12932_ & (new_n12922_ | (~new_n12926_ & ~new_n12942_))));
  assign new_n12942_ = ~new_n12920_ & (new_n12927_ | (new_n12918_ & (~new_n12924_ | (~new_n12943_ & new_n12913_))));
  assign new_n12943_ = ~\all_features[3253]  & \all_features[3254]  & \all_features[3255]  & (\all_features[3252]  ? new_n12916_ : (new_n12917_ | ~new_n12916_));
  assign new_n12944_ = ~new_n12907_ & ~new_n9547_ & ~new_n9129_ & (new_n7866_ | new_n7833_);
  assign new_n12945_ = new_n7407_ & new_n9760_ & new_n12946_;
  assign new_n12946_ = new_n12977_ & new_n12947_ & new_n12968_;
  assign new_n12947_ = ~new_n12948_ & (\all_features[4595]  | \all_features[4596]  | \all_features[4597]  | \all_features[4598]  | \all_features[4599] );
  assign new_n12948_ = ~new_n12962_ & (new_n12964_ | (~new_n12965_ & (new_n12966_ | (~new_n12949_ & ~new_n12967_))));
  assign new_n12949_ = ~new_n12950_ & (new_n12952_ | (new_n12961_ & (~new_n12956_ | (~new_n12960_ & new_n12959_))));
  assign new_n12950_ = ~new_n12951_ & ~\all_features[4599] ;
  assign new_n12951_ = \all_features[4597]  & \all_features[4598]  & (\all_features[4596]  | (\all_features[4594]  & \all_features[4595]  & \all_features[4593] ));
  assign new_n12952_ = ~\all_features[4599]  & (~\all_features[4598]  | ~new_n12953_ | ~new_n12954_ | ~new_n12955_);
  assign new_n12953_ = \all_features[4592]  & \all_features[4593] ;
  assign new_n12954_ = \all_features[4596]  & \all_features[4597] ;
  assign new_n12955_ = \all_features[4594]  & \all_features[4595] ;
  assign new_n12956_ = \all_features[4599]  & (\all_features[4598]  | (\all_features[4597]  & (\all_features[4596]  | ~new_n12958_ | ~new_n12957_)));
  assign new_n12957_ = ~\all_features[4592]  & ~\all_features[4593] ;
  assign new_n12958_ = ~\all_features[4594]  & ~\all_features[4595] ;
  assign new_n12959_ = \all_features[4599]  & (\all_features[4598]  | (new_n12954_ & (\all_features[4594]  | \all_features[4595]  | \all_features[4593] )));
  assign new_n12960_ = ~\all_features[4597]  & \all_features[4598]  & \all_features[4599]  & (\all_features[4596]  ? new_n12958_ : (new_n12953_ | ~new_n12958_));
  assign new_n12961_ = \all_features[4599]  & (\all_features[4597]  | \all_features[4598]  | \all_features[4596] );
  assign new_n12962_ = ~\all_features[4597]  & new_n12963_ & ((~\all_features[4594]  & new_n12957_) | ~\all_features[4596]  | ~\all_features[4595] );
  assign new_n12963_ = ~\all_features[4598]  & ~\all_features[4599] ;
  assign new_n12964_ = new_n12963_ & (~\all_features[4597]  | (~\all_features[4596]  & (~\all_features[4595]  | (~\all_features[4594]  & ~\all_features[4593] ))));
  assign new_n12965_ = new_n12963_ & (~\all_features[4595]  | ~new_n12954_ | (~\all_features[4594]  & ~new_n12953_));
  assign new_n12966_ = ~\all_features[4599]  & (~\all_features[4598]  | (~\all_features[4596]  & ~\all_features[4597]  & ~new_n12955_));
  assign new_n12967_ = ~\all_features[4599]  & (~\all_features[4598]  | (~\all_features[4597]  & (new_n12957_ | ~new_n12955_ | ~\all_features[4596] )));
  assign new_n12968_ = new_n12976_ & (~new_n12974_ | (~new_n12969_ & new_n12975_));
  assign new_n12969_ = new_n12972_ & ((~new_n12970_ & new_n12959_ & new_n12973_) | ~new_n12961_ | ~new_n12956_);
  assign new_n12970_ = \all_features[4599]  & \all_features[4598]  & ~new_n12971_ & \all_features[4597] ;
  assign new_n12971_ = ~\all_features[4595]  & ~\all_features[4596]  & (~\all_features[4594]  | new_n12957_);
  assign new_n12972_ = ~new_n12950_ & ~new_n12952_;
  assign new_n12973_ = \all_features[4598]  & \all_features[4599]  & (\all_features[4596]  | \all_features[4597]  | new_n12953_ | ~new_n12958_);
  assign new_n12974_ = ~new_n12964_ & ~new_n12965_;
  assign new_n12975_ = ~new_n12966_ & ~new_n12967_;
  assign new_n12976_ = ~new_n12962_ & (\all_features[4595]  | \all_features[4596]  | \all_features[4597]  | \all_features[4598]  | \all_features[4599] );
  assign new_n12977_ = new_n12978_ & new_n12980_;
  assign new_n12978_ = new_n12974_ & new_n12976_ & (~new_n12972_ | ~new_n12975_ | (new_n12979_ & new_n12956_));
  assign new_n12979_ = new_n12961_ & new_n12959_ & new_n12973_;
  assign new_n12980_ = new_n12976_ & new_n12974_ & ~new_n12952_ & ~new_n12950_ & ~new_n12966_ & ~new_n12967_;
  assign new_n12981_ = ~new_n13013_ | ((new_n10438_ | new_n12982_ | (new_n13057_ & new_n13040_)) & (new_n9689_ | ~new_n12982_));
  assign new_n12982_ = ~new_n12983_ & new_n13012_;
  assign new_n12983_ = ~new_n12984_ & ~new_n13009_;
  assign new_n12984_ = new_n13007_ & (~new_n12995_ | (new_n12999_ & (~new_n13003_ | new_n12985_)));
  assign new_n12985_ = new_n12986_ & (~new_n12989_ | (~new_n12994_ & \all_features[1453]  & \all_features[1454]  & \all_features[1455] ));
  assign new_n12986_ = \all_features[1455]  & (\all_features[1454]  | (~new_n12987_ & \all_features[1453] ));
  assign new_n12987_ = new_n12988_ & ~\all_features[1452]  & ~\all_features[1450]  & ~\all_features[1451] ;
  assign new_n12988_ = ~\all_features[1448]  & ~\all_features[1449] ;
  assign new_n12989_ = \all_features[1455]  & \all_features[1454]  & ~new_n12992_ & new_n12990_;
  assign new_n12990_ = \all_features[1455]  & (\all_features[1454]  | (new_n12991_ & (\all_features[1450]  | \all_features[1451]  | \all_features[1449] )));
  assign new_n12991_ = \all_features[1452]  & \all_features[1453] ;
  assign new_n12992_ = ~\all_features[1453]  & ~\all_features[1452]  & ~\all_features[1451]  & ~new_n12993_ & ~\all_features[1450] ;
  assign new_n12993_ = \all_features[1448]  & \all_features[1449] ;
  assign new_n12994_ = ~\all_features[1451]  & ~\all_features[1452]  & (~\all_features[1450]  | new_n12988_);
  assign new_n12995_ = ~new_n12996_ & ~new_n12997_;
  assign new_n12996_ = ~\all_features[1454]  & ~\all_features[1455]  & (~\all_features[1451]  | ~new_n12991_ | (~\all_features[1450]  & ~new_n12993_));
  assign new_n12997_ = ~\all_features[1455]  & ~new_n12998_ & ~\all_features[1454] ;
  assign new_n12998_ = \all_features[1453]  & (\all_features[1452]  | (\all_features[1451]  & (\all_features[1450]  | \all_features[1449] )));
  assign new_n12999_ = ~new_n13000_ & ~new_n13002_;
  assign new_n13000_ = ~\all_features[1455]  & (~\all_features[1454]  | (~\all_features[1452]  & ~\all_features[1453]  & ~new_n13001_));
  assign new_n13001_ = \all_features[1450]  & \all_features[1451] ;
  assign new_n13002_ = ~\all_features[1455]  & (~\all_features[1454]  | (~\all_features[1453]  & (new_n12988_ | ~new_n13001_ | ~\all_features[1452] )));
  assign new_n13003_ = ~new_n13004_ & ~new_n13005_;
  assign new_n13004_ = ~\all_features[1455]  & (~\all_features[1454]  | ~new_n12993_ | ~new_n12991_ | ~new_n13001_);
  assign new_n13005_ = ~new_n13006_ & ~\all_features[1455] ;
  assign new_n13006_ = \all_features[1453]  & \all_features[1454]  & (\all_features[1452]  | (\all_features[1450]  & \all_features[1451]  & \all_features[1449] ));
  assign new_n13007_ = ~new_n13008_ | (\all_features[1451]  & \all_features[1452]  & (\all_features[1450]  | ~new_n12988_));
  assign new_n13008_ = ~\all_features[1455]  & ~\all_features[1453]  & ~\all_features[1454] ;
  assign new_n13009_ = new_n13010_ & (new_n13002_ | new_n13005_ | ~new_n13011_ | (new_n12989_ & new_n12986_));
  assign new_n13010_ = new_n12995_ & new_n13007_;
  assign new_n13011_ = ~new_n13000_ & ~new_n13004_;
  assign new_n13012_ = new_n13003_ & new_n13010_ & new_n12999_;
  assign new_n13013_ = new_n13014_ & new_n9129_;
  assign new_n13014_ = new_n13015_ & new_n13038_;
  assign new_n13015_ = new_n13033_ & ~new_n13037_ & ~new_n13016_ & ~new_n13036_;
  assign new_n13016_ = ~new_n13031_ & ~new_n13032_ & new_n13024_ & (~new_n13029_ | ~new_n13017_);
  assign new_n13017_ = new_n13023_ & new_n13018_ & new_n13020_;
  assign new_n13018_ = \all_features[2607]  & (\all_features[2606]  | (new_n13019_ & (\all_features[2602]  | \all_features[2603]  | \all_features[2601] )));
  assign new_n13019_ = \all_features[2604]  & \all_features[2605] ;
  assign new_n13020_ = \all_features[2606]  & \all_features[2607]  & (\all_features[2604]  | \all_features[2605]  | new_n13022_ | ~new_n13021_);
  assign new_n13021_ = ~\all_features[2602]  & ~\all_features[2603] ;
  assign new_n13022_ = \all_features[2600]  & \all_features[2601] ;
  assign new_n13023_ = \all_features[2607]  & (\all_features[2605]  | \all_features[2606]  | \all_features[2604] );
  assign new_n13024_ = ~new_n13025_ & ~new_n13027_;
  assign new_n13025_ = ~new_n13026_ & ~\all_features[2607] ;
  assign new_n13026_ = \all_features[2605]  & \all_features[2606]  & (\all_features[2604]  | (\all_features[2602]  & \all_features[2603]  & \all_features[2601] ));
  assign new_n13027_ = ~\all_features[2607]  & (~\all_features[2606]  | (~\all_features[2604]  & ~\all_features[2605]  & ~new_n13028_));
  assign new_n13028_ = \all_features[2602]  & \all_features[2603] ;
  assign new_n13029_ = \all_features[2607]  & (\all_features[2606]  | (\all_features[2605]  & (\all_features[2604]  | ~new_n13030_ | ~new_n13021_)));
  assign new_n13030_ = ~\all_features[2600]  & ~\all_features[2601] ;
  assign new_n13031_ = ~\all_features[2607]  & (~\all_features[2606]  | (~\all_features[2605]  & (new_n13030_ | ~new_n13028_ | ~\all_features[2604] )));
  assign new_n13032_ = ~\all_features[2607]  & (~\all_features[2606]  | ~new_n13019_ | ~new_n13022_ | ~new_n13028_);
  assign new_n13033_ = ~new_n13034_ & (\all_features[2603]  | \all_features[2604]  | \all_features[2605]  | \all_features[2606]  | \all_features[2607] );
  assign new_n13034_ = ~\all_features[2605]  & new_n13035_ & ((~\all_features[2602]  & new_n13030_) | ~\all_features[2604]  | ~\all_features[2603] );
  assign new_n13035_ = ~\all_features[2606]  & ~\all_features[2607] ;
  assign new_n13036_ = new_n13035_ & (~\all_features[2605]  | (~\all_features[2604]  & (~\all_features[2603]  | (~\all_features[2602]  & ~\all_features[2601] ))));
  assign new_n13037_ = new_n13035_ & (~\all_features[2603]  | ~new_n13019_ | (~\all_features[2602]  & ~new_n13022_));
  assign new_n13038_ = new_n13033_ & new_n13024_ & new_n13039_ & ~new_n13031_ & ~new_n13032_;
  assign new_n13039_ = ~new_n13036_ & ~new_n13037_;
  assign new_n13040_ = new_n13041_ & new_n13055_;
  assign new_n13041_ = new_n13053_ & (~new_n13054_ | (new_n13051_ & (~new_n13052_ | new_n13042_)));
  assign new_n13042_ = new_n13050_ & ~new_n13043_ & new_n13049_;
  assign new_n13043_ = new_n13045_ & new_n13044_ & (~\all_features[4797]  | ~new_n13047_ | new_n13048_);
  assign new_n13044_ = \all_features[4799]  & (\all_features[4798]  | (new_n10446_ & (\all_features[4794]  | \all_features[4795]  | \all_features[4793] )));
  assign new_n13045_ = new_n13047_ & (new_n10445_ | \all_features[4796]  | \all_features[4797]  | ~new_n13046_);
  assign new_n13046_ = ~\all_features[4794]  & ~\all_features[4795] ;
  assign new_n13047_ = \all_features[4798]  & \all_features[4799] ;
  assign new_n13048_ = ~\all_features[4795]  & ~\all_features[4796]  & (~\all_features[4794]  | new_n10450_);
  assign new_n13049_ = \all_features[4799]  & (\all_features[4798]  | (\all_features[4797]  & (\all_features[4796]  | ~new_n13046_ | ~new_n10450_)));
  assign new_n13050_ = \all_features[4799]  & (\all_features[4797]  | \all_features[4798]  | \all_features[4796] );
  assign new_n13051_ = ~new_n10449_ & ~new_n10451_;
  assign new_n13052_ = ~new_n10440_ & ~new_n10444_;
  assign new_n13053_ = ~new_n10452_ & ~new_n10448_;
  assign new_n13054_ = ~new_n10442_ & ~new_n10453_;
  assign new_n13055_ = new_n13054_ & new_n13053_ & (~new_n13052_ | ~new_n13051_ | (new_n13056_ & new_n13049_));
  assign new_n13056_ = new_n13050_ & new_n13044_ & new_n13045_;
  assign new_n13057_ = ~new_n10448_ & (new_n10452_ | (~new_n10442_ & (new_n10453_ | (~new_n10451_ & ~new_n13058_))));
  assign new_n13058_ = ~new_n10449_ & (new_n10440_ | (~new_n10444_ & (~new_n13050_ | (~new_n13059_ & new_n13049_))));
  assign new_n13059_ = new_n13044_ & (\all_features[4797]  | ~new_n13047_ | (~new_n10445_ & ~\all_features[4796]  & new_n13046_) | (\all_features[4796]  & ~new_n13046_));
  assign new_n13060_ = ~new_n13096_ & new_n13061_ & (~new_n13130_ | new_n13099_);
  assign new_n13061_ = (~new_n13065_ | new_n13064_ | ~new_n11635_) & (new_n13062_ | ~new_n13063_ | ~new_n9724_ | new_n11635_);
  assign new_n13062_ = ~new_n9690_ & ~new_n9721_;
  assign new_n13063_ = ~new_n6630_ & new_n6604_;
  assign new_n13064_ = ~new_n11236_ & (~new_n11233_ | new_n11203_);
  assign new_n13065_ = ~new_n13066_ & new_n13095_;
  assign new_n13066_ = ~new_n13067_ & ~new_n13090_;
  assign new_n13067_ = new_n13085_ & ~new_n13089_ & ~new_n13068_ & ~new_n13088_;
  assign new_n13068_ = ~new_n13083_ & ~new_n13084_ & new_n13076_ & (~new_n13081_ | ~new_n13069_);
  assign new_n13069_ = new_n13075_ & new_n13070_ & new_n13072_;
  assign new_n13070_ = \all_features[5031]  & (\all_features[5030]  | (new_n13071_ & (\all_features[5026]  | \all_features[5027]  | \all_features[5025] )));
  assign new_n13071_ = \all_features[5028]  & \all_features[5029] ;
  assign new_n13072_ = \all_features[5030]  & \all_features[5031]  & (\all_features[5028]  | \all_features[5029]  | new_n13074_ | ~new_n13073_);
  assign new_n13073_ = ~\all_features[5026]  & ~\all_features[5027] ;
  assign new_n13074_ = \all_features[5024]  & \all_features[5025] ;
  assign new_n13075_ = \all_features[5031]  & (\all_features[5029]  | \all_features[5030]  | \all_features[5028] );
  assign new_n13076_ = ~new_n13077_ & ~new_n13079_;
  assign new_n13077_ = ~new_n13078_ & ~\all_features[5031] ;
  assign new_n13078_ = \all_features[5029]  & \all_features[5030]  & (\all_features[5028]  | (\all_features[5026]  & \all_features[5027]  & \all_features[5025] ));
  assign new_n13079_ = ~\all_features[5031]  & (~\all_features[5030]  | (~\all_features[5028]  & ~\all_features[5029]  & ~new_n13080_));
  assign new_n13080_ = \all_features[5026]  & \all_features[5027] ;
  assign new_n13081_ = \all_features[5031]  & (\all_features[5030]  | (\all_features[5029]  & (\all_features[5028]  | ~new_n13082_ | ~new_n13073_)));
  assign new_n13082_ = ~\all_features[5024]  & ~\all_features[5025] ;
  assign new_n13083_ = ~\all_features[5031]  & (~\all_features[5030]  | (~\all_features[5029]  & (new_n13082_ | ~new_n13080_ | ~\all_features[5028] )));
  assign new_n13084_ = ~\all_features[5031]  & (~\all_features[5030]  | ~new_n13071_ | ~new_n13074_ | ~new_n13080_);
  assign new_n13085_ = ~new_n13086_ & (\all_features[5027]  | \all_features[5028]  | \all_features[5029]  | \all_features[5030]  | \all_features[5031] );
  assign new_n13086_ = ~\all_features[5029]  & new_n13087_ & ((~\all_features[5026]  & new_n13082_) | ~\all_features[5028]  | ~\all_features[5027] );
  assign new_n13087_ = ~\all_features[5030]  & ~\all_features[5031] ;
  assign new_n13088_ = new_n13087_ & (~\all_features[5029]  | (~\all_features[5028]  & (~\all_features[5027]  | (~\all_features[5026]  & ~\all_features[5025] ))));
  assign new_n13089_ = new_n13087_ & (~\all_features[5027]  | ~new_n13071_ | (~\all_features[5026]  & ~new_n13074_));
  assign new_n13090_ = new_n13085_ & (~new_n13094_ | (~new_n13091_ & ~new_n13079_ & ~new_n13083_));
  assign new_n13091_ = ~new_n13084_ & ~new_n13077_ & (~new_n13075_ | ~new_n13081_ | new_n13092_);
  assign new_n13092_ = new_n13070_ & new_n13072_ & (new_n13093_ | ~\all_features[5029]  | ~\all_features[5030]  | ~\all_features[5031] );
  assign new_n13093_ = ~\all_features[5027]  & ~\all_features[5028]  & (~\all_features[5026]  | new_n13082_);
  assign new_n13094_ = ~new_n13088_ & ~new_n13089_;
  assign new_n13095_ = new_n13085_ & new_n13076_ & new_n13094_ & ~new_n13083_ & ~new_n13084_;
  assign new_n13096_ = (new_n7949_ & ~new_n13063_ & ~new_n11635_) | (~new_n13065_ & ~new_n13097_ & new_n13098_ & new_n11635_);
  assign new_n13097_ = new_n10169_ & new_n10190_;
  assign new_n13098_ = ~new_n10201_ & ~new_n10204_;
  assign new_n13099_ = ~new_n13100_ & ~new_n13127_;
  assign new_n13100_ = new_n13112_ & (~new_n13116_ | (new_n13119_ & (~new_n13123_ | new_n13101_)));
  assign new_n13101_ = new_n13102_ & (~new_n13106_ | (~new_n13111_ & \all_features[5685]  & \all_features[5686]  & \all_features[5687] ));
  assign new_n13102_ = \all_features[5687]  & (\all_features[5686]  | (~new_n13103_ & \all_features[5685] ));
  assign new_n13103_ = new_n13104_ & ~\all_features[5684]  & new_n13105_;
  assign new_n13104_ = ~\all_features[5680]  & ~\all_features[5681] ;
  assign new_n13105_ = ~\all_features[5682]  & ~\all_features[5683] ;
  assign new_n13106_ = \all_features[5687]  & \all_features[5686]  & ~new_n13109_ & new_n13107_;
  assign new_n13107_ = \all_features[5687]  & (\all_features[5686]  | (new_n13108_ & (\all_features[5682]  | \all_features[5683]  | \all_features[5681] )));
  assign new_n13108_ = \all_features[5684]  & \all_features[5685] ;
  assign new_n13109_ = new_n13105_ & ~\all_features[5685]  & ~new_n13110_ & ~\all_features[5684] ;
  assign new_n13110_ = \all_features[5680]  & \all_features[5681] ;
  assign new_n13111_ = ~\all_features[5683]  & ~\all_features[5684]  & (~\all_features[5682]  | new_n13104_);
  assign new_n13112_ = ~new_n13113_ & ~new_n13115_;
  assign new_n13113_ = ~\all_features[5685]  & new_n13114_ & ((~\all_features[5682]  & new_n13104_) | ~\all_features[5684]  | ~\all_features[5683] );
  assign new_n13114_ = ~\all_features[5686]  & ~\all_features[5687] ;
  assign new_n13115_ = ~\all_features[5687]  & ~\all_features[5686]  & ~\all_features[5685]  & ~\all_features[5683]  & ~\all_features[5684] ;
  assign new_n13116_ = ~new_n13117_ & ~new_n13118_;
  assign new_n13117_ = new_n13114_ & (~\all_features[5683]  | ~new_n13108_ | (~\all_features[5682]  & ~new_n13110_));
  assign new_n13118_ = new_n13114_ & (~\all_features[5685]  | (~\all_features[5684]  & (~\all_features[5683]  | (~\all_features[5682]  & ~\all_features[5681] ))));
  assign new_n13119_ = ~new_n13120_ & ~new_n13122_;
  assign new_n13120_ = ~\all_features[5687]  & (~\all_features[5686]  | (~\all_features[5684]  & ~\all_features[5685]  & ~new_n13121_));
  assign new_n13121_ = \all_features[5682]  & \all_features[5683] ;
  assign new_n13122_ = ~\all_features[5687]  & (~\all_features[5686]  | (~\all_features[5685]  & (new_n13104_ | ~new_n13121_ | ~\all_features[5684] )));
  assign new_n13123_ = ~new_n13124_ & ~new_n13125_;
  assign new_n13124_ = ~\all_features[5687]  & (~\all_features[5686]  | ~new_n13110_ | ~new_n13108_ | ~new_n13121_);
  assign new_n13125_ = ~new_n13126_ & ~\all_features[5687] ;
  assign new_n13126_ = \all_features[5685]  & \all_features[5686]  & (\all_features[5684]  | (\all_features[5682]  & \all_features[5683]  & \all_features[5681] ));
  assign new_n13127_ = new_n13128_ & (new_n13122_ | new_n13125_ | ~new_n13129_ | (new_n13106_ & new_n13102_));
  assign new_n13128_ = new_n13112_ & new_n13116_;
  assign new_n13129_ = ~new_n13120_ & ~new_n13124_;
  assign new_n13130_ = new_n13123_ & new_n13128_ & new_n13119_;
  assign new_n13131_ = new_n13132_ & (new_n10939_ | ~new_n10911_ | (new_n13243_ ? new_n13208_ : new_n13201_));
  assign new_n13132_ = (new_n13133_ & ~new_n7600_) | (new_n10911_ & ~new_n10939_) | (new_n6354_ & new_n6953_ & new_n7600_);
  assign new_n13133_ = (~new_n13134_ | ~new_n13168_) & (~new_n12334_ | ~new_n12337_ | new_n13168_);
  assign new_n13134_ = new_n13135_ & new_n13159_;
  assign new_n13135_ = ~new_n13136_ & ~new_n13158_;
  assign new_n13136_ = new_n13137_ & (~new_n13146_ | (new_n13156_ & new_n13157_ & new_n13153_ & new_n13155_));
  assign new_n13137_ = new_n13138_ & ~new_n13142_ & ~new_n13143_;
  assign new_n13138_ = ~new_n13139_ & (\all_features[3195]  | \all_features[3196]  | \all_features[3197]  | \all_features[3198]  | \all_features[3199] );
  assign new_n13139_ = ~\all_features[3197]  & new_n13141_ & ((~\all_features[3194]  & new_n13140_) | ~\all_features[3196]  | ~\all_features[3195] );
  assign new_n13140_ = ~\all_features[3192]  & ~\all_features[3193] ;
  assign new_n13141_ = ~\all_features[3198]  & ~\all_features[3199] ;
  assign new_n13142_ = new_n13141_ & (~\all_features[3197]  | (~\all_features[3196]  & (~\all_features[3195]  | (~\all_features[3194]  & ~\all_features[3193] ))));
  assign new_n13143_ = new_n13141_ & (~\all_features[3195]  | ~new_n13144_ | (~\all_features[3194]  & ~new_n13145_));
  assign new_n13144_ = \all_features[3196]  & \all_features[3197] ;
  assign new_n13145_ = \all_features[3192]  & \all_features[3193] ;
  assign new_n13146_ = ~new_n13152_ & ~new_n13151_ & ~new_n13147_ & ~new_n13149_;
  assign new_n13147_ = ~\all_features[3199]  & (~\all_features[3198]  | (~\all_features[3197]  & (new_n13140_ | ~new_n13148_ | ~\all_features[3196] )));
  assign new_n13148_ = \all_features[3194]  & \all_features[3195] ;
  assign new_n13149_ = ~new_n13150_ & ~\all_features[3199] ;
  assign new_n13150_ = \all_features[3197]  & \all_features[3198]  & (\all_features[3196]  | (\all_features[3194]  & \all_features[3195]  & \all_features[3193] ));
  assign new_n13151_ = ~\all_features[3199]  & (~\all_features[3198]  | ~new_n13144_ | ~new_n13145_ | ~new_n13148_);
  assign new_n13152_ = ~\all_features[3199]  & (~\all_features[3198]  | (~\all_features[3196]  & ~\all_features[3197]  & ~new_n13148_));
  assign new_n13153_ = \all_features[3199]  & (\all_features[3198]  | (\all_features[3197]  & (\all_features[3196]  | ~new_n13140_ | ~new_n13154_)));
  assign new_n13154_ = ~\all_features[3194]  & ~\all_features[3195] ;
  assign new_n13155_ = \all_features[3199]  & (\all_features[3198]  | (new_n13144_ & (\all_features[3194]  | \all_features[3195]  | \all_features[3193] )));
  assign new_n13156_ = \all_features[3198]  & \all_features[3199]  & (\all_features[3196]  | \all_features[3197]  | new_n13145_ | ~new_n13154_);
  assign new_n13157_ = \all_features[3199]  & (\all_features[3197]  | \all_features[3198]  | \all_features[3196] );
  assign new_n13158_ = new_n13137_ & new_n13146_;
  assign new_n13159_ = ~new_n13160_ & ~new_n13164_;
  assign new_n13160_ = new_n13138_ & (new_n13143_ | new_n13142_ | (~new_n13147_ & ~new_n13152_ & ~new_n13161_));
  assign new_n13161_ = ~new_n13151_ & ~new_n13149_ & (~new_n13157_ | ~new_n13153_ | new_n13162_);
  assign new_n13162_ = new_n13155_ & new_n13156_ & (new_n13163_ | ~\all_features[3197]  | ~\all_features[3198]  | ~\all_features[3199] );
  assign new_n13163_ = ~\all_features[3195]  & ~\all_features[3196]  & (~\all_features[3194]  | new_n13140_);
  assign new_n13164_ = ~new_n13165_ & (\all_features[3195]  | \all_features[3196]  | \all_features[3197]  | \all_features[3198]  | \all_features[3199] );
  assign new_n13165_ = ~new_n13139_ & (new_n13142_ | (~new_n13143_ & (new_n13152_ | (~new_n13147_ & ~new_n13166_))));
  assign new_n13166_ = ~new_n13149_ & (new_n13151_ | (new_n13157_ & (~new_n13153_ | (~new_n13167_ & new_n13155_))));
  assign new_n13167_ = ~\all_features[3197]  & \all_features[3198]  & \all_features[3199]  & (\all_features[3196]  ? new_n13154_ : (new_n13145_ | ~new_n13154_));
  assign new_n13168_ = ~new_n13197_ & new_n13169_;
  assign new_n13169_ = ~new_n13170_ & ~new_n13196_;
  assign new_n13170_ = new_n13183_ & (~new_n13171_ | (new_n13194_ & new_n13195_ & new_n13191_ & new_n13192_));
  assign new_n13171_ = new_n13172_ & new_n13179_;
  assign new_n13172_ = ~new_n13173_ & ~new_n13175_;
  assign new_n13173_ = ~new_n13174_ & ~\all_features[3895] ;
  assign new_n13174_ = \all_features[3893]  & \all_features[3894]  & (\all_features[3892]  | (\all_features[3890]  & \all_features[3891]  & \all_features[3889] ));
  assign new_n13175_ = ~\all_features[3895]  & (~\all_features[3894]  | ~new_n13176_ | ~new_n13177_ | ~new_n13178_);
  assign new_n13176_ = \all_features[3892]  & \all_features[3893] ;
  assign new_n13177_ = \all_features[3888]  & \all_features[3889] ;
  assign new_n13178_ = \all_features[3890]  & \all_features[3891] ;
  assign new_n13179_ = ~new_n13180_ & ~new_n13181_;
  assign new_n13180_ = ~\all_features[3895]  & (~\all_features[3894]  | (~\all_features[3892]  & ~\all_features[3893]  & ~new_n13178_));
  assign new_n13181_ = ~\all_features[3895]  & (~\all_features[3894]  | (~\all_features[3893]  & (new_n13182_ | ~new_n13178_ | ~\all_features[3892] )));
  assign new_n13182_ = ~\all_features[3888]  & ~\all_features[3889] ;
  assign new_n13183_ = new_n13184_ & new_n13188_;
  assign new_n13184_ = ~new_n13185_ & ~new_n13187_;
  assign new_n13185_ = new_n13186_ & (~\all_features[3893]  | (~\all_features[3892]  & (~\all_features[3891]  | (~\all_features[3890]  & ~\all_features[3889] ))));
  assign new_n13186_ = ~\all_features[3894]  & ~\all_features[3895] ;
  assign new_n13187_ = new_n13186_ & (~\all_features[3891]  | ~new_n13176_ | (~\all_features[3890]  & ~new_n13177_));
  assign new_n13188_ = ~new_n13189_ & ~new_n13190_;
  assign new_n13189_ = ~\all_features[3893]  & new_n13186_ & ((~\all_features[3890]  & new_n13182_) | ~\all_features[3892]  | ~\all_features[3891] );
  assign new_n13190_ = ~\all_features[3895]  & ~\all_features[3894]  & ~\all_features[3893]  & ~\all_features[3891]  & ~\all_features[3892] ;
  assign new_n13191_ = \all_features[3895]  & (\all_features[3894]  | (new_n13176_ & (\all_features[3890]  | \all_features[3891]  | \all_features[3889] )));
  assign new_n13192_ = \all_features[3894]  & \all_features[3895]  & (\all_features[3892]  | \all_features[3893]  | new_n13177_ | ~new_n13193_);
  assign new_n13193_ = ~\all_features[3890]  & ~\all_features[3891] ;
  assign new_n13194_ = \all_features[3895]  & (\all_features[3894]  | (\all_features[3893]  & (\all_features[3892]  | ~new_n13193_ | ~new_n13182_)));
  assign new_n13195_ = \all_features[3895]  & (\all_features[3893]  | \all_features[3894]  | \all_features[3892] );
  assign new_n13196_ = new_n13171_ & new_n13183_;
  assign new_n13197_ = new_n13188_ & (~new_n13184_ | (~new_n13198_ & new_n13179_));
  assign new_n13198_ = new_n13172_ & ((~new_n13199_ & new_n13192_ & new_n13191_) | ~new_n13195_ | ~new_n13194_);
  assign new_n13199_ = \all_features[3895]  & \all_features[3894]  & ~new_n13200_ & \all_features[3893] ;
  assign new_n13200_ = ~\all_features[3891]  & ~\all_features[3892]  & (~\all_features[3890]  | new_n13182_);
  assign new_n13201_ = new_n13202_ ? new_n10873_ : new_n9689_;
  assign new_n13202_ = new_n13203_ & ~new_n11675_ & ~new_n11699_;
  assign new_n13203_ = ~new_n11700_ & ~new_n13204_;
  assign new_n13204_ = ~new_n11696_ & (new_n11694_ | (~new_n11697_ & ~new_n13205_));
  assign new_n13205_ = ~new_n11698_ & (new_n11685_ | (~new_n11686_ & (new_n11683_ | (~new_n13206_ & ~new_n11692_))));
  assign new_n13206_ = new_n11681_ & (~new_n11678_ | (new_n11690_ & (new_n13207_ | ~new_n11688_)));
  assign new_n13207_ = \all_features[3638]  & \all_features[3639]  & (\all_features[3637]  | (~new_n11679_ & \all_features[3636] ));
  assign new_n13208_ = (new_n7409_ & new_n13242_ & (new_n13238_ | ~new_n13209_)) | (new_n10130_ & new_n10153_ & (~new_n13242_ | (~new_n13238_ & new_n13209_)));
  assign new_n13209_ = ~new_n13210_ & ~new_n13234_;
  assign new_n13210_ = ~new_n13232_ & ~new_n13231_ & (~new_n13225_ | (~new_n13211_ & ~new_n13229_ & ~new_n13233_));
  assign new_n13211_ = ~new_n13220_ & ~new_n13221_ & (~new_n13224_ | ~new_n13223_ | new_n13212_);
  assign new_n13212_ = new_n13213_ & new_n13215_ & (new_n13218_ | ~\all_features[4349]  | ~\all_features[4350]  | ~\all_features[4351] );
  assign new_n13213_ = \all_features[4351]  & (\all_features[4350]  | (new_n13214_ & (\all_features[4346]  | \all_features[4347]  | \all_features[4345] )));
  assign new_n13214_ = \all_features[4348]  & \all_features[4349] ;
  assign new_n13215_ = \all_features[4350]  & \all_features[4351]  & (\all_features[4348]  | \all_features[4349]  | new_n13216_ | ~new_n13217_);
  assign new_n13216_ = \all_features[4344]  & \all_features[4345] ;
  assign new_n13217_ = ~\all_features[4346]  & ~\all_features[4347] ;
  assign new_n13218_ = ~\all_features[4347]  & ~\all_features[4348]  & (~\all_features[4346]  | new_n13219_);
  assign new_n13219_ = ~\all_features[4344]  & ~\all_features[4345] ;
  assign new_n13220_ = ~\all_features[4351]  & (~new_n13214_ | ~\all_features[4346]  | ~\all_features[4347]  | ~\all_features[4350]  | ~new_n13216_);
  assign new_n13221_ = ~new_n13222_ & ~\all_features[4351] ;
  assign new_n13222_ = \all_features[4349]  & \all_features[4350]  & (\all_features[4348]  | (\all_features[4346]  & \all_features[4347]  & \all_features[4345] ));
  assign new_n13223_ = \all_features[4351]  & (\all_features[4350]  | (\all_features[4349]  & (\all_features[4348]  | ~new_n13217_ | ~new_n13219_)));
  assign new_n13224_ = \all_features[4351]  & (\all_features[4349]  | \all_features[4350]  | \all_features[4348] );
  assign new_n13225_ = ~new_n13226_ & ~new_n13228_;
  assign new_n13226_ = new_n13227_ & (~\all_features[4347]  | ~new_n13214_ | (~\all_features[4346]  & ~new_n13216_));
  assign new_n13227_ = ~\all_features[4350]  & ~\all_features[4351] ;
  assign new_n13228_ = new_n13227_ & (~\all_features[4349]  | (~\all_features[4348]  & (~\all_features[4347]  | (~\all_features[4346]  & ~\all_features[4345] ))));
  assign new_n13229_ = ~\all_features[4351]  & (~\all_features[4350]  | new_n13230_);
  assign new_n13230_ = ~\all_features[4349]  & (new_n13219_ | ~\all_features[4347]  | ~\all_features[4348]  | ~\all_features[4346] );
  assign new_n13231_ = ~\all_features[4349]  & new_n13227_ & ((~\all_features[4346]  & new_n13219_) | ~\all_features[4348]  | ~\all_features[4347] );
  assign new_n13232_ = ~\all_features[4351]  & ~\all_features[4350]  & ~\all_features[4349]  & ~\all_features[4347]  & ~\all_features[4348] ;
  assign new_n13233_ = ~\all_features[4351]  & (~\all_features[4350]  | (~\all_features[4349]  & ~\all_features[4348]  & (~\all_features[4347]  | ~\all_features[4346] )));
  assign new_n13234_ = ~new_n13235_ & ~new_n13232_;
  assign new_n13235_ = ~new_n13231_ & (new_n13228_ | (~new_n13226_ & (new_n13233_ | (~new_n13229_ & ~new_n13236_))));
  assign new_n13236_ = ~new_n13221_ & (new_n13220_ | (new_n13224_ & (~new_n13223_ | (~new_n13237_ & new_n13213_))));
  assign new_n13237_ = ~\all_features[4349]  & \all_features[4350]  & \all_features[4351]  & (\all_features[4348]  ? new_n13217_ : (new_n13216_ | ~new_n13217_));
  assign new_n13238_ = ~new_n13232_ & ~new_n13231_ & ~new_n13228_ & ~new_n13239_ & ~new_n13226_;
  assign new_n13239_ = ~new_n13229_ & ~new_n13220_ & new_n13240_ & (~new_n13223_ | ~new_n13241_);
  assign new_n13240_ = ~new_n13221_ & ~new_n13233_;
  assign new_n13241_ = new_n13224_ & new_n13213_ & new_n13215_;
  assign new_n13242_ = new_n13225_ & new_n13240_ & ~new_n13232_ & ~new_n13220_ & ~new_n13229_ & ~new_n13231_;
  assign new_n13243_ = new_n13244_ & new_n13270_;
  assign new_n13244_ = ~new_n13245_ & ~new_n13269_;
  assign new_n13245_ = new_n13263_ & ~new_n13268_ & ~new_n13246_ & ~new_n13267_;
  assign new_n13246_ = ~new_n13256_ & ~new_n13262_ & new_n13252_ & (~new_n13260_ | ~new_n13258_ | ~new_n13247_);
  assign new_n13247_ = \all_features[4991]  & (\all_features[4990]  | (~new_n13251_ & new_n13248_));
  assign new_n13248_ = \all_features[4989]  & (\all_features[4988]  | ~new_n13250_ | ~new_n13249_);
  assign new_n13249_ = ~\all_features[4986]  & ~\all_features[4987] ;
  assign new_n13250_ = ~\all_features[4984]  & ~\all_features[4985] ;
  assign new_n13251_ = ~\all_features[4988]  & ~\all_features[4989] ;
  assign new_n13252_ = ~new_n13253_ & ~new_n13255_;
  assign new_n13253_ = ~new_n13254_ & ~\all_features[4991] ;
  assign new_n13254_ = \all_features[4989]  & \all_features[4990]  & (\all_features[4988]  | (\all_features[4986]  & \all_features[4987]  & \all_features[4985] ));
  assign new_n13255_ = ~\all_features[4991]  & (~\all_features[4990]  | (new_n13251_ & (~\all_features[4987]  | ~\all_features[4986] )));
  assign new_n13256_ = ~\all_features[4991]  & (~\all_features[4990]  | new_n13257_);
  assign new_n13257_ = ~\all_features[4989]  & (new_n13250_ | ~\all_features[4987]  | ~\all_features[4988]  | ~\all_features[4986] );
  assign new_n13258_ = \all_features[4990]  & \all_features[4991]  & (new_n13259_ | ~new_n13251_ | ~new_n13249_);
  assign new_n13259_ = \all_features[4984]  & \all_features[4985] ;
  assign new_n13260_ = \all_features[4991]  & (\all_features[4990]  | (new_n13261_ & (\all_features[4986]  | \all_features[4987]  | \all_features[4985] )));
  assign new_n13261_ = \all_features[4988]  & \all_features[4989] ;
  assign new_n13262_ = ~\all_features[4991]  & (~new_n13261_ | ~\all_features[4986]  | ~\all_features[4987]  | ~\all_features[4990]  | ~new_n13259_);
  assign new_n13263_ = ~new_n13264_ & ~new_n13266_;
  assign new_n13264_ = ~\all_features[4989]  & new_n13265_ & ((~\all_features[4986]  & new_n13250_) | ~\all_features[4988]  | ~\all_features[4987] );
  assign new_n13265_ = ~\all_features[4990]  & ~\all_features[4991] ;
  assign new_n13266_ = ~\all_features[4991]  & ~\all_features[4990]  & ~\all_features[4989]  & ~\all_features[4987]  & ~\all_features[4988] ;
  assign new_n13267_ = new_n13265_ & (~\all_features[4989]  | (~\all_features[4988]  & (~\all_features[4987]  | (~\all_features[4986]  & ~\all_features[4985] ))));
  assign new_n13268_ = new_n13265_ & (~\all_features[4987]  | ~new_n13261_ | (~\all_features[4986]  & ~new_n13259_));
  assign new_n13269_ = new_n13252_ & new_n13263_ & ~new_n13268_ & ~new_n13267_ & ~new_n13256_ & ~new_n13262_;
  assign new_n13270_ = ~new_n13271_ & (new_n13266_ | (~new_n13264_ & (new_n13267_ | new_n13275_)));
  assign new_n13271_ = new_n13263_ & (new_n13268_ | new_n13267_ | (~new_n13255_ & ~new_n13272_ & ~new_n13256_));
  assign new_n13272_ = ~new_n13253_ & ~new_n13262_ & (~new_n13247_ | (~new_n13273_ & new_n13258_ & new_n13260_));
  assign new_n13273_ = \all_features[4991]  & \all_features[4990]  & ~new_n13274_ & \all_features[4989] ;
  assign new_n13274_ = ~\all_features[4987]  & ~\all_features[4988]  & (~\all_features[4986]  | new_n13250_);
  assign new_n13275_ = ~new_n13268_ & (new_n13255_ | (~new_n13256_ & (new_n13253_ | (~new_n13276_ & ~new_n13262_))));
  assign new_n13276_ = \all_features[4991]  & ((~new_n13277_ & \all_features[4990]  & new_n13260_) | (~new_n13251_ & ((~new_n13277_ & new_n13260_) | (~new_n13248_ & ~\all_features[4990] ))));
  assign new_n13277_ = ~\all_features[4989]  & \all_features[4990]  & \all_features[4991]  & (\all_features[4988]  ? new_n13249_ : (new_n13259_ | ~new_n13249_));
  assign new_n13278_ = ~new_n13279_ & new_n13442_;
  assign new_n13279_ = new_n13280_ & new_n13351_ & (~new_n13404_ | ~new_n13405_) & (~new_n13403_ | ~new_n13407_);
  assign new_n13280_ = ~new_n13281_ & (~new_n13346_ | (~new_n13347_ & ~new_n13349_) | (~new_n12118_ & new_n13349_));
  assign new_n13281_ = new_n13329_ & new_n13282_ & new_n13318_;
  assign new_n13282_ = ~new_n6884_ & new_n13283_;
  assign new_n13283_ = new_n13316_ & (new_n13314_ | ~new_n13284_);
  assign new_n13284_ = ~new_n13285_ & (new_n13310_ | (~new_n13311_ & ~new_n13309_));
  assign new_n13285_ = ~new_n13309_ & ~new_n13310_ & (~new_n13302_ | (~new_n13286_ & new_n13306_));
  assign new_n13286_ = new_n13290_ & ((~new_n13300_ & new_n13298_ & new_n13297_) | ~new_n13301_ | ~new_n13287_);
  assign new_n13287_ = \all_features[3311]  & (\all_features[3310]  | new_n13288_);
  assign new_n13288_ = \all_features[3309]  & (\all_features[3306]  | \all_features[3307]  | \all_features[3308]  | ~new_n13289_);
  assign new_n13289_ = ~\all_features[3304]  & ~\all_features[3305] ;
  assign new_n13290_ = ~new_n13291_ & ~new_n13293_;
  assign new_n13291_ = ~new_n13292_ & ~\all_features[3311] ;
  assign new_n13292_ = \all_features[3309]  & \all_features[3310]  & (\all_features[3308]  | (\all_features[3306]  & \all_features[3307]  & \all_features[3305] ));
  assign new_n13293_ = ~\all_features[3311]  & (~\all_features[3310]  | ~new_n13294_ | ~new_n13295_ | ~new_n13296_);
  assign new_n13294_ = \all_features[3304]  & \all_features[3305] ;
  assign new_n13295_ = \all_features[3308]  & \all_features[3309] ;
  assign new_n13296_ = \all_features[3306]  & \all_features[3307] ;
  assign new_n13297_ = \all_features[3311]  & (\all_features[3310]  | (new_n13295_ & (\all_features[3306]  | \all_features[3307]  | \all_features[3305] )));
  assign new_n13298_ = new_n13299_ & (new_n13294_ | \all_features[3306]  | \all_features[3307]  | \all_features[3308]  | \all_features[3309] );
  assign new_n13299_ = \all_features[3310]  & \all_features[3311] ;
  assign new_n13300_ = new_n13299_ & \all_features[3309]  & ((~new_n13289_ & \all_features[3306] ) | \all_features[3308]  | \all_features[3307] );
  assign new_n13301_ = \all_features[3311]  & (\all_features[3309]  | \all_features[3310]  | \all_features[3308] );
  assign new_n13302_ = ~new_n13303_ & ~new_n13305_;
  assign new_n13303_ = new_n13304_ & (~\all_features[3309]  | (~\all_features[3308]  & (~\all_features[3307]  | (~\all_features[3306]  & ~\all_features[3305] ))));
  assign new_n13304_ = ~\all_features[3310]  & ~\all_features[3311] ;
  assign new_n13305_ = new_n13304_ & (~\all_features[3307]  | ~new_n13295_ | (~\all_features[3306]  & ~new_n13294_));
  assign new_n13306_ = ~new_n13307_ & ~new_n13308_;
  assign new_n13307_ = ~\all_features[3311]  & (~\all_features[3310]  | (~\all_features[3308]  & ~\all_features[3309]  & ~new_n13296_));
  assign new_n13308_ = ~\all_features[3311]  & (~\all_features[3310]  | (~\all_features[3309]  & (new_n13289_ | ~\all_features[3308]  | ~new_n13296_)));
  assign new_n13309_ = ~\all_features[3309]  & new_n13304_ & ((~\all_features[3306]  & new_n13289_) | ~\all_features[3308]  | ~\all_features[3307] );
  assign new_n13310_ = ~\all_features[3311]  & ~\all_features[3310]  & ~\all_features[3309]  & ~\all_features[3307]  & ~\all_features[3308] ;
  assign new_n13311_ = ~new_n13303_ & (new_n13305_ | (~new_n13307_ & (new_n13308_ | (~new_n13312_ & ~new_n13291_))));
  assign new_n13312_ = ~new_n13293_ & (~new_n13301_ | (new_n13287_ & (~new_n13297_ | (~new_n13313_ & new_n13298_))));
  assign new_n13313_ = new_n13299_ & (\all_features[3309]  | (\all_features[3308]  & (\all_features[3307]  | \all_features[3306] )));
  assign new_n13314_ = ~new_n13310_ & ~new_n13305_ & ~new_n13303_ & ~new_n13315_ & ~new_n13309_;
  assign new_n13315_ = new_n13306_ & new_n13290_ & (~new_n13298_ | ~new_n13301_ | ~new_n13287_ | ~new_n13297_);
  assign new_n13316_ = new_n13302_ & new_n13317_ & ~new_n13308_ & ~new_n13309_ & ~new_n13291_ & ~new_n13307_;
  assign new_n13317_ = ~new_n13293_ & ~new_n13310_;
  assign new_n13318_ = ~new_n13319_ & new_n13328_;
  assign new_n13319_ = ~new_n13320_ & ~new_n13324_;
  assign new_n13320_ = ~new_n13321_ & (\all_features[3451]  | \all_features[3452]  | \all_features[3453]  | \all_features[3454]  | \all_features[3455] );
  assign new_n13321_ = ~new_n10980_ & (new_n10983_ | (~new_n10984_ & (new_n10993_ | (~new_n10988_ & ~new_n13322_))));
  assign new_n13322_ = ~new_n10990_ & (new_n10992_ | (new_n10998_ & (~new_n10994_ | (~new_n13323_ & new_n10996_))));
  assign new_n13323_ = ~\all_features[3453]  & \all_features[3454]  & \all_features[3455]  & (\all_features[3452]  ? new_n10995_ : (new_n10986_ | ~new_n10995_));
  assign new_n13324_ = new_n10979_ & (new_n10984_ | new_n10983_ | (~new_n10988_ & ~new_n10993_ & ~new_n13325_));
  assign new_n13325_ = ~new_n10992_ & ~new_n10990_ & (~new_n10998_ | ~new_n10994_ | new_n13326_);
  assign new_n13326_ = new_n10996_ & new_n10997_ & (new_n13327_ | ~\all_features[3453]  | ~\all_features[3454]  | ~\all_features[3455] );
  assign new_n13327_ = ~\all_features[3451]  & ~\all_features[3452]  & (~\all_features[3450]  | new_n10981_);
  assign new_n13328_ = new_n10977_ & new_n10999_;
  assign new_n13329_ = new_n13336_ & new_n13330_ & ~new_n13345_ & ~new_n13343_ & ~new_n13340_ & ~new_n13342_;
  assign new_n13330_ = ~new_n13331_ & ~new_n13335_;
  assign new_n13331_ = ~\all_features[1735]  & (~\all_features[1734]  | ~new_n13332_ | ~new_n13333_ | ~new_n13334_);
  assign new_n13332_ = \all_features[1728]  & \all_features[1729] ;
  assign new_n13333_ = \all_features[1732]  & \all_features[1733] ;
  assign new_n13334_ = \all_features[1730]  & \all_features[1731] ;
  assign new_n13335_ = ~\all_features[1735]  & ~\all_features[1734]  & ~\all_features[1733]  & ~\all_features[1731]  & ~\all_features[1732] ;
  assign new_n13336_ = ~new_n13337_ & ~new_n13339_;
  assign new_n13337_ = new_n13338_ & (~\all_features[1731]  | ~new_n13333_ | (~\all_features[1730]  & ~new_n13332_));
  assign new_n13338_ = ~\all_features[1734]  & ~\all_features[1735] ;
  assign new_n13339_ = new_n13338_ & (~\all_features[1733]  | (~\all_features[1732]  & (~\all_features[1731]  | (~\all_features[1730]  & ~\all_features[1729] ))));
  assign new_n13340_ = ~new_n13341_ & ~\all_features[1735] ;
  assign new_n13341_ = \all_features[1733]  & \all_features[1734]  & (\all_features[1732]  | (\all_features[1730]  & \all_features[1731]  & \all_features[1729] ));
  assign new_n13342_ = ~\all_features[1735]  & (~\all_features[1734]  | (~\all_features[1732]  & ~\all_features[1733]  & ~new_n13334_));
  assign new_n13343_ = ~\all_features[1733]  & new_n13338_ & ((~\all_features[1730]  & new_n13344_) | ~\all_features[1732]  | ~\all_features[1731] );
  assign new_n13344_ = ~\all_features[1728]  & ~\all_features[1729] ;
  assign new_n13345_ = ~\all_features[1735]  & (~\all_features[1734]  | (~\all_features[1733]  & (new_n13344_ | ~\all_features[1732]  | ~new_n13334_)));
  assign new_n13346_ = ~new_n9312_ & new_n6884_;
  assign new_n13347_ = ~new_n12269_ & new_n13348_;
  assign new_n13348_ = ~new_n12298_ & ~new_n12301_;
  assign new_n13349_ = new_n13350_ & ~new_n11944_ & ~new_n11965_;
  assign new_n13350_ = ~new_n11975_ & ~new_n11972_;
  assign new_n13351_ = (~new_n13352_ | ~new_n13401_) & (~new_n13365_ | ~new_n13364_);
  assign new_n13352_ = ~new_n13354_ & new_n13353_;
  assign new_n13353_ = ~new_n6884_ & ~new_n13283_;
  assign new_n13354_ = new_n7159_ & (new_n7137_ | ~new_n13355_);
  assign new_n13355_ = ~new_n13356_ & ~new_n13360_;
  assign new_n13356_ = new_n7154_ & (~new_n7160_ | (~new_n13357_ & ~new_n7152_ & ~new_n7142_));
  assign new_n13357_ = ~new_n7144_ & ~new_n7140_ & (~new_n7153_ | ~new_n7147_ | new_n13358_);
  assign new_n13358_ = new_n7150_ & new_n7151_ & (new_n13359_ | ~\all_features[4333]  | ~\all_features[4334]  | ~\all_features[4335] );
  assign new_n13359_ = ~\all_features[4331]  & ~\all_features[4332]  & (~\all_features[4330]  | new_n7149_);
  assign new_n13360_ = ~new_n13361_ & (\all_features[4331]  | \all_features[4332]  | \all_features[4333]  | \all_features[4334]  | \all_features[4335] );
  assign new_n13361_ = ~new_n7155_ & (new_n7157_ | (~new_n7158_ & (new_n7142_ | (~new_n7152_ & ~new_n13362_))));
  assign new_n13362_ = ~new_n7140_ & (new_n7144_ | (new_n7153_ & (~new_n7147_ | (~new_n13363_ & new_n7150_))));
  assign new_n13363_ = ~\all_features[4333]  & \all_features[4334]  & \all_features[4335]  & (\all_features[4332]  ? new_n7148_ : (new_n7146_ | ~new_n7148_));
  assign new_n13364_ = new_n6884_ & new_n9312_;
  assign new_n13365_ = new_n13367_ ? ~new_n13366_ : ~new_n7581_;
  assign new_n13366_ = ~new_n7991_ & (~new_n7988_ | ~new_n7958_);
  assign new_n13367_ = new_n13368_ & new_n13392_;
  assign new_n13368_ = ~new_n13369_ & ~new_n13391_;
  assign new_n13369_ = new_n13370_ & (~new_n13379_ | (new_n13389_ & new_n13390_ & new_n13386_ & new_n13388_));
  assign new_n13370_ = new_n13371_ & ~new_n13375_ & ~new_n13376_;
  assign new_n13371_ = ~new_n13372_ & (\all_features[1963]  | \all_features[1964]  | \all_features[1965]  | \all_features[1966]  | \all_features[1967] );
  assign new_n13372_ = ~\all_features[1965]  & new_n13374_ & ((~\all_features[1962]  & new_n13373_) | ~\all_features[1964]  | ~\all_features[1963] );
  assign new_n13373_ = ~\all_features[1960]  & ~\all_features[1961] ;
  assign new_n13374_ = ~\all_features[1966]  & ~\all_features[1967] ;
  assign new_n13375_ = new_n13374_ & (~\all_features[1965]  | (~\all_features[1964]  & (~\all_features[1963]  | (~\all_features[1962]  & ~\all_features[1961] ))));
  assign new_n13376_ = new_n13374_ & (~\all_features[1963]  | ~new_n13377_ | (~\all_features[1962]  & ~new_n13378_));
  assign new_n13377_ = \all_features[1964]  & \all_features[1965] ;
  assign new_n13378_ = \all_features[1960]  & \all_features[1961] ;
  assign new_n13379_ = ~new_n13385_ & ~new_n13384_ & ~new_n13380_ & ~new_n13382_;
  assign new_n13380_ = ~\all_features[1967]  & (~\all_features[1966]  | (~\all_features[1965]  & (new_n13373_ | ~new_n13381_ | ~\all_features[1964] )));
  assign new_n13381_ = \all_features[1962]  & \all_features[1963] ;
  assign new_n13382_ = ~new_n13383_ & ~\all_features[1967] ;
  assign new_n13383_ = \all_features[1965]  & \all_features[1966]  & (\all_features[1964]  | (\all_features[1962]  & \all_features[1963]  & \all_features[1961] ));
  assign new_n13384_ = ~\all_features[1967]  & (~\all_features[1966]  | ~new_n13377_ | ~new_n13378_ | ~new_n13381_);
  assign new_n13385_ = ~\all_features[1967]  & (~\all_features[1966]  | (~\all_features[1964]  & ~\all_features[1965]  & ~new_n13381_));
  assign new_n13386_ = \all_features[1967]  & (\all_features[1966]  | (\all_features[1965]  & (\all_features[1964]  | ~new_n13373_ | ~new_n13387_)));
  assign new_n13387_ = ~\all_features[1962]  & ~\all_features[1963] ;
  assign new_n13388_ = \all_features[1967]  & (\all_features[1966]  | (new_n13377_ & (\all_features[1962]  | \all_features[1963]  | \all_features[1961] )));
  assign new_n13389_ = \all_features[1966]  & \all_features[1967]  & (\all_features[1964]  | \all_features[1965]  | new_n13378_ | ~new_n13387_);
  assign new_n13390_ = \all_features[1967]  & (\all_features[1965]  | \all_features[1966]  | \all_features[1964] );
  assign new_n13391_ = new_n13370_ & new_n13379_;
  assign new_n13392_ = ~new_n13393_ & ~new_n13397_;
  assign new_n13393_ = new_n13371_ & (new_n13376_ | new_n13375_ | (~new_n13380_ & ~new_n13385_ & ~new_n13394_));
  assign new_n13394_ = ~new_n13384_ & ~new_n13382_ & (~new_n13390_ | ~new_n13386_ | new_n13395_);
  assign new_n13395_ = new_n13388_ & new_n13389_ & (new_n13396_ | ~\all_features[1965]  | ~\all_features[1966]  | ~\all_features[1967] );
  assign new_n13396_ = ~\all_features[1963]  & ~\all_features[1964]  & (~\all_features[1962]  | new_n13373_);
  assign new_n13397_ = ~new_n13398_ & (\all_features[1963]  | \all_features[1964]  | \all_features[1965]  | \all_features[1966]  | \all_features[1967] );
  assign new_n13398_ = ~new_n13372_ & (new_n13375_ | (~new_n13376_ & (new_n13385_ | (~new_n13380_ & ~new_n13399_))));
  assign new_n13399_ = ~new_n13382_ & (new_n13384_ | (new_n13390_ & (~new_n13386_ | (~new_n13400_ & new_n13388_))));
  assign new_n13400_ = ~\all_features[1965]  & \all_features[1966]  & \all_features[1967]  & (\all_features[1964]  ? new_n13387_ : (new_n13378_ | ~new_n13387_));
  assign new_n13401_ = new_n13402_ & new_n9203_;
  assign new_n13402_ = new_n9172_ & new_n9193_;
  assign new_n13403_ = new_n13353_ & new_n13354_;
  assign new_n13404_ = ~new_n13329_ & new_n13282_;
  assign new_n13405_ = new_n8061_ & new_n13406_;
  assign new_n13406_ = new_n8094_ & new_n8097_;
  assign new_n13407_ = ~new_n13408_ & new_n13437_;
  assign new_n13408_ = ~new_n13409_ & ~new_n13433_;
  assign new_n13409_ = new_n13430_ & (~new_n13424_ | (~new_n13410_ & ~new_n13428_ & ~new_n13432_));
  assign new_n13410_ = ~new_n13421_ & ~new_n13420_ & (~new_n13423_ | ~new_n13419_ | new_n13411_);
  assign new_n13411_ = new_n13412_ & new_n13414_ & (new_n13417_ | ~\all_features[3429]  | ~\all_features[3430]  | ~\all_features[3431] );
  assign new_n13412_ = \all_features[3431]  & (\all_features[3430]  | (new_n13413_ & (\all_features[3426]  | \all_features[3427]  | \all_features[3425] )));
  assign new_n13413_ = \all_features[3428]  & \all_features[3429] ;
  assign new_n13414_ = \all_features[3430]  & \all_features[3431]  & (\all_features[3428]  | \all_features[3429]  | new_n13415_ | ~new_n13416_);
  assign new_n13415_ = \all_features[3424]  & \all_features[3425] ;
  assign new_n13416_ = ~\all_features[3426]  & ~\all_features[3427] ;
  assign new_n13417_ = ~\all_features[3427]  & ~\all_features[3428]  & (~\all_features[3426]  | new_n13418_);
  assign new_n13418_ = ~\all_features[3424]  & ~\all_features[3425] ;
  assign new_n13419_ = \all_features[3431]  & (\all_features[3430]  | (\all_features[3429]  & (\all_features[3428]  | ~new_n13418_ | ~new_n13416_)));
  assign new_n13420_ = ~\all_features[3431]  & (~new_n13413_ | ~\all_features[3426]  | ~\all_features[3427]  | ~\all_features[3430]  | ~new_n13415_);
  assign new_n13421_ = ~new_n13422_ & ~\all_features[3431] ;
  assign new_n13422_ = \all_features[3429]  & \all_features[3430]  & (\all_features[3428]  | (\all_features[3426]  & \all_features[3427]  & \all_features[3425] ));
  assign new_n13423_ = \all_features[3431]  & (\all_features[3429]  | \all_features[3430]  | \all_features[3428] );
  assign new_n13424_ = ~new_n13425_ & ~new_n13427_;
  assign new_n13425_ = new_n13426_ & (~\all_features[3427]  | ~new_n13413_ | (~\all_features[3426]  & ~new_n13415_));
  assign new_n13426_ = ~\all_features[3430]  & ~\all_features[3431] ;
  assign new_n13427_ = new_n13426_ & (~\all_features[3429]  | (~\all_features[3428]  & (~\all_features[3427]  | (~\all_features[3426]  & ~\all_features[3425] ))));
  assign new_n13428_ = ~\all_features[3431]  & (~\all_features[3430]  | new_n13429_);
  assign new_n13429_ = ~\all_features[3429]  & (new_n13418_ | ~\all_features[3427]  | ~\all_features[3428]  | ~\all_features[3426] );
  assign new_n13430_ = ~new_n13431_ & (\all_features[3427]  | \all_features[3428]  | \all_features[3429]  | \all_features[3430]  | \all_features[3431] );
  assign new_n13431_ = ~\all_features[3429]  & new_n13426_ & ((~\all_features[3426]  & new_n13418_) | ~\all_features[3428]  | ~\all_features[3427] );
  assign new_n13432_ = ~\all_features[3431]  & (~\all_features[3430]  | (~\all_features[3429]  & ~\all_features[3428]  & (~\all_features[3427]  | ~\all_features[3426] )));
  assign new_n13433_ = ~new_n13434_ & (\all_features[3427]  | \all_features[3428]  | \all_features[3429]  | \all_features[3430]  | \all_features[3431] );
  assign new_n13434_ = ~new_n13431_ & (new_n13427_ | (~new_n13425_ & (new_n13432_ | (~new_n13428_ & ~new_n13435_))));
  assign new_n13435_ = ~new_n13421_ & (new_n13420_ | (new_n13423_ & (~new_n13419_ | (~new_n13436_ & new_n13412_))));
  assign new_n13436_ = ~\all_features[3429]  & \all_features[3430]  & \all_features[3431]  & (\all_features[3428]  ? new_n13416_ : (new_n13415_ | ~new_n13416_));
  assign new_n13437_ = new_n13438_ & new_n13441_;
  assign new_n13438_ = new_n13424_ & new_n13430_ & (new_n13428_ | new_n13439_ | new_n13420_ | ~new_n13440_);
  assign new_n13439_ = new_n13423_ & new_n13419_ & new_n13412_ & new_n13414_;
  assign new_n13440_ = ~new_n13421_ & ~new_n13432_;
  assign new_n13441_ = new_n13424_ & new_n13440_ & new_n13430_ & ~new_n13428_ & ~new_n13420_;
  assign new_n13442_ = new_n13443_ & new_n13444_;
  assign new_n13443_ = (~new_n13346_ | (new_n13349_ ? new_n12118_ : new_n13347_)) & (~new_n13352_ | new_n13401_);
  assign new_n13444_ = (new_n13407_ | ~new_n13403_) & (new_n13365_ | ~new_n13364_) & (new_n13405_ | ~new_n13404_);
  assign new_n13445_ = ~new_n13446_ & ~new_n13561_;
  assign new_n13446_ = new_n13558_ & ~new_n13515_ & new_n13447_;
  assign new_n13447_ = new_n13448_ & (new_n6354_ | new_n13514_ | new_n8188_ | ~new_n13450_);
  assign new_n13448_ = (~new_n13449_ | new_n6533_) & (new_n10000_ | new_n13478_ | ~new_n6354_);
  assign new_n13449_ = ~new_n8188_ & ~new_n6354_ & ~new_n13450_;
  assign new_n13450_ = ~new_n13451_ & new_n13475_;
  assign new_n13451_ = new_n13471_ & (~new_n13467_ | (~new_n13452_ & ~new_n13473_ & ~new_n13474_));
  assign new_n13452_ = ~new_n13464_ & ~new_n13462_ & (~new_n13466_ | ~new_n13461_ | new_n13453_);
  assign new_n13453_ = new_n13454_ & new_n13458_ & (new_n13456_ | ~\all_features[3109]  | ~\all_features[3110]  | ~\all_features[3111] );
  assign new_n13454_ = \all_features[3111]  & (\all_features[3110]  | (new_n13455_ & (\all_features[3106]  | \all_features[3107]  | \all_features[3105] )));
  assign new_n13455_ = \all_features[3108]  & \all_features[3109] ;
  assign new_n13456_ = ~\all_features[3107]  & ~\all_features[3108]  & (~\all_features[3106]  | new_n13457_);
  assign new_n13457_ = ~\all_features[3104]  & ~\all_features[3105] ;
  assign new_n13458_ = \all_features[3110]  & \all_features[3111]  & (\all_features[3108]  | \all_features[3109]  | new_n13459_ | ~new_n13460_);
  assign new_n13459_ = \all_features[3104]  & \all_features[3105] ;
  assign new_n13460_ = ~\all_features[3106]  & ~\all_features[3107] ;
  assign new_n13461_ = \all_features[3111]  & (\all_features[3110]  | (\all_features[3109]  & (\all_features[3108]  | ~new_n13460_ | ~new_n13457_)));
  assign new_n13462_ = ~\all_features[3111]  & (~\all_features[3110]  | ~new_n13459_ | ~new_n13455_ | ~new_n13463_);
  assign new_n13463_ = \all_features[3106]  & \all_features[3107] ;
  assign new_n13464_ = ~new_n13465_ & ~\all_features[3111] ;
  assign new_n13465_ = \all_features[3109]  & \all_features[3110]  & (\all_features[3108]  | (\all_features[3106]  & \all_features[3107]  & \all_features[3105] ));
  assign new_n13466_ = \all_features[3111]  & (\all_features[3109]  | \all_features[3110]  | \all_features[3108] );
  assign new_n13467_ = ~new_n13468_ & ~new_n13470_;
  assign new_n13468_ = new_n13469_ & (~\all_features[3107]  | ~new_n13455_ | (~\all_features[3106]  & ~new_n13459_));
  assign new_n13469_ = ~\all_features[3110]  & ~\all_features[3111] ;
  assign new_n13470_ = new_n13469_ & (~\all_features[3109]  | (~\all_features[3108]  & (~\all_features[3107]  | (~\all_features[3106]  & ~\all_features[3105] ))));
  assign new_n13471_ = ~new_n13472_ & (\all_features[3107]  | \all_features[3108]  | \all_features[3109]  | \all_features[3110]  | \all_features[3111] );
  assign new_n13472_ = ~\all_features[3109]  & new_n13469_ & ((~\all_features[3106]  & new_n13457_) | ~\all_features[3108]  | ~\all_features[3107] );
  assign new_n13473_ = ~\all_features[3111]  & (~\all_features[3110]  | (~\all_features[3108]  & ~\all_features[3109]  & ~new_n13463_));
  assign new_n13474_ = ~\all_features[3111]  & (~\all_features[3110]  | (~\all_features[3109]  & (new_n13457_ | ~new_n13463_ | ~\all_features[3108] )));
  assign new_n13475_ = ~new_n13467_ | ~new_n13471_;
  assign new_n13476_ = ~new_n13462_ & ~new_n13473_;
  assign new_n13478_ = new_n13479_ & new_n13505_;
  assign new_n13479_ = new_n13480_ & new_n13503_;
  assign new_n13480_ = new_n13498_ & ~new_n13502_ & ~new_n13481_ & ~new_n13501_;
  assign new_n13481_ = ~new_n13496_ & ~new_n13497_ & new_n13489_ & (~new_n13494_ | ~new_n13482_);
  assign new_n13482_ = new_n13488_ & new_n13483_ & new_n13485_;
  assign new_n13483_ = \all_features[4783]  & (\all_features[4782]  | (new_n13484_ & (\all_features[4778]  | \all_features[4779]  | \all_features[4777] )));
  assign new_n13484_ = \all_features[4780]  & \all_features[4781] ;
  assign new_n13485_ = \all_features[4782]  & \all_features[4783]  & (\all_features[4780]  | \all_features[4781]  | new_n13487_ | ~new_n13486_);
  assign new_n13486_ = ~\all_features[4778]  & ~\all_features[4779] ;
  assign new_n13487_ = \all_features[4776]  & \all_features[4777] ;
  assign new_n13488_ = \all_features[4783]  & (\all_features[4781]  | \all_features[4782]  | \all_features[4780] );
  assign new_n13489_ = ~new_n13490_ & ~new_n13492_;
  assign new_n13490_ = ~new_n13491_ & ~\all_features[4783] ;
  assign new_n13491_ = \all_features[4781]  & \all_features[4782]  & (\all_features[4780]  | (\all_features[4778]  & \all_features[4779]  & \all_features[4777] ));
  assign new_n13492_ = ~\all_features[4783]  & (~\all_features[4782]  | (~\all_features[4780]  & ~\all_features[4781]  & ~new_n13493_));
  assign new_n13493_ = \all_features[4778]  & \all_features[4779] ;
  assign new_n13494_ = \all_features[4783]  & (\all_features[4782]  | (\all_features[4781]  & (\all_features[4780]  | ~new_n13495_ | ~new_n13486_)));
  assign new_n13495_ = ~\all_features[4776]  & ~\all_features[4777] ;
  assign new_n13496_ = ~\all_features[4783]  & (~\all_features[4782]  | (~\all_features[4781]  & (new_n13495_ | ~new_n13493_ | ~\all_features[4780] )));
  assign new_n13497_ = ~\all_features[4783]  & (~\all_features[4782]  | ~new_n13484_ | ~new_n13487_ | ~new_n13493_);
  assign new_n13498_ = ~new_n13499_ & (\all_features[4779]  | \all_features[4780]  | \all_features[4781]  | \all_features[4782]  | \all_features[4783] );
  assign new_n13499_ = ~\all_features[4781]  & new_n13500_ & ((~\all_features[4778]  & new_n13495_) | ~\all_features[4780]  | ~\all_features[4779] );
  assign new_n13500_ = ~\all_features[4782]  & ~\all_features[4783] ;
  assign new_n13501_ = new_n13500_ & (~\all_features[4781]  | (~\all_features[4780]  & (~\all_features[4779]  | (~\all_features[4778]  & ~\all_features[4777] ))));
  assign new_n13502_ = new_n13500_ & (~\all_features[4779]  | ~new_n13484_ | (~\all_features[4778]  & ~new_n13487_));
  assign new_n13503_ = new_n13498_ & new_n13489_ & new_n13504_ & ~new_n13496_ & ~new_n13497_;
  assign new_n13504_ = ~new_n13501_ & ~new_n13502_;
  assign new_n13505_ = new_n13506_ & new_n13510_;
  assign new_n13506_ = new_n13498_ & (~new_n13504_ | (~new_n13507_ & ~new_n13492_ & ~new_n13496_));
  assign new_n13507_ = ~new_n13497_ & ~new_n13490_ & (~new_n13488_ | ~new_n13494_ | new_n13508_);
  assign new_n13508_ = new_n13483_ & new_n13485_ & (new_n13509_ | ~\all_features[4781]  | ~\all_features[4782]  | ~\all_features[4783] );
  assign new_n13509_ = ~\all_features[4779]  & ~\all_features[4780]  & (~\all_features[4778]  | new_n13495_);
  assign new_n13510_ = ~new_n13511_ & (\all_features[4779]  | \all_features[4780]  | \all_features[4781]  | \all_features[4782]  | \all_features[4783] );
  assign new_n13511_ = ~new_n13499_ & (new_n13501_ | (~new_n13502_ & (new_n13492_ | (~new_n13496_ & ~new_n13512_))));
  assign new_n13512_ = ~new_n13490_ & (new_n13497_ | (new_n13488_ & (~new_n13494_ | (~new_n13513_ & new_n13483_))));
  assign new_n13513_ = ~\all_features[4781]  & \all_features[4782]  & \all_features[4783]  & (\all_features[4780]  ? new_n13486_ : (new_n13487_ | ~new_n13486_));
  assign new_n13514_ = new_n13097_ & new_n10200_;
  assign new_n13515_ = new_n6354_ & new_n10000_ & (new_n13522_ ? new_n13523_ : new_n13516_);
  assign new_n13516_ = new_n13517_ & ~new_n13067_ & ~new_n13095_;
  assign new_n13517_ = ~new_n13090_ & ~new_n13518_;
  assign new_n13518_ = ~new_n13519_ & (\all_features[5027]  | \all_features[5028]  | \all_features[5029]  | \all_features[5030]  | \all_features[5031] );
  assign new_n13519_ = ~new_n13086_ & (new_n13088_ | (~new_n13089_ & (new_n13079_ | (~new_n13083_ & ~new_n13520_))));
  assign new_n13520_ = ~new_n13077_ & (new_n13084_ | (new_n13075_ & (~new_n13081_ | (~new_n13521_ & new_n13070_))));
  assign new_n13521_ = ~\all_features[5029]  & \all_features[5030]  & \all_features[5031]  & (\all_features[5028]  ? new_n13073_ : (new_n13074_ | ~new_n13073_));
  assign new_n13522_ = new_n8132_ & (new_n8129_ | new_n8099_);
  assign new_n13523_ = ~new_n13556_ & ~new_n13545_ & ~new_n13553_ & (new_n13551_ | (~new_n13550_ & ~new_n13524_));
  assign new_n13524_ = ~new_n13538_ & (new_n13540_ | (~new_n13541_ & (new_n13542_ | (~new_n13525_ & ~new_n13543_))));
  assign new_n13525_ = ~new_n13532_ & (~new_n13536_ | (new_n13526_ & (~new_n13535_ | (~new_n13537_ & new_n13529_))));
  assign new_n13526_ = \all_features[2191]  & (\all_features[2190]  | new_n13527_);
  assign new_n13527_ = \all_features[2189]  & (\all_features[2186]  | \all_features[2187]  | \all_features[2188]  | ~new_n13528_);
  assign new_n13528_ = ~\all_features[2184]  & ~\all_features[2185] ;
  assign new_n13529_ = \all_features[2191]  & ~new_n13530_ & \all_features[2190] ;
  assign new_n13530_ = ~\all_features[2189]  & ~\all_features[2188]  & ~\all_features[2187]  & ~new_n13531_ & ~\all_features[2186] ;
  assign new_n13531_ = \all_features[2184]  & \all_features[2185] ;
  assign new_n13532_ = ~\all_features[2191]  & (~\all_features[2190]  | ~new_n13531_ | ~new_n13533_ | ~new_n13534_);
  assign new_n13533_ = \all_features[2188]  & \all_features[2189] ;
  assign new_n13534_ = \all_features[2186]  & \all_features[2187] ;
  assign new_n13535_ = \all_features[2191]  & (\all_features[2190]  | (new_n13533_ & (\all_features[2186]  | \all_features[2187]  | \all_features[2185] )));
  assign new_n13536_ = \all_features[2191]  & (\all_features[2189]  | \all_features[2190]  | \all_features[2188] );
  assign new_n13537_ = \all_features[2190]  & \all_features[2191]  & (\all_features[2189]  | (\all_features[2188]  & (\all_features[2187]  | \all_features[2186] )));
  assign new_n13538_ = new_n13539_ & (~\all_features[2189]  | (~\all_features[2188]  & (~\all_features[2187]  | (~\all_features[2186]  & ~\all_features[2185] ))));
  assign new_n13539_ = ~\all_features[2190]  & ~\all_features[2191] ;
  assign new_n13540_ = new_n13539_ & (~\all_features[2187]  | ~new_n13533_ | (~\all_features[2186]  & ~new_n13531_));
  assign new_n13541_ = ~\all_features[2191]  & (~\all_features[2190]  | (~\all_features[2188]  & ~\all_features[2189]  & ~new_n13534_));
  assign new_n13542_ = ~\all_features[2191]  & (~\all_features[2190]  | (~\all_features[2189]  & (new_n13528_ | ~new_n13534_ | ~\all_features[2188] )));
  assign new_n13543_ = ~new_n13544_ & ~\all_features[2191] ;
  assign new_n13544_ = \all_features[2189]  & \all_features[2190]  & (\all_features[2188]  | (\all_features[2186]  & \all_features[2187]  & \all_features[2185] ));
  assign new_n13545_ = new_n13549_ & (~new_n13552_ | (~new_n13546_ & ~new_n13541_ & ~new_n13542_));
  assign new_n13546_ = ~new_n13532_ & ~new_n13543_ & (~new_n13536_ | new_n13547_ | ~new_n13526_);
  assign new_n13547_ = ~new_n13530_ & new_n13535_ & \all_features[2190]  & \all_features[2191]  & (~\all_features[2189]  | new_n13548_);
  assign new_n13548_ = ~\all_features[2187]  & ~\all_features[2188]  & (~\all_features[2186]  | new_n13528_);
  assign new_n13549_ = ~new_n13550_ & ~new_n13551_;
  assign new_n13550_ = ~\all_features[2189]  & new_n13539_ & ((~\all_features[2186]  & new_n13528_) | ~\all_features[2188]  | ~\all_features[2187] );
  assign new_n13551_ = ~\all_features[2191]  & ~\all_features[2190]  & ~\all_features[2189]  & ~\all_features[2187]  & ~\all_features[2188] ;
  assign new_n13552_ = ~new_n13538_ & ~new_n13540_;
  assign new_n13553_ = new_n13552_ & ~new_n13554_ & new_n13549_;
  assign new_n13554_ = new_n13555_ & (~new_n13535_ | ~new_n13536_ | ~new_n13529_ | ~new_n13526_);
  assign new_n13555_ = ~new_n13532_ & ~new_n13543_ & ~new_n13541_ & ~new_n13542_;
  assign new_n13556_ = new_n13557_ & new_n13549_ & ~new_n13538_ & ~new_n13543_;
  assign new_n13557_ = ~new_n13532_ & ~new_n13542_ & ~new_n13540_ & ~new_n13541_;
  assign new_n13558_ = (~new_n8188_ | new_n13559_ | new_n6354_) & (new_n10000_ | ~new_n13478_ | ~new_n13560_ | ~new_n6354_);
  assign new_n13559_ = new_n7304_ ? new_n8477_ : new_n13514_;
  assign new_n13560_ = ~new_n8927_ & (~new_n8924_ | new_n8893_);
  assign new_n13561_ = new_n13449_ & new_n6533_;
  assign \o[1]  = ~new_n13563_ ^ new_n13609_;
  assign new_n13563_ = new_n13564_ ? (~new_n13607_ ^ new_n13608_) : (new_n13607_ ^ new_n13608_);
  assign new_n13564_ = new_n13565_ ? (new_n13599_ ^ new_n13600_) : (~new_n13599_ ^ new_n13600_);
  assign new_n13565_ = new_n13566_ ? (new_n13585_ ^ new_n13586_) : (~new_n13585_ ^ new_n13586_);
  assign new_n13566_ = new_n13567_ ? (new_n13577_ ^ new_n13578_) : (~new_n13577_ ^ new_n13578_);
  assign new_n13567_ = new_n13568_ ? (new_n13572_ ^ new_n13573_) : (~new_n13572_ ^ new_n13573_);
  assign new_n13568_ = new_n13569_ ? (new_n13570_ ^ new_n13571_) : (~new_n13570_ ^ new_n13571_);
  assign new_n13569_ = ~new_n13561_ & new_n13446_;
  assign new_n13570_ = new_n6351_ & new_n6767_;
  assign new_n13571_ = new_n7263_ & new_n7551_ & (new_n7514_ | (~new_n7592_ & new_n7593_));
  assign new_n13572_ = (new_n6843_ & new_n7261_) | (new_n6350_ & (new_n6843_ | new_n7261_));
  assign new_n13573_ = new_n13574_ ? (new_n13575_ ^ new_n13576_) : (~new_n13575_ ^ new_n13576_);
  assign new_n13574_ = new_n6844_ & new_n7223_;
  assign new_n13575_ = new_n7952_ & new_n8348_;
  assign new_n13576_ = new_n13279_ & new_n13442_;
  assign new_n13577_ = (~new_n7594_ & new_n8538_) | (~new_n6349_ & (~new_n7594_ | new_n8538_));
  assign new_n13578_ = new_n13579_ ? (~new_n13583_ ^ new_n13584_) : (new_n13583_ ^ new_n13584_);
  assign new_n13579_ = new_n13580_ ? (new_n13581_ ^ new_n13582_) : (~new_n13581_ ^ new_n13582_);
  assign new_n13580_ = new_n7596_ & new_n7947_;
  assign new_n13581_ = new_n8351_ & new_n8536_;
  assign new_n13582_ = new_n12724_ & new_n12799_;
  assign new_n13583_ = (new_n7951_ & new_n8350_) | (new_n7595_ & (new_n7951_ | new_n8350_));
  assign new_n13584_ = (new_n9061_ & new_n9383_) | (new_n8814_ & (new_n9061_ | new_n9383_));
  assign new_n13585_ = (~new_n8812_ & new_n10163_) | (~new_n6348_ & (~new_n8812_ | new_n10163_));
  assign new_n13586_ = new_n13587_ ? (~new_n13597_ ^ new_n13598_) : (new_n13597_ ^ new_n13598_);
  assign new_n13587_ = new_n13588_ ? (new_n13592_ ^ new_n13593_) : (~new_n13592_ ^ new_n13593_);
  assign new_n13588_ = new_n13589_ ? (new_n13590_ ^ new_n13591_) : (~new_n13590_ ^ new_n13591_);
  assign new_n13589_ = new_n10164_ & new_n10369_;
  assign new_n13590_ = new_n12261_ & new_n12449_;
  assign new_n13591_ = new_n9062_ & new_n9381_;
  assign new_n13592_ = (new_n10641_ & new_n10835_) | (new_n10374_ & (new_n10641_ | new_n10835_));
  assign new_n13593_ = new_n13594_ ? (new_n13595_ ^ new_n13596_) : (~new_n13595_ ^ new_n13596_);
  assign new_n13594_ = new_n8815_ & new_n9059_;
  assign new_n13595_ = new_n12044_ & new_n12258_;
  assign new_n13596_ = ~new_n9607_ & new_n9384_;
  assign new_n13597_ = (~new_n11126_ & new_n11721_) | (new_n10373_ & (~new_n11126_ | new_n11721_));
  assign new_n13598_ = (new_n9608_ & new_n9895_) | (~new_n8813_ & (new_n9608_ | new_n9895_));
  assign new_n13599_ = (~new_n10371_ & new_n12451_) | (~new_n6347_ & (~new_n10371_ | new_n12451_));
  assign new_n13600_ = new_n13601_ ? (~new_n13602_ ^ new_n13606_) : (new_n13602_ ^ new_n13606_);
  assign new_n13601_ = (new_n12043_ & new_n12260_) | (~new_n10372_ & (new_n12043_ | new_n12260_));
  assign new_n13602_ = new_n13603_ ? (new_n13604_ ^ new_n13605_) : (~new_n13604_ ^ new_n13605_);
  assign new_n13603_ = (new_n11374_ & new_n11574_) | (new_n11127_ & (new_n11374_ | new_n11574_));
  assign new_n13604_ = new_n10375_ & new_n10638_;
  assign new_n13605_ = new_n11722_ & new_n12039_;
  assign new_n13606_ = (new_n12867_ & new_n13060_) | (new_n12838_ & (new_n12867_ | new_n13060_));
  assign new_n13607_ = (~new_n12722_ & new_n13278_) | (~new_n6346_ & (~new_n12722_ | new_n13278_));
  assign new_n13608_ = (~new_n12837_ & new_n13131_) | (new_n12723_ & (~new_n12837_ | new_n13131_));
  assign new_n13609_ = new_n6345_ & new_n13445_;
  assign \o[2]  = ~new_n13611_ ^ new_n13612_;
  assign new_n13611_ = ~new_n13563_ & new_n13609_;
  assign new_n13612_ = new_n13613_ ^ new_n13614_;
  assign new_n13613_ = (new_n13607_ & new_n13608_) | (~new_n13564_ & (new_n13607_ | new_n13608_));
  assign new_n13614_ = new_n13615_ ? (~new_n13616_ ^ new_n13636_) : (new_n13616_ ^ new_n13636_);
  assign new_n13615_ = (~new_n13600_ & new_n13599_) | (~new_n13565_ & (~new_n13600_ | new_n13599_));
  assign new_n13616_ = new_n13617_ ? (new_n13618_ ^ new_n13632_) : (~new_n13618_ ^ new_n13632_);
  assign new_n13617_ = (~new_n13586_ & new_n13585_) | (~new_n13566_ & (~new_n13586_ | new_n13585_));
  assign new_n13618_ = new_n13619_ ? (new_n13620_ ^ new_n13628_) : (~new_n13620_ ^ new_n13628_);
  assign new_n13619_ = (~new_n13578_ & new_n13577_) | (~new_n13567_ & (~new_n13578_ | new_n13577_));
  assign new_n13620_ = new_n13621_ ? (new_n13622_ ^ new_n13625_) : (~new_n13622_ ^ new_n13625_);
  assign new_n13621_ = (~new_n13573_ & new_n13572_) | (~new_n13568_ & (~new_n13573_ | new_n13572_));
  assign new_n13622_ = new_n13623_ ^ new_n13624_;
  assign new_n13623_ = (new_n13570_ & new_n13571_) | (new_n13569_ & (new_n13570_ | new_n13571_));
  assign new_n13624_ = new_n7262_ & new_n7551_;
  assign new_n13625_ = ~new_n13626_ ^ new_n13627_;
  assign new_n13626_ = (new_n13581_ & new_n13582_) | (new_n13580_ & (new_n13581_ | new_n13582_));
  assign new_n13627_ = (new_n13575_ & new_n13576_) | (new_n13574_ & (new_n13575_ | new_n13576_));
  assign new_n13628_ = new_n13629_ ? (new_n13630_ ^ new_n13631_) : (~new_n13630_ ^ new_n13631_);
  assign new_n13629_ = (new_n13583_ & new_n13584_) | (~new_n13579_ & (new_n13583_ | new_n13584_));
  assign new_n13630_ = (~new_n13593_ & new_n13592_) | (~new_n13588_ & (~new_n13593_ | new_n13592_));
  assign new_n13631_ = (new_n13595_ & new_n13596_) | (new_n13594_ & (new_n13595_ | new_n13596_));
  assign new_n13632_ = new_n13633_ ? (new_n13634_ ^ new_n13635_) : (~new_n13634_ ^ new_n13635_);
  assign new_n13633_ = (new_n13597_ & new_n13598_) | (~new_n13587_ & (new_n13597_ | new_n13598_));
  assign new_n13634_ = (new_n13604_ & new_n13605_) | (new_n13603_ & (new_n13604_ | new_n13605_));
  assign new_n13635_ = (new_n13590_ & new_n13591_) | (new_n13589_ & (new_n13590_ | new_n13591_));
  assign new_n13636_ = (~new_n13602_ & new_n13606_) | (new_n13601_ & (~new_n13602_ | new_n13606_));
  assign \o[3]  = ((new_n13638_ | new_n13639_) & (new_n13640_ ^ new_n13641_)) | (~new_n13638_ & ~new_n13639_ & (~new_n13640_ ^ new_n13641_));
  assign new_n13638_ = ~new_n13612_ & new_n13611_;
  assign new_n13639_ = ~new_n13614_ & new_n13613_;
  assign new_n13640_ = (~new_n13616_ & new_n13636_) | (new_n13615_ & (~new_n13616_ | new_n13636_));
  assign new_n13641_ = new_n13642_ ? (~new_n13643_ ^ new_n13650_) : (new_n13643_ ^ new_n13650_);
  assign new_n13642_ = (~new_n13618_ & ~new_n13632_) | (new_n13617_ & (~new_n13618_ | ~new_n13632_));
  assign new_n13643_ = new_n13644_ ? (~new_n13645_ ^ new_n13649_) : (new_n13645_ ^ new_n13649_);
  assign new_n13644_ = (~new_n13620_ & ~new_n13628_) | (new_n13619_ & (~new_n13620_ | ~new_n13628_));
  assign new_n13645_ = new_n13646_ ? (~new_n13647_ ^ new_n13648_) : (new_n13647_ ^ new_n13648_);
  assign new_n13646_ = (~new_n13622_ & ~new_n13625_) | (new_n13621_ & (~new_n13622_ | ~new_n13625_));
  assign new_n13647_ = ~new_n13623_ & ~new_n13624_;
  assign new_n13648_ = new_n13626_ & new_n13627_;
  assign new_n13649_ = (new_n13630_ & new_n13631_) | (new_n13629_ & (new_n13630_ | new_n13631_));
  assign new_n13650_ = (new_n13634_ & new_n13635_) | (new_n13633_ & (new_n13634_ | new_n13635_));
  assign \o[4]  = ~new_n13652_ ^ new_n13653_;
  assign new_n13652_ = (new_n13640_ | (~new_n13641_ & (new_n13639_ | new_n13638_))) & (new_n13639_ | new_n13638_ | ~new_n13641_);
  assign new_n13653_ = new_n13654_ ^ new_n13655_;
  assign new_n13654_ = (~new_n13643_ & new_n13650_) | (new_n13642_ & (~new_n13643_ | new_n13650_));
  assign new_n13655_ = ~new_n13656_ ^ new_n13657_;
  assign new_n13656_ = (~new_n13645_ & new_n13649_) | (new_n13644_ & (~new_n13645_ | new_n13649_));
  assign new_n13657_ = (~new_n13647_ & new_n13648_) | (new_n13646_ & (~new_n13647_ | new_n13648_));
  assign \o[5]  = (~new_n13661_ & (new_n13659_ | new_n13660_)) | (~new_n13659_ & ~new_n13660_ & new_n13661_);
  assign new_n13659_ = ~new_n13653_ & new_n13652_;
  assign new_n13660_ = ~new_n13655_ & new_n13654_;
  assign new_n13661_ = new_n13656_ & new_n13657_;
  assign \o[6]  = new_n13661_ & (new_n13660_ | new_n13659_);
  assign \o[7]  = new_n13664_ ? (new_n16895_ ^ new_n16953_) : (~new_n16895_ ^ new_n16953_);
  assign new_n13664_ = new_n13665_ ? (new_n16324_ ^ new_n16771_) : (~new_n16324_ ^ new_n16771_);
  assign new_n13665_ = new_n13666_ ? (new_n15400_ ^ new_n16149_) : (~new_n15400_ ^ new_n16149_);
  assign new_n13666_ = new_n13667_ ? (~new_n14869_ ^ new_n15350_) : (new_n14869_ ^ new_n15350_);
  assign new_n13667_ = new_n13668_ ? (new_n14284_ ^ new_n14613_) : (~new_n14284_ ^ new_n14613_);
  assign new_n13668_ = new_n13669_ ? (new_n13884_ ^ new_n14081_) : (~new_n13884_ ^ new_n14081_);
  assign new_n13669_ = ~new_n13670_ & new_n13847_;
  assign new_n13670_ = new_n13671_ & (~new_n13842_ | (~new_n13843_ & new_n13516_) | (~new_n13846_ & ~new_n13516_));
  assign new_n13671_ = new_n13672_ & (~new_n13803_ | (~new_n13806_ & new_n7600_) | (~new_n13807_ & ~new_n7600_));
  assign new_n13672_ = new_n12117_ | ((~new_n13734_ | ~new_n13774_ | new_n13766_) & (new_n13673_ | ~new_n13766_));
  assign new_n13673_ = new_n13674_ ? ~new_n8991_ : ~new_n13708_;
  assign new_n13674_ = ~new_n13675_ & ~new_n13707_;
  assign new_n13675_ = new_n13676_ & new_n13703_;
  assign new_n13676_ = ~new_n13677_ & (\all_features[3507]  | \all_features[3508]  | \all_features[3509]  | \all_features[3510]  | \all_features[3511] );
  assign new_n13677_ = new_n13678_ & (new_n13700_ | (~new_n13698_ & (new_n13691_ | (~new_n13701_ & ~new_n13693_))));
  assign new_n13678_ = ~new_n13695_ & ~new_n13699_ & ~new_n13697_ & (new_n13700_ | new_n13698_ | new_n13679_);
  assign new_n13679_ = ~new_n13691_ & ~new_n13693_ & (~new_n13689_ | (~new_n13680_ & new_n13683_));
  assign new_n13680_ = \all_features[3511]  & \all_features[3510]  & ~new_n13681_ & \all_features[3509] ;
  assign new_n13681_ = ~\all_features[3507]  & ~\all_features[3508]  & (~\all_features[3506]  | new_n13682_);
  assign new_n13682_ = ~\all_features[3504]  & ~\all_features[3505] ;
  assign new_n13683_ = new_n13684_ & \all_features[3510]  & \all_features[3511]  & (~new_n13688_ | ~new_n13687_ | new_n13686_);
  assign new_n13684_ = \all_features[3511]  & (\all_features[3510]  | (new_n13685_ & (\all_features[3506]  | \all_features[3507]  | \all_features[3505] )));
  assign new_n13685_ = \all_features[3508]  & \all_features[3509] ;
  assign new_n13686_ = \all_features[3504]  & \all_features[3505] ;
  assign new_n13687_ = ~\all_features[3508]  & ~\all_features[3509] ;
  assign new_n13688_ = ~\all_features[3506]  & ~\all_features[3507] ;
  assign new_n13689_ = \all_features[3511]  & (\all_features[3510]  | (~new_n13687_ & new_n13690_));
  assign new_n13690_ = \all_features[3509]  & (\all_features[3508]  | ~new_n13688_ | ~new_n13682_);
  assign new_n13691_ = ~new_n13692_ & ~\all_features[3511] ;
  assign new_n13692_ = \all_features[3509]  & \all_features[3510]  & (\all_features[3508]  | (\all_features[3506]  & \all_features[3507]  & \all_features[3505] ));
  assign new_n13693_ = ~\all_features[3511]  & (~\all_features[3510]  | ~new_n13694_ | ~new_n13686_ | ~new_n13685_);
  assign new_n13694_ = \all_features[3506]  & \all_features[3507] ;
  assign new_n13695_ = new_n13696_ & (~\all_features[3509]  | (~\all_features[3508]  & (~\all_features[3507]  | (~\all_features[3506]  & ~\all_features[3505] ))));
  assign new_n13696_ = ~\all_features[3510]  & ~\all_features[3511] ;
  assign new_n13697_ = ~\all_features[3509]  & new_n13696_ & ((~\all_features[3506]  & new_n13682_) | ~\all_features[3508]  | ~\all_features[3507] );
  assign new_n13698_ = ~\all_features[3511]  & (~\all_features[3510]  | (~\all_features[3509]  & (new_n13682_ | ~new_n13694_ | ~\all_features[3508] )));
  assign new_n13699_ = new_n13696_ & (~\all_features[3507]  | ~new_n13685_ | (~\all_features[3506]  & ~new_n13686_));
  assign new_n13700_ = ~\all_features[3511]  & (~\all_features[3510]  | (~new_n13694_ & new_n13687_));
  assign new_n13701_ = \all_features[3511]  & ((~new_n13702_ & \all_features[3510]  & new_n13684_) | (~new_n13687_ & ((~new_n13702_ & new_n13684_) | (~new_n13690_ & ~\all_features[3510] ))));
  assign new_n13702_ = ~\all_features[3509]  & \all_features[3510]  & \all_features[3511]  & (\all_features[3508]  ? new_n13688_ : (new_n13686_ | ~new_n13688_));
  assign new_n13703_ = new_n13706_ & ~new_n13699_ & ~new_n13704_ & ~new_n13695_;
  assign new_n13704_ = ~new_n13691_ & ~new_n13698_ & new_n13705_ & (~new_n13689_ | ~new_n13683_);
  assign new_n13705_ = ~new_n13693_ & ~new_n13700_;
  assign new_n13706_ = ~new_n13697_ & (\all_features[3507]  | \all_features[3508]  | \all_features[3509]  | \all_features[3510]  | \all_features[3511] );
  assign new_n13707_ = new_n13705_ & new_n13706_ & ~new_n13699_ & ~new_n13698_ & ~new_n13691_ & ~new_n13695_;
  assign new_n13708_ = new_n13709_ & new_n13733_;
  assign new_n13709_ = new_n13727_ & (~new_n13720_ | (new_n13716_ & new_n13710_));
  assign new_n13710_ = \all_features[4671]  & \all_features[4670]  & ~new_n13711_ & new_n13714_;
  assign new_n13711_ = new_n13712_ & ~\all_features[4669]  & ~new_n13713_ & ~\all_features[4668] ;
  assign new_n13712_ = ~\all_features[4666]  & ~\all_features[4667] ;
  assign new_n13713_ = \all_features[4664]  & \all_features[4665] ;
  assign new_n13714_ = \all_features[4671]  & (\all_features[4670]  | (new_n13715_ & (\all_features[4666]  | \all_features[4667]  | \all_features[4665] )));
  assign new_n13715_ = \all_features[4668]  & \all_features[4669] ;
  assign new_n13716_ = new_n13717_ & new_n13719_;
  assign new_n13717_ = \all_features[4671]  & (\all_features[4670]  | (\all_features[4669]  & (\all_features[4668]  | ~new_n13718_ | ~new_n13712_)));
  assign new_n13718_ = ~\all_features[4664]  & ~\all_features[4665] ;
  assign new_n13719_ = \all_features[4671]  & (\all_features[4669]  | \all_features[4670]  | \all_features[4668] );
  assign new_n13720_ = ~new_n13726_ & ~new_n13725_ & ~new_n13721_ & ~new_n13723_;
  assign new_n13721_ = ~\all_features[4671]  & (~\all_features[4670]  | (~\all_features[4669]  & (new_n13718_ | ~new_n13722_ | ~\all_features[4668] )));
  assign new_n13722_ = \all_features[4666]  & \all_features[4667] ;
  assign new_n13723_ = ~new_n13724_ & ~\all_features[4671] ;
  assign new_n13724_ = \all_features[4669]  & \all_features[4670]  & (\all_features[4668]  | (\all_features[4666]  & \all_features[4667]  & \all_features[4665] ));
  assign new_n13725_ = ~\all_features[4671]  & (~\all_features[4670]  | ~new_n13713_ | ~new_n13715_ | ~new_n13722_);
  assign new_n13726_ = ~\all_features[4671]  & (~\all_features[4670]  | (~\all_features[4668]  & ~\all_features[4669]  & ~new_n13722_));
  assign new_n13727_ = ~new_n13732_ & ~new_n13731_ & ~new_n13728_ & ~new_n13730_;
  assign new_n13728_ = new_n13729_ & (~\all_features[4669]  | (~\all_features[4668]  & (~\all_features[4667]  | (~\all_features[4666]  & ~\all_features[4665] ))));
  assign new_n13729_ = ~\all_features[4670]  & ~\all_features[4671] ;
  assign new_n13730_ = new_n13729_ & (~\all_features[4667]  | ~new_n13715_ | (~\all_features[4666]  & ~new_n13713_));
  assign new_n13731_ = ~\all_features[4669]  & new_n13729_ & ((~\all_features[4666]  & new_n13718_) | ~\all_features[4668]  | ~\all_features[4667] );
  assign new_n13732_ = ~\all_features[4671]  & ~\all_features[4670]  & ~\all_features[4669]  & ~\all_features[4667]  & ~\all_features[4668] ;
  assign new_n13733_ = new_n13720_ & new_n13727_;
  assign new_n13734_ = new_n13735_ & new_n13765_;
  assign new_n13735_ = new_n13736_ & new_n13758_;
  assign new_n13736_ = new_n13753_ & ~new_n13757_ & ~new_n13737_ & ~new_n13756_;
  assign new_n13737_ = new_n13738_ & (~new_n13751_ | ~new_n13752_ | ~new_n13748_ | ~new_n13750_);
  assign new_n13738_ = ~new_n13747_ & ~new_n13744_ & ~new_n13739_ & ~new_n13742_;
  assign new_n13739_ = ~\all_features[5551]  & (~\all_features[5550]  | (~\all_features[5549]  & (new_n13740_ | ~new_n13741_ | ~\all_features[5548] )));
  assign new_n13740_ = ~\all_features[5544]  & ~\all_features[5545] ;
  assign new_n13741_ = \all_features[5546]  & \all_features[5547] ;
  assign new_n13742_ = ~new_n13743_ & ~\all_features[5551] ;
  assign new_n13743_ = \all_features[5549]  & \all_features[5550]  & (\all_features[5548]  | (\all_features[5546]  & \all_features[5547]  & \all_features[5545] ));
  assign new_n13744_ = ~\all_features[5551]  & (~\all_features[5550]  | ~new_n13745_ | ~new_n13746_ | ~new_n13741_);
  assign new_n13745_ = \all_features[5548]  & \all_features[5549] ;
  assign new_n13746_ = \all_features[5544]  & \all_features[5545] ;
  assign new_n13747_ = ~\all_features[5551]  & (~\all_features[5550]  | (~\all_features[5548]  & ~\all_features[5549]  & ~new_n13741_));
  assign new_n13748_ = \all_features[5551]  & (\all_features[5550]  | (\all_features[5549]  & (\all_features[5548]  | ~new_n13740_ | ~new_n13749_)));
  assign new_n13749_ = ~\all_features[5546]  & ~\all_features[5547] ;
  assign new_n13750_ = \all_features[5551]  & (\all_features[5550]  | (new_n13745_ & (\all_features[5546]  | \all_features[5547]  | \all_features[5545] )));
  assign new_n13751_ = \all_features[5550]  & \all_features[5551]  & (\all_features[5548]  | \all_features[5549]  | new_n13746_ | ~new_n13749_);
  assign new_n13752_ = \all_features[5551]  & (\all_features[5549]  | \all_features[5550]  | \all_features[5548] );
  assign new_n13753_ = ~new_n13754_ & (\all_features[5547]  | \all_features[5548]  | \all_features[5549]  | \all_features[5550]  | \all_features[5551] );
  assign new_n13754_ = ~\all_features[5549]  & new_n13755_ & ((~\all_features[5546]  & new_n13740_) | ~\all_features[5548]  | ~\all_features[5547] );
  assign new_n13755_ = ~\all_features[5550]  & ~\all_features[5551] ;
  assign new_n13756_ = new_n13755_ & (~\all_features[5549]  | (~\all_features[5548]  & (~\all_features[5547]  | (~\all_features[5546]  & ~\all_features[5545] ))));
  assign new_n13757_ = new_n13755_ & (~\all_features[5547]  | ~new_n13745_ | (~\all_features[5546]  & ~new_n13746_));
  assign new_n13758_ = new_n13753_ & (~new_n13764_ | (~new_n13759_ & new_n13763_));
  assign new_n13759_ = new_n13762_ & ((~new_n13760_ & new_n13750_ & new_n13751_) | ~new_n13752_ | ~new_n13748_);
  assign new_n13760_ = \all_features[5551]  & \all_features[5550]  & ~new_n13761_ & \all_features[5549] ;
  assign new_n13761_ = ~\all_features[5547]  & ~\all_features[5548]  & (~\all_features[5546]  | new_n13740_);
  assign new_n13762_ = ~new_n13742_ & ~new_n13744_;
  assign new_n13763_ = ~new_n13739_ & ~new_n13747_;
  assign new_n13764_ = ~new_n13756_ & ~new_n13757_;
  assign new_n13765_ = new_n13764_ & new_n13763_ & new_n13753_ & new_n13762_;
  assign new_n13766_ = new_n13767_ & new_n13773_;
  assign new_n13767_ = new_n11297_ & new_n13768_;
  assign new_n13768_ = ~new_n11293_ & (new_n11290_ | (~new_n11296_ & (new_n11295_ | (~new_n11283_ & ~new_n13769_))));
  assign new_n13769_ = ~new_n11285_ & (new_n11286_ | (~new_n11288_ & (~new_n13772_ | new_n13770_)));
  assign new_n13770_ = \all_features[3911]  & ((~new_n13771_ & ~\all_features[3909]  & \all_features[3910] ) | (~new_n11280_ & (\all_features[3910]  | (~new_n11277_ & \all_features[3909] ))));
  assign new_n13771_ = (~\all_features[3906]  & ~\all_features[3907]  & ~\all_features[3908]  & (~\all_features[3905]  | ~\all_features[3904] )) | (\all_features[3908]  & (\all_features[3906]  | \all_features[3907] ));
  assign new_n13772_ = \all_features[3911]  & (\all_features[3909]  | \all_features[3910]  | \all_features[3908] );
  assign new_n13773_ = new_n11274_ & new_n11301_;
  assign new_n13774_ = ~new_n13775_ & new_n13799_;
  assign new_n13775_ = new_n13791_ & (~new_n13794_ | (~new_n13776_ & ~new_n13797_ & ~new_n13798_));
  assign new_n13776_ = ~new_n13787_ & ~new_n13789_ & (~new_n13777_ | (~new_n13780_ & new_n13782_));
  assign new_n13777_ = \all_features[1087]  & (\all_features[1086]  | (~new_n13778_ & \all_features[1085] ));
  assign new_n13778_ = new_n13779_ & ~\all_features[1084]  & ~\all_features[1082]  & ~\all_features[1083] ;
  assign new_n13779_ = ~\all_features[1080]  & ~\all_features[1081] ;
  assign new_n13780_ = \all_features[1087]  & \all_features[1086]  & ~new_n13781_ & \all_features[1085] ;
  assign new_n13781_ = ~\all_features[1083]  & ~\all_features[1084]  & (~\all_features[1082]  | new_n13779_);
  assign new_n13782_ = \all_features[1087]  & \all_features[1086]  & ~new_n13785_ & new_n13783_;
  assign new_n13783_ = \all_features[1087]  & (\all_features[1086]  | (new_n13784_ & (\all_features[1082]  | \all_features[1083]  | \all_features[1081] )));
  assign new_n13784_ = \all_features[1084]  & \all_features[1085] ;
  assign new_n13785_ = ~\all_features[1085]  & ~\all_features[1084]  & ~\all_features[1083]  & ~new_n13786_ & ~\all_features[1082] ;
  assign new_n13786_ = \all_features[1080]  & \all_features[1081] ;
  assign new_n13787_ = ~\all_features[1087]  & (~\all_features[1086]  | ~new_n13784_ | ~new_n13786_ | ~new_n13788_);
  assign new_n13788_ = \all_features[1082]  & \all_features[1083] ;
  assign new_n13789_ = ~new_n13790_ & ~\all_features[1087] ;
  assign new_n13790_ = \all_features[1085]  & \all_features[1086]  & (\all_features[1084]  | (\all_features[1082]  & \all_features[1083]  & \all_features[1081] ));
  assign new_n13791_ = ~new_n13792_ & (\all_features[1083]  | \all_features[1084]  | \all_features[1085]  | \all_features[1086]  | \all_features[1087] );
  assign new_n13792_ = ~\all_features[1085]  & new_n13793_ & ((~\all_features[1082]  & new_n13779_) | ~\all_features[1084]  | ~\all_features[1083] );
  assign new_n13793_ = ~\all_features[1086]  & ~\all_features[1087] ;
  assign new_n13794_ = ~new_n13795_ & ~new_n13796_;
  assign new_n13795_ = new_n13793_ & (~\all_features[1085]  | (~\all_features[1084]  & (~\all_features[1083]  | (~\all_features[1082]  & ~\all_features[1081] ))));
  assign new_n13796_ = new_n13793_ & (~\all_features[1083]  | ~new_n13784_ | (~new_n13786_ & ~\all_features[1082] ));
  assign new_n13797_ = ~\all_features[1087]  & (~\all_features[1086]  | (~\all_features[1084]  & ~\all_features[1085]  & ~new_n13788_));
  assign new_n13798_ = ~\all_features[1087]  & (~\all_features[1086]  | (~\all_features[1085]  & (new_n13779_ | ~new_n13788_ | ~\all_features[1084] )));
  assign new_n13799_ = ~new_n13800_ & (new_n13802_ | ~new_n13791_ | ~new_n13794_);
  assign new_n13800_ = new_n13801_ & new_n13791_ & ~new_n13789_ & ~new_n13795_;
  assign new_n13801_ = ~new_n13796_ & ~new_n13798_ & ~new_n13787_ & ~new_n13797_;
  assign new_n13802_ = ~new_n13787_ & ~new_n13789_ & ~new_n13797_ & ~new_n13798_ & (~new_n13782_ | ~new_n13777_);
  assign new_n13803_ = ~new_n13804_ & new_n12117_;
  assign new_n13804_ = new_n6908_ & new_n13805_ & new_n6886_;
  assign new_n13805_ = new_n6910_ & new_n6914_;
  assign new_n13806_ = new_n10976_ & new_n13319_;
  assign new_n13807_ = new_n13808_ & new_n13837_;
  assign new_n13808_ = new_n13809_ & new_n13830_;
  assign new_n13809_ = ~new_n13810_ & (\all_features[2363]  | \all_features[2364]  | \all_features[2365]  | \all_features[2366]  | \all_features[2367] );
  assign new_n13810_ = ~new_n13826_ & (new_n13824_ | (~new_n13828_ & (new_n13829_ | (~new_n13827_ & ~new_n13811_))));
  assign new_n13811_ = ~new_n13812_ & (new_n13814_ | (new_n13823_ & (~new_n13818_ | (~new_n13822_ & new_n13821_))));
  assign new_n13812_ = ~new_n13813_ & ~\all_features[2367] ;
  assign new_n13813_ = \all_features[2365]  & \all_features[2366]  & (\all_features[2364]  | (\all_features[2362]  & \all_features[2363]  & \all_features[2361] ));
  assign new_n13814_ = ~\all_features[2367]  & (~\all_features[2366]  | ~new_n13815_ | ~new_n13816_ | ~new_n13817_);
  assign new_n13815_ = \all_features[2362]  & \all_features[2363] ;
  assign new_n13816_ = \all_features[2360]  & \all_features[2361] ;
  assign new_n13817_ = \all_features[2364]  & \all_features[2365] ;
  assign new_n13818_ = \all_features[2367]  & (\all_features[2366]  | (\all_features[2365]  & (\all_features[2364]  | ~new_n13820_ | ~new_n13819_)));
  assign new_n13819_ = ~\all_features[2360]  & ~\all_features[2361] ;
  assign new_n13820_ = ~\all_features[2362]  & ~\all_features[2363] ;
  assign new_n13821_ = \all_features[2367]  & (\all_features[2366]  | (new_n13817_ & (\all_features[2362]  | \all_features[2363]  | \all_features[2361] )));
  assign new_n13822_ = ~\all_features[2365]  & \all_features[2366]  & \all_features[2367]  & (\all_features[2364]  ? new_n13820_ : (new_n13816_ | ~new_n13820_));
  assign new_n13823_ = \all_features[2367]  & (\all_features[2365]  | \all_features[2366]  | \all_features[2364] );
  assign new_n13824_ = new_n13825_ & (~\all_features[2365]  | (~\all_features[2364]  & (~\all_features[2363]  | (~\all_features[2362]  & ~\all_features[2361] ))));
  assign new_n13825_ = ~\all_features[2366]  & ~\all_features[2367] ;
  assign new_n13826_ = ~\all_features[2365]  & new_n13825_ & ((~\all_features[2362]  & new_n13819_) | ~\all_features[2364]  | ~\all_features[2363] );
  assign new_n13827_ = ~\all_features[2367]  & (~\all_features[2366]  | (~\all_features[2365]  & (new_n13819_ | ~new_n13815_ | ~\all_features[2364] )));
  assign new_n13828_ = new_n13825_ & (~\all_features[2363]  | ~new_n13817_ | (~\all_features[2362]  & ~new_n13816_));
  assign new_n13829_ = ~\all_features[2367]  & (~\all_features[2366]  | (~\all_features[2364]  & ~\all_features[2365]  & ~new_n13815_));
  assign new_n13830_ = new_n13835_ & (~new_n13836_ | (~new_n13831_ & ~new_n13827_ & ~new_n13829_));
  assign new_n13831_ = ~new_n13812_ & ~new_n13814_ & (~new_n13823_ | ~new_n13818_ | new_n13832_);
  assign new_n13832_ = new_n13821_ & new_n13833_ & (new_n13834_ | ~\all_features[2365]  | ~\all_features[2366]  | ~\all_features[2367] );
  assign new_n13833_ = \all_features[2366]  & \all_features[2367]  & (\all_features[2364]  | \all_features[2365]  | new_n13816_ | ~new_n13820_);
  assign new_n13834_ = ~\all_features[2363]  & ~\all_features[2364]  & (~\all_features[2362]  | new_n13819_);
  assign new_n13835_ = ~new_n13826_ & (\all_features[2363]  | \all_features[2364]  | \all_features[2365]  | \all_features[2366]  | \all_features[2367] );
  assign new_n13836_ = ~new_n13824_ & ~new_n13828_;
  assign new_n13837_ = new_n13838_ & new_n13840_;
  assign new_n13838_ = new_n13839_ & new_n13835_ & ~new_n13828_ & ~new_n13827_ & ~new_n13812_ & ~new_n13824_;
  assign new_n13839_ = ~new_n13814_ & ~new_n13829_;
  assign new_n13840_ = new_n13835_ & new_n13836_ & (new_n13841_ | new_n13812_ | new_n13827_ | ~new_n13839_);
  assign new_n13841_ = new_n13823_ & new_n13833_ & new_n13818_ & new_n13821_;
  assign new_n13842_ = new_n12117_ & new_n13804_;
  assign new_n13843_ = new_n13844_ & new_n13845_;
  assign new_n13844_ = ~new_n11379_ & ~new_n11403_;
  assign new_n13845_ = ~new_n11407_ & ~new_n11409_;
  assign new_n13846_ = new_n13838_ & (new_n13840_ | new_n13808_);
  assign new_n13847_ = new_n13848_ & (~new_n13842_ | (new_n13843_ & new_n13516_) | (new_n13846_ & ~new_n13516_));
  assign new_n13848_ = new_n13849_ & (~new_n13803_ | (new_n13806_ & new_n7600_) | (new_n13807_ & ~new_n7600_));
  assign new_n13849_ = new_n12117_ | (new_n13766_ ? ~new_n13673_ : (new_n13774_ ? new_n13734_ : new_n13850_));
  assign new_n13850_ = new_n13882_ & new_n13880_ & new_n13851_ & new_n13873_;
  assign new_n13851_ = ~new_n13872_ & (new_n13867_ | (~new_n13869_ & (new_n13870_ | (~new_n13852_ & ~new_n13871_))));
  assign new_n13852_ = ~new_n13859_ & (new_n13862_ | (~new_n13864_ & (~new_n13866_ | (~new_n13853_ & new_n13865_))));
  assign new_n13853_ = new_n13854_ & (\all_features[4757]  | ~new_n13858_ | (~new_n13856_ & ~\all_features[4756]  & new_n13857_) | (\all_features[4756]  & ~new_n13857_));
  assign new_n13854_ = \all_features[4759]  & (\all_features[4758]  | (new_n13855_ & (\all_features[4754]  | \all_features[4755]  | \all_features[4753] )));
  assign new_n13855_ = \all_features[4756]  & \all_features[4757] ;
  assign new_n13856_ = \all_features[4752]  & \all_features[4753] ;
  assign new_n13857_ = ~\all_features[4754]  & ~\all_features[4755] ;
  assign new_n13858_ = \all_features[4758]  & \all_features[4759] ;
  assign new_n13859_ = ~\all_features[4759]  & (~\all_features[4758]  | (~\all_features[4757]  & (new_n13860_ | ~new_n13861_ | ~\all_features[4756] )));
  assign new_n13860_ = ~\all_features[4752]  & ~\all_features[4753] ;
  assign new_n13861_ = \all_features[4754]  & \all_features[4755] ;
  assign new_n13862_ = ~new_n13863_ & ~\all_features[4759] ;
  assign new_n13863_ = \all_features[4757]  & \all_features[4758]  & (\all_features[4756]  | (\all_features[4754]  & \all_features[4755]  & \all_features[4753] ));
  assign new_n13864_ = ~\all_features[4759]  & (~\all_features[4758]  | ~new_n13856_ | ~new_n13855_ | ~new_n13861_);
  assign new_n13865_ = \all_features[4759]  & (\all_features[4758]  | (\all_features[4757]  & (\all_features[4756]  | ~new_n13857_ | ~new_n13860_)));
  assign new_n13866_ = \all_features[4759]  & (\all_features[4757]  | \all_features[4758]  | \all_features[4756] );
  assign new_n13867_ = ~\all_features[4757]  & new_n13868_ & ((~\all_features[4754]  & new_n13860_) | ~\all_features[4756]  | ~\all_features[4755] );
  assign new_n13868_ = ~\all_features[4758]  & ~\all_features[4759] ;
  assign new_n13869_ = new_n13868_ & (~\all_features[4757]  | (~\all_features[4756]  & (~\all_features[4755]  | (~\all_features[4754]  & ~\all_features[4753] ))));
  assign new_n13870_ = new_n13868_ & (~\all_features[4755]  | ~new_n13855_ | (~\all_features[4754]  & ~new_n13856_));
  assign new_n13871_ = ~\all_features[4759]  & (~\all_features[4758]  | (~\all_features[4756]  & ~\all_features[4757]  & ~new_n13861_));
  assign new_n13872_ = ~\all_features[4759]  & ~\all_features[4758]  & ~\all_features[4757]  & ~\all_features[4755]  & ~\all_features[4756] ;
  assign new_n13873_ = ~new_n13867_ & ~new_n13872_ & (~new_n13878_ | (~new_n13874_ & new_n13879_));
  assign new_n13874_ = new_n13875_ & ((~new_n13877_ & new_n13876_ & new_n13854_) | ~new_n13866_ | ~new_n13865_);
  assign new_n13875_ = ~new_n13862_ & ~new_n13864_;
  assign new_n13876_ = new_n13858_ & (new_n13856_ | \all_features[4756]  | \all_features[4757]  | ~new_n13857_);
  assign new_n13877_ = new_n13858_ & \all_features[4757]  & ((~new_n13860_ & \all_features[4754] ) | \all_features[4756]  | \all_features[4755] );
  assign new_n13878_ = ~new_n13869_ & ~new_n13870_;
  assign new_n13879_ = ~new_n13871_ & ~new_n13859_;
  assign new_n13880_ = ~new_n13872_ & ~new_n13870_ & ~new_n13869_ & ~new_n13881_ & ~new_n13867_;
  assign new_n13881_ = new_n13879_ & new_n13875_ & (~new_n13876_ | ~new_n13866_ | ~new_n13865_ | ~new_n13854_);
  assign new_n13882_ = new_n13883_ & new_n13878_ & ~new_n13862_ & ~new_n13859_ & ~new_n13867_ & ~new_n13871_;
  assign new_n13883_ = ~new_n13864_ & ~new_n13872_;
  assign new_n13884_ = new_n13885_ & ~new_n14012_ & ~new_n14043_;
  assign new_n13885_ = new_n13886_ & (new_n13976_ | ~new_n12849_ | ~new_n13922_ | (new_n14008_ & new_n13982_));
  assign new_n13886_ = (new_n13922_ | new_n13887_ | new_n6460_ | ~new_n12849_) & (new_n13943_ | new_n13941_ | new_n12849_);
  assign new_n13887_ = new_n13888_ & ~new_n13918_ & ~new_n13921_;
  assign new_n13888_ = ~new_n13889_ & ~new_n13909_;
  assign new_n13889_ = (new_n13890_ | (~new_n13908_ & ~\all_features[1677]  & new_n13905_)) & (\all_features[1675]  | \all_features[1676]  | \all_features[1677]  | ~new_n13905_);
  assign new_n13890_ = ~new_n13904_ & (new_n13906_ | (~new_n13891_ & ~new_n13907_));
  assign new_n13891_ = ~new_n13898_ & (new_n13900_ | (~new_n13902_ & (~new_n13903_ | new_n13892_)));
  assign new_n13892_ = \all_features[1679]  & ((~new_n13897_ & ~\all_features[1677]  & \all_features[1678] ) | (~new_n13895_ & (\all_features[1678]  | (~new_n13893_ & \all_features[1677] ))));
  assign new_n13893_ = new_n13894_ & ~\all_features[1676]  & ~\all_features[1674]  & ~\all_features[1675] ;
  assign new_n13894_ = ~\all_features[1672]  & ~\all_features[1673] ;
  assign new_n13895_ = \all_features[1679]  & (\all_features[1678]  | (new_n13896_ & (\all_features[1674]  | \all_features[1675]  | \all_features[1673] )));
  assign new_n13896_ = \all_features[1676]  & \all_features[1677] ;
  assign new_n13897_ = (~\all_features[1674]  & ~\all_features[1675]  & ~\all_features[1676]  & (~\all_features[1673]  | ~\all_features[1672] )) | (\all_features[1676]  & (\all_features[1674]  | \all_features[1675] ));
  assign new_n13898_ = ~\all_features[1679]  & (~\all_features[1678]  | (~\all_features[1677]  & (new_n13894_ | ~new_n13899_ | ~\all_features[1676] )));
  assign new_n13899_ = \all_features[1674]  & \all_features[1675] ;
  assign new_n13900_ = ~new_n13901_ & ~\all_features[1679] ;
  assign new_n13901_ = \all_features[1677]  & \all_features[1678]  & (\all_features[1676]  | (\all_features[1674]  & \all_features[1675]  & \all_features[1673] ));
  assign new_n13902_ = ~\all_features[1679]  & (~new_n13899_ | ~\all_features[1672]  | ~\all_features[1673]  | ~\all_features[1678]  | ~new_n13896_);
  assign new_n13903_ = \all_features[1679]  & (\all_features[1677]  | \all_features[1678]  | \all_features[1676] );
  assign new_n13904_ = new_n13905_ & (~\all_features[1677]  | (~\all_features[1676]  & (~\all_features[1675]  | (~\all_features[1674]  & ~\all_features[1673] ))));
  assign new_n13905_ = ~\all_features[1678]  & ~\all_features[1679] ;
  assign new_n13906_ = new_n13905_ & (~new_n13896_ | ~\all_features[1675]  | (~\all_features[1674]  & (~\all_features[1672]  | ~\all_features[1673] )));
  assign new_n13907_ = ~\all_features[1679]  & (~\all_features[1678]  | (~\all_features[1676]  & ~\all_features[1677]  & ~new_n13899_));
  assign new_n13908_ = \all_features[1675]  & \all_features[1676]  & (\all_features[1674]  | ~new_n13894_);
  assign new_n13909_ = new_n13916_ & (~new_n13917_ | (~new_n13910_ & ~new_n13907_ & ~new_n13898_));
  assign new_n13910_ = ~new_n13900_ & ~new_n13902_ & (~new_n13911_ | (~new_n13914_ & new_n13912_));
  assign new_n13911_ = \all_features[1679]  & (\all_features[1678]  | (~new_n13893_ & \all_features[1677] ));
  assign new_n13912_ = \all_features[1679]  & \all_features[1678]  & ~new_n13913_ & new_n13895_;
  assign new_n13913_ = ~\all_features[1674]  & ~\all_features[1675]  & ~\all_features[1676]  & ~\all_features[1677]  & (~\all_features[1673]  | ~\all_features[1672] );
  assign new_n13914_ = \all_features[1679]  & \all_features[1678]  & ~new_n13915_ & \all_features[1677] ;
  assign new_n13915_ = ~\all_features[1675]  & ~\all_features[1676]  & (~\all_features[1674]  | new_n13894_);
  assign new_n13916_ = \all_features[1677]  | ~new_n13905_ | (new_n13908_ & (\all_features[1675]  | \all_features[1676] ));
  assign new_n13917_ = ~new_n13904_ & ~new_n13906_;
  assign new_n13918_ = new_n13919_ & (~new_n13920_ | (new_n13911_ & new_n13912_));
  assign new_n13919_ = new_n13916_ & new_n13917_;
  assign new_n13920_ = ~new_n13902_ & ~new_n13900_ & ~new_n13907_ & ~new_n13898_;
  assign new_n13921_ = new_n13919_ & new_n13920_;
  assign new_n13922_ = new_n13923_ & new_n13932_;
  assign new_n13923_ = ~new_n13924_ & ~new_n10682_;
  assign new_n13924_ = ~new_n10695_ & ~new_n10691_ & ~new_n10687_ & ~new_n13925_ & ~new_n10697_;
  assign new_n13925_ = ~new_n10696_ & ~new_n10698_ & ~new_n10692_ & ~new_n10683_ & ~new_n13926_;
  assign new_n13926_ = new_n13931_ & new_n13930_ & new_n13927_ & new_n13929_;
  assign new_n13927_ = \all_features[2383]  & (\all_features[2382]  | (\all_features[2381]  & (\all_features[2380]  | ~new_n13928_ | ~new_n10685_)));
  assign new_n13928_ = ~\all_features[2378]  & ~\all_features[2379] ;
  assign new_n13929_ = \all_features[2383]  & (\all_features[2382]  | (new_n10690_ & (\all_features[2378]  | \all_features[2379]  | \all_features[2377] )));
  assign new_n13930_ = \all_features[2382]  & \all_features[2383]  & (\all_features[2380]  | \all_features[2381]  | new_n10689_ | ~new_n13928_);
  assign new_n13931_ = \all_features[2383]  & (\all_features[2381]  | \all_features[2382]  | \all_features[2380] );
  assign new_n13932_ = ~new_n13933_ & ~new_n13937_;
  assign new_n13933_ = ~new_n10695_ & ~new_n10697_ & (~new_n10686_ | (~new_n10683_ & ~new_n13934_ & ~new_n10696_));
  assign new_n13934_ = ~new_n10692_ & ~new_n10698_ & (~new_n13931_ | ~new_n13927_ | new_n13935_);
  assign new_n13935_ = new_n13929_ & new_n13930_ & (new_n13936_ | ~\all_features[2381]  | ~\all_features[2382]  | ~\all_features[2383] );
  assign new_n13936_ = ~\all_features[2379]  & ~\all_features[2380]  & (~\all_features[2378]  | new_n10685_);
  assign new_n13937_ = ~new_n13938_ & ~new_n10695_;
  assign new_n13938_ = ~new_n10697_ & (new_n10691_ | (~new_n10687_ & (new_n10696_ | (~new_n10683_ & ~new_n13939_))));
  assign new_n13939_ = ~new_n10692_ & (new_n10698_ | (new_n13931_ & (~new_n13927_ | (~new_n13940_ & new_n13929_))));
  assign new_n13940_ = ~\all_features[2381]  & \all_features[2382]  & \all_features[2383]  & (\all_features[2380]  ? new_n13928_ : (new_n10689_ | ~new_n13928_));
  assign new_n13941_ = ~new_n13942_ & new_n10677_;
  assign new_n13942_ = ~new_n10670_ & ~new_n10679_;
  assign new_n13943_ = new_n13971_ & new_n13974_ & new_n13964_ & (new_n13970_ | new_n13944_);
  assign new_n13944_ = ~new_n13957_ & (new_n13959_ | (~new_n13960_ & (new_n13961_ | (~new_n13945_ & ~new_n13962_))));
  assign new_n13945_ = ~new_n13949_ & (~new_n13955_ | (new_n13946_ & (~new_n13954_ | (~new_n13956_ & new_n13952_))));
  assign new_n13946_ = \all_features[4975]  & (\all_features[4974]  | new_n13947_);
  assign new_n13947_ = \all_features[4973]  & (\all_features[4970]  | \all_features[4971]  | \all_features[4972]  | ~new_n13948_);
  assign new_n13948_ = ~\all_features[4968]  & ~\all_features[4969] ;
  assign new_n13949_ = ~\all_features[4975]  & (~new_n13951_ | ~\all_features[4968]  | ~\all_features[4969]  | ~\all_features[4974]  | ~new_n13950_);
  assign new_n13950_ = \all_features[4972]  & \all_features[4973] ;
  assign new_n13951_ = \all_features[4970]  & \all_features[4971] ;
  assign new_n13952_ = \all_features[4975]  & ~new_n13953_ & \all_features[4974] ;
  assign new_n13953_ = ~\all_features[4970]  & ~\all_features[4971]  & ~\all_features[4972]  & ~\all_features[4973]  & (~\all_features[4969]  | ~\all_features[4968] );
  assign new_n13954_ = \all_features[4975]  & (\all_features[4974]  | (new_n13950_ & (\all_features[4970]  | \all_features[4971]  | \all_features[4969] )));
  assign new_n13955_ = \all_features[4975]  & (\all_features[4973]  | \all_features[4974]  | \all_features[4972] );
  assign new_n13956_ = \all_features[4974]  & \all_features[4975]  & (\all_features[4973]  | (\all_features[4972]  & (\all_features[4971]  | \all_features[4970] )));
  assign new_n13957_ = new_n13958_ & (~\all_features[4973]  | (~\all_features[4972]  & (~\all_features[4971]  | (~\all_features[4970]  & ~\all_features[4969] ))));
  assign new_n13958_ = ~\all_features[4974]  & ~\all_features[4975] ;
  assign new_n13959_ = new_n13958_ & (~new_n13950_ | ~\all_features[4971]  | (~\all_features[4970]  & (~\all_features[4968]  | ~\all_features[4969] )));
  assign new_n13960_ = ~\all_features[4975]  & (~\all_features[4974]  | (~\all_features[4972]  & ~\all_features[4973]  & ~new_n13951_));
  assign new_n13961_ = ~\all_features[4975]  & (~\all_features[4974]  | (~\all_features[4973]  & (new_n13948_ | ~new_n13951_ | ~\all_features[4972] )));
  assign new_n13962_ = ~new_n13963_ & ~\all_features[4975] ;
  assign new_n13963_ = \all_features[4973]  & \all_features[4974]  & (\all_features[4972]  | (\all_features[4970]  & \all_features[4971]  & \all_features[4969] ));
  assign new_n13964_ = new_n13969_ & (~new_n13968_ | (~new_n13965_ & ~new_n13960_ & ~new_n13961_));
  assign new_n13965_ = ~new_n13949_ & ~new_n13962_ & (~new_n13955_ | new_n13966_ | ~new_n13946_);
  assign new_n13966_ = ~new_n13953_ & new_n13954_ & \all_features[4974]  & \all_features[4975]  & (~\all_features[4973]  | new_n13967_);
  assign new_n13967_ = ~\all_features[4971]  & ~\all_features[4972]  & (~\all_features[4970]  | new_n13948_);
  assign new_n13968_ = ~new_n13957_ & ~new_n13959_;
  assign new_n13969_ = ~new_n13970_ & (\all_features[4971]  | \all_features[4972]  | \all_features[4973]  | \all_features[4974]  | \all_features[4975] );
  assign new_n13970_ = ~\all_features[4973]  & new_n13958_ & ((~\all_features[4970]  & new_n13948_) | ~\all_features[4972]  | ~\all_features[4971] );
  assign new_n13971_ = new_n13968_ & new_n13969_ & (new_n13972_ | new_n13961_ | new_n13949_ | ~new_n13973_);
  assign new_n13972_ = new_n13955_ & new_n13954_ & new_n13946_ & new_n13952_;
  assign new_n13973_ = ~new_n13960_ & ~new_n13962_;
  assign new_n13974_ = new_n13975_ & (\all_features[4971]  | \all_features[4972]  | \all_features[4973]  | \all_features[4974]  | \all_features[4975] );
  assign new_n13975_ = new_n13969_ & new_n13968_ & new_n13973_ & ~new_n13961_ & ~new_n13949_;
  assign new_n13976_ = new_n13169_ & new_n13977_;
  assign new_n13977_ = ~new_n13197_ & ~new_n13978_;
  assign new_n13978_ = ~new_n13190_ & (new_n13189_ | new_n13979_);
  assign new_n13979_ = ~new_n13185_ & (new_n13187_ | (~new_n13180_ & (new_n13181_ | (~new_n13173_ & ~new_n13980_))));
  assign new_n13980_ = ~new_n13175_ & (~new_n13195_ | (new_n13194_ & (~new_n13191_ | (~new_n13981_ & new_n13192_))));
  assign new_n13981_ = \all_features[3894]  & \all_features[3895]  & (\all_features[3893]  | (~new_n13193_ & \all_features[3892] ));
  assign new_n13982_ = new_n13983_ & new_n14006_;
  assign new_n13983_ = new_n14001_ & ~new_n14005_ & ~new_n13984_ & ~new_n14004_;
  assign new_n13984_ = ~new_n13999_ & ~new_n14000_ & new_n13992_ & (~new_n13997_ | ~new_n13985_);
  assign new_n13985_ = new_n13991_ & new_n13986_ & new_n13988_;
  assign new_n13986_ = \all_features[4631]  & (\all_features[4630]  | (new_n13987_ & (\all_features[4626]  | \all_features[4627]  | \all_features[4625] )));
  assign new_n13987_ = \all_features[4628]  & \all_features[4629] ;
  assign new_n13988_ = \all_features[4630]  & \all_features[4631]  & (\all_features[4628]  | \all_features[4629]  | new_n13990_ | ~new_n13989_);
  assign new_n13989_ = ~\all_features[4626]  & ~\all_features[4627] ;
  assign new_n13990_ = \all_features[4624]  & \all_features[4625] ;
  assign new_n13991_ = \all_features[4631]  & (\all_features[4629]  | \all_features[4630]  | \all_features[4628] );
  assign new_n13992_ = ~new_n13993_ & ~new_n13995_;
  assign new_n13993_ = ~new_n13994_ & ~\all_features[4631] ;
  assign new_n13994_ = \all_features[4629]  & \all_features[4630]  & (\all_features[4628]  | (\all_features[4626]  & \all_features[4627]  & \all_features[4625] ));
  assign new_n13995_ = ~\all_features[4631]  & (~\all_features[4630]  | (~\all_features[4628]  & ~\all_features[4629]  & ~new_n13996_));
  assign new_n13996_ = \all_features[4626]  & \all_features[4627] ;
  assign new_n13997_ = \all_features[4631]  & (\all_features[4630]  | (\all_features[4629]  & (\all_features[4628]  | ~new_n13998_ | ~new_n13989_)));
  assign new_n13998_ = ~\all_features[4624]  & ~\all_features[4625] ;
  assign new_n13999_ = ~\all_features[4631]  & (~\all_features[4630]  | (~\all_features[4629]  & (new_n13998_ | ~new_n13996_ | ~\all_features[4628] )));
  assign new_n14000_ = ~\all_features[4631]  & (~\all_features[4630]  | ~new_n13987_ | ~new_n13990_ | ~new_n13996_);
  assign new_n14001_ = ~new_n14002_ & (\all_features[4627]  | \all_features[4628]  | \all_features[4629]  | \all_features[4630]  | \all_features[4631] );
  assign new_n14002_ = ~\all_features[4629]  & new_n14003_ & ((~\all_features[4626]  & new_n13998_) | ~\all_features[4628]  | ~\all_features[4627] );
  assign new_n14003_ = ~\all_features[4630]  & ~\all_features[4631] ;
  assign new_n14004_ = new_n14003_ & (~\all_features[4629]  | (~\all_features[4628]  & (~\all_features[4627]  | (~\all_features[4626]  & ~\all_features[4625] ))));
  assign new_n14005_ = new_n14003_ & (~\all_features[4627]  | ~new_n13987_ | (~\all_features[4626]  & ~new_n13990_));
  assign new_n14006_ = new_n14001_ & new_n13992_ & new_n14007_ & ~new_n13999_ & ~new_n14000_;
  assign new_n14007_ = ~new_n14004_ & ~new_n14005_;
  assign new_n14008_ = new_n14001_ & (~new_n14007_ | (~new_n14009_ & ~new_n13995_ & ~new_n13999_));
  assign new_n14009_ = ~new_n14000_ & ~new_n13993_ & (~new_n13991_ | ~new_n13997_ | new_n14010_);
  assign new_n14010_ = new_n13986_ & new_n13988_ & (new_n14011_ | ~\all_features[4629]  | ~\all_features[4630]  | ~\all_features[4631] );
  assign new_n14011_ = ~\all_features[4627]  & ~\all_features[4628]  & (~\all_features[4626]  | new_n13998_);
  assign new_n14012_ = new_n12849_ & ((~new_n6603_ & new_n13976_ & new_n13922_) | (~new_n14013_ & new_n13887_ & ~new_n13922_));
  assign new_n14013_ = ~new_n14014_ & new_n14038_;
  assign new_n14014_ = new_n14035_ & (~new_n14029_ | (~new_n14015_ & ~new_n14033_ & ~new_n14037_));
  assign new_n14015_ = ~new_n14026_ & ~new_n14025_ & (~new_n14028_ | ~new_n14024_ | new_n14016_);
  assign new_n14016_ = new_n14017_ & new_n14019_ & (new_n14022_ | ~\all_features[2557]  | ~\all_features[2558]  | ~\all_features[2559] );
  assign new_n14017_ = \all_features[2559]  & (\all_features[2558]  | (new_n14018_ & (\all_features[2554]  | \all_features[2555]  | \all_features[2553] )));
  assign new_n14018_ = \all_features[2556]  & \all_features[2557] ;
  assign new_n14019_ = \all_features[2558]  & \all_features[2559]  & (\all_features[2556]  | \all_features[2557]  | new_n14020_ | ~new_n14021_);
  assign new_n14020_ = \all_features[2552]  & \all_features[2553] ;
  assign new_n14021_ = ~\all_features[2554]  & ~\all_features[2555] ;
  assign new_n14022_ = ~\all_features[2555]  & ~\all_features[2556]  & (~\all_features[2554]  | new_n14023_);
  assign new_n14023_ = ~\all_features[2552]  & ~\all_features[2553] ;
  assign new_n14024_ = \all_features[2559]  & (\all_features[2558]  | (\all_features[2557]  & (\all_features[2556]  | ~new_n14023_ | ~new_n14021_)));
  assign new_n14025_ = ~\all_features[2559]  & (~new_n14018_ | ~\all_features[2554]  | ~\all_features[2555]  | ~\all_features[2558]  | ~new_n14020_);
  assign new_n14026_ = ~new_n14027_ & ~\all_features[2559] ;
  assign new_n14027_ = \all_features[2557]  & \all_features[2558]  & (\all_features[2556]  | (\all_features[2554]  & \all_features[2555]  & \all_features[2553] ));
  assign new_n14028_ = \all_features[2559]  & (\all_features[2557]  | \all_features[2558]  | \all_features[2556] );
  assign new_n14029_ = ~new_n14030_ & ~new_n14032_;
  assign new_n14030_ = new_n14031_ & (~\all_features[2555]  | ~new_n14018_ | (~\all_features[2554]  & ~new_n14020_));
  assign new_n14031_ = ~\all_features[2558]  & ~\all_features[2559] ;
  assign new_n14032_ = new_n14031_ & (~\all_features[2557]  | (~\all_features[2556]  & (~\all_features[2555]  | (~\all_features[2554]  & ~\all_features[2553] ))));
  assign new_n14033_ = ~\all_features[2559]  & (~\all_features[2558]  | new_n14034_);
  assign new_n14034_ = ~\all_features[2557]  & (new_n14023_ | ~\all_features[2555]  | ~\all_features[2556]  | ~\all_features[2554] );
  assign new_n14035_ = ~new_n14036_ & (\all_features[2555]  | \all_features[2556]  | \all_features[2557]  | \all_features[2558]  | \all_features[2559] );
  assign new_n14036_ = ~\all_features[2557]  & new_n14031_ & ((~\all_features[2554]  & new_n14023_) | ~\all_features[2556]  | ~\all_features[2555] );
  assign new_n14037_ = ~\all_features[2559]  & (~\all_features[2558]  | (~\all_features[2557]  & ~\all_features[2556]  & (~\all_features[2555]  | ~\all_features[2554] )));
  assign new_n14038_ = ~new_n14039_ & ~new_n14042_;
  assign new_n14039_ = new_n14029_ & new_n14035_ & (new_n14033_ | new_n14040_ | new_n14025_ | ~new_n14041_);
  assign new_n14040_ = new_n14028_ & new_n14024_ & new_n14017_ & new_n14019_;
  assign new_n14041_ = ~new_n14026_ & ~new_n14037_;
  assign new_n14042_ = new_n14029_ & new_n14041_ & new_n14035_ & ~new_n14033_ & ~new_n14025_;
  assign new_n14043_ = ~new_n12849_ & new_n13941_ & (new_n14044_ ? ~new_n12755_ : (~new_n14072_ | ~new_n14046_));
  assign new_n14044_ = new_n14045_ & ~new_n12978_ & ~new_n12980_;
  assign new_n14045_ = ~new_n12947_ & ~new_n12968_;
  assign new_n14046_ = new_n14047_ & new_n14070_;
  assign new_n14047_ = new_n14065_ & ~new_n14069_ & ~new_n14048_ & ~new_n14068_;
  assign new_n14048_ = ~new_n14063_ & ~new_n14064_ & new_n14056_ & (~new_n14061_ | ~new_n14049_);
  assign new_n14049_ = new_n14055_ & new_n14050_ & new_n14052_;
  assign new_n14050_ = \all_features[5487]  & (\all_features[5486]  | (new_n14051_ & (\all_features[5482]  | \all_features[5483]  | \all_features[5481] )));
  assign new_n14051_ = \all_features[5484]  & \all_features[5485] ;
  assign new_n14052_ = \all_features[5486]  & \all_features[5487]  & (\all_features[5484]  | \all_features[5485]  | new_n14054_ | ~new_n14053_);
  assign new_n14053_ = ~\all_features[5482]  & ~\all_features[5483] ;
  assign new_n14054_ = \all_features[5480]  & \all_features[5481] ;
  assign new_n14055_ = \all_features[5487]  & (\all_features[5485]  | \all_features[5486]  | \all_features[5484] );
  assign new_n14056_ = ~new_n14057_ & ~new_n14059_;
  assign new_n14057_ = ~new_n14058_ & ~\all_features[5487] ;
  assign new_n14058_ = \all_features[5485]  & \all_features[5486]  & (\all_features[5484]  | (\all_features[5482]  & \all_features[5483]  & \all_features[5481] ));
  assign new_n14059_ = ~\all_features[5487]  & (~\all_features[5486]  | (~\all_features[5484]  & ~\all_features[5485]  & ~new_n14060_));
  assign new_n14060_ = \all_features[5482]  & \all_features[5483] ;
  assign new_n14061_ = \all_features[5487]  & (\all_features[5486]  | (\all_features[5485]  & (\all_features[5484]  | ~new_n14062_ | ~new_n14053_)));
  assign new_n14062_ = ~\all_features[5480]  & ~\all_features[5481] ;
  assign new_n14063_ = ~\all_features[5487]  & (~\all_features[5486]  | (~\all_features[5485]  & (new_n14062_ | ~new_n14060_ | ~\all_features[5484] )));
  assign new_n14064_ = ~\all_features[5487]  & (~\all_features[5486]  | ~new_n14051_ | ~new_n14054_ | ~new_n14060_);
  assign new_n14065_ = ~new_n14066_ & (\all_features[5483]  | \all_features[5484]  | \all_features[5485]  | \all_features[5486]  | \all_features[5487] );
  assign new_n14066_ = ~\all_features[5485]  & new_n14067_ & ((~\all_features[5482]  & new_n14062_) | ~\all_features[5484]  | ~\all_features[5483] );
  assign new_n14067_ = ~\all_features[5486]  & ~\all_features[5487] ;
  assign new_n14068_ = new_n14067_ & (~\all_features[5485]  | (~\all_features[5484]  & (~\all_features[5483]  | (~\all_features[5482]  & ~\all_features[5481] ))));
  assign new_n14069_ = new_n14067_ & (~\all_features[5483]  | ~new_n14051_ | (~\all_features[5482]  & ~new_n14054_));
  assign new_n14070_ = new_n14065_ & new_n14056_ & new_n14071_ & ~new_n14063_ & ~new_n14064_;
  assign new_n14071_ = ~new_n14068_ & ~new_n14069_;
  assign new_n14072_ = new_n14073_ & new_n14077_;
  assign new_n14073_ = ~new_n14074_ & (\all_features[5483]  | \all_features[5484]  | \all_features[5485]  | \all_features[5486]  | \all_features[5487] );
  assign new_n14074_ = ~new_n14066_ & (new_n14068_ | (~new_n14069_ & (new_n14059_ | (~new_n14063_ & ~new_n14075_))));
  assign new_n14075_ = ~new_n14057_ & (new_n14064_ | (new_n14055_ & (~new_n14061_ | (~new_n14076_ & new_n14050_))));
  assign new_n14076_ = ~\all_features[5485]  & \all_features[5486]  & \all_features[5487]  & (\all_features[5484]  ? new_n14053_ : (new_n14054_ | ~new_n14053_));
  assign new_n14077_ = new_n14065_ & (~new_n14071_ | (~new_n14078_ & ~new_n14059_ & ~new_n14063_));
  assign new_n14078_ = ~new_n14064_ & ~new_n14057_ & (~new_n14055_ | ~new_n14061_ | new_n14079_);
  assign new_n14079_ = new_n14050_ & new_n14052_ & (new_n14080_ | ~\all_features[5485]  | ~\all_features[5486]  | ~\all_features[5487] );
  assign new_n14080_ = ~\all_features[5483]  & ~\all_features[5484]  & (~\all_features[5482]  | new_n14062_);
  assign new_n14081_ = (new_n14161_ & new_n14278_ & (~new_n14275_ | new_n13887_)) | (new_n14082_ & ~new_n14241_ & ~new_n14278_);
  assign new_n14082_ = new_n14158_ ? new_n14083_ : (~new_n14124_ | (~new_n10999_ & new_n14160_));
  assign new_n14083_ = (new_n14119_ & new_n13887_ & (new_n14122_ | ~new_n14090_)) | (new_n14084_ & ~new_n13887_);
  assign new_n14084_ = new_n11977_ & new_n14085_;
  assign new_n14085_ = ~new_n12002_ & ~new_n14086_;
  assign new_n14086_ = ~new_n14087_ & (\all_features[3459]  | \all_features[3460]  | \all_features[3461]  | \all_features[3462]  | \all_features[3463] );
  assign new_n14087_ = ~new_n11995_ & (new_n11993_ | (~new_n11991_ & (new_n11988_ | (~new_n11980_ & ~new_n14088_))));
  assign new_n14088_ = ~new_n11986_ & (new_n11983_ | (new_n12000_ & (~new_n11999_ | (~new_n14089_ & new_n11996_))));
  assign new_n14089_ = ~\all_features[3461]  & \all_features[3462]  & \all_features[3463]  & (\all_features[3460]  ? new_n11998_ : (new_n11984_ | ~new_n11998_));
  assign new_n14090_ = ~new_n14091_ & ~new_n14115_;
  assign new_n14091_ = new_n14112_ & (~new_n14106_ | (~new_n14092_ & ~new_n14110_ & ~new_n14114_));
  assign new_n14092_ = ~new_n14103_ & ~new_n14102_ & (~new_n14105_ | ~new_n14101_ | new_n14093_);
  assign new_n14093_ = new_n14094_ & new_n14096_ & (new_n14099_ | ~\all_features[1941]  | ~\all_features[1942]  | ~\all_features[1943] );
  assign new_n14094_ = \all_features[1943]  & (\all_features[1942]  | (new_n14095_ & (\all_features[1938]  | \all_features[1939]  | \all_features[1937] )));
  assign new_n14095_ = \all_features[1940]  & \all_features[1941] ;
  assign new_n14096_ = \all_features[1942]  & \all_features[1943]  & (\all_features[1940]  | \all_features[1941]  | new_n14097_ | ~new_n14098_);
  assign new_n14097_ = \all_features[1936]  & \all_features[1937] ;
  assign new_n14098_ = ~\all_features[1938]  & ~\all_features[1939] ;
  assign new_n14099_ = ~\all_features[1939]  & ~\all_features[1940]  & (~\all_features[1938]  | new_n14100_);
  assign new_n14100_ = ~\all_features[1936]  & ~\all_features[1937] ;
  assign new_n14101_ = \all_features[1943]  & (\all_features[1942]  | (\all_features[1941]  & (\all_features[1940]  | ~new_n14100_ | ~new_n14098_)));
  assign new_n14102_ = ~\all_features[1943]  & (~new_n14095_ | ~\all_features[1938]  | ~\all_features[1939]  | ~\all_features[1942]  | ~new_n14097_);
  assign new_n14103_ = ~new_n14104_ & ~\all_features[1943] ;
  assign new_n14104_ = \all_features[1941]  & \all_features[1942]  & (\all_features[1940]  | (\all_features[1938]  & \all_features[1939]  & \all_features[1937] ));
  assign new_n14105_ = \all_features[1943]  & (\all_features[1941]  | \all_features[1942]  | \all_features[1940] );
  assign new_n14106_ = ~new_n14107_ & ~new_n14109_;
  assign new_n14107_ = new_n14108_ & (~\all_features[1939]  | ~new_n14095_ | (~\all_features[1938]  & ~new_n14097_));
  assign new_n14108_ = ~\all_features[1942]  & ~\all_features[1943] ;
  assign new_n14109_ = new_n14108_ & (~\all_features[1941]  | (~\all_features[1940]  & (~\all_features[1939]  | (~\all_features[1938]  & ~\all_features[1937] ))));
  assign new_n14110_ = ~\all_features[1943]  & (~\all_features[1942]  | new_n14111_);
  assign new_n14111_ = ~\all_features[1941]  & (new_n14100_ | ~\all_features[1939]  | ~\all_features[1940]  | ~\all_features[1938] );
  assign new_n14112_ = ~new_n14113_ & (\all_features[1939]  | \all_features[1940]  | \all_features[1941]  | \all_features[1942]  | \all_features[1943] );
  assign new_n14113_ = ~\all_features[1941]  & new_n14108_ & ((~\all_features[1938]  & new_n14100_) | ~\all_features[1940]  | ~\all_features[1939] );
  assign new_n14114_ = ~\all_features[1943]  & (~\all_features[1942]  | (~\all_features[1941]  & ~\all_features[1940]  & (~\all_features[1939]  | ~\all_features[1938] )));
  assign new_n14115_ = ~new_n14116_ & (\all_features[1939]  | \all_features[1940]  | \all_features[1941]  | \all_features[1942]  | \all_features[1943] );
  assign new_n14116_ = ~new_n14113_ & (new_n14109_ | (~new_n14107_ & (new_n14114_ | (~new_n14110_ & ~new_n14117_))));
  assign new_n14117_ = ~new_n14103_ & (new_n14102_ | (new_n14105_ & (~new_n14101_ | (~new_n14118_ & new_n14094_))));
  assign new_n14118_ = ~\all_features[1941]  & \all_features[1942]  & \all_features[1943]  & (\all_features[1940]  ? new_n14098_ : (new_n14097_ | ~new_n14098_));
  assign new_n14119_ = new_n14106_ & new_n14121_ & new_n14120_ & ~new_n14110_ & ~new_n14113_;
  assign new_n14120_ = ~new_n14102_ & (\all_features[1939]  | \all_features[1940]  | \all_features[1941]  | \all_features[1942]  | \all_features[1943] );
  assign new_n14121_ = ~new_n14103_ & ~new_n14114_;
  assign new_n14122_ = new_n14106_ & new_n14112_ & (new_n14110_ | new_n14123_ | new_n14102_ | ~new_n14121_);
  assign new_n14123_ = new_n14105_ & new_n14101_ & new_n14094_ & new_n14096_;
  assign new_n14124_ = new_n14156_ & new_n14125_ & new_n14154_;
  assign new_n14125_ = new_n14126_ & new_n14147_;
  assign new_n14126_ = ~new_n14127_ & (\all_features[4827]  | \all_features[4828]  | \all_features[4829]  | \all_features[4830]  | \all_features[4831] );
  assign new_n14127_ = ~new_n14143_ & (new_n14141_ | (~new_n14145_ & (new_n14146_ | (~new_n14144_ & ~new_n14128_))));
  assign new_n14128_ = ~new_n14129_ & (new_n14131_ | (new_n14140_ & (~new_n14135_ | (~new_n14139_ & new_n14138_))));
  assign new_n14129_ = ~new_n14130_ & ~\all_features[4831] ;
  assign new_n14130_ = \all_features[4829]  & \all_features[4830]  & (\all_features[4828]  | (\all_features[4826]  & \all_features[4827]  & \all_features[4825] ));
  assign new_n14131_ = ~\all_features[4831]  & (~\all_features[4830]  | ~new_n14132_ | ~new_n14133_ | ~new_n14134_);
  assign new_n14132_ = \all_features[4826]  & \all_features[4827] ;
  assign new_n14133_ = \all_features[4824]  & \all_features[4825] ;
  assign new_n14134_ = \all_features[4828]  & \all_features[4829] ;
  assign new_n14135_ = \all_features[4831]  & (\all_features[4830]  | (\all_features[4829]  & (\all_features[4828]  | ~new_n14137_ | ~new_n14136_)));
  assign new_n14136_ = ~\all_features[4824]  & ~\all_features[4825] ;
  assign new_n14137_ = ~\all_features[4826]  & ~\all_features[4827] ;
  assign new_n14138_ = \all_features[4831]  & (\all_features[4830]  | (new_n14134_ & (\all_features[4826]  | \all_features[4827]  | \all_features[4825] )));
  assign new_n14139_ = ~\all_features[4829]  & \all_features[4830]  & \all_features[4831]  & (\all_features[4828]  ? new_n14137_ : (new_n14133_ | ~new_n14137_));
  assign new_n14140_ = \all_features[4831]  & (\all_features[4829]  | \all_features[4830]  | \all_features[4828] );
  assign new_n14141_ = new_n14142_ & (~\all_features[4829]  | (~\all_features[4828]  & (~\all_features[4827]  | (~\all_features[4826]  & ~\all_features[4825] ))));
  assign new_n14142_ = ~\all_features[4830]  & ~\all_features[4831] ;
  assign new_n14143_ = ~\all_features[4829]  & new_n14142_ & ((~\all_features[4826]  & new_n14136_) | ~\all_features[4828]  | ~\all_features[4827] );
  assign new_n14144_ = ~\all_features[4831]  & (~\all_features[4830]  | (~\all_features[4829]  & (new_n14136_ | ~new_n14132_ | ~\all_features[4828] )));
  assign new_n14145_ = new_n14142_ & (~\all_features[4827]  | ~new_n14134_ | (~\all_features[4826]  & ~new_n14133_));
  assign new_n14146_ = ~\all_features[4831]  & (~\all_features[4830]  | (~\all_features[4828]  & ~\all_features[4829]  & ~new_n14132_));
  assign new_n14147_ = new_n14152_ & (~new_n14153_ | (~new_n14148_ & ~new_n14144_ & ~new_n14146_));
  assign new_n14148_ = ~new_n14129_ & ~new_n14131_ & (~new_n14140_ | ~new_n14135_ | new_n14149_);
  assign new_n14149_ = new_n14138_ & new_n14150_ & (new_n14151_ | ~\all_features[4829]  | ~\all_features[4830]  | ~\all_features[4831] );
  assign new_n14150_ = \all_features[4830]  & \all_features[4831]  & (\all_features[4828]  | \all_features[4829]  | new_n14133_ | ~new_n14137_);
  assign new_n14151_ = ~\all_features[4827]  & ~\all_features[4828]  & (~\all_features[4826]  | new_n14136_);
  assign new_n14152_ = ~new_n14143_ & (\all_features[4827]  | \all_features[4828]  | \all_features[4829]  | \all_features[4830]  | \all_features[4831] );
  assign new_n14153_ = ~new_n14141_ & ~new_n14145_;
  assign new_n14154_ = new_n14155_ & new_n14152_ & ~new_n14145_ & ~new_n14144_ & ~new_n14129_ & ~new_n14141_;
  assign new_n14155_ = ~new_n14131_ & ~new_n14146_;
  assign new_n14156_ = new_n14152_ & new_n14153_ & (new_n14157_ | new_n14129_ | new_n14144_ | ~new_n14155_);
  assign new_n14157_ = new_n14140_ & new_n14150_ & new_n14135_ & new_n14138_;
  assign new_n14158_ = new_n14159_ & new_n6521_;
  assign new_n14159_ = new_n6529_ & new_n6532_;
  assign new_n14160_ = ~new_n10977_ & ~new_n13324_;
  assign new_n14161_ = (~new_n6384_ | ~new_n13887_ | new_n14162_) & (new_n14181_ | ~new_n14162_ | (~new_n14237_ & new_n14211_));
  assign new_n14162_ = new_n14163_ & new_n14172_;
  assign new_n14163_ = ~new_n14164_ & ~new_n12354_;
  assign new_n14164_ = ~new_n12367_ & ~new_n12363_ & ~new_n12359_ & ~new_n14165_ & ~new_n12369_;
  assign new_n14165_ = ~new_n12368_ & ~new_n12370_ & ~new_n12364_ & ~new_n12355_ & ~new_n14166_;
  assign new_n14166_ = new_n14171_ & new_n14170_ & new_n14167_ & new_n14169_;
  assign new_n14167_ = \all_features[2391]  & (\all_features[2390]  | (\all_features[2389]  & (\all_features[2388]  | ~new_n14168_ | ~new_n12357_)));
  assign new_n14168_ = ~\all_features[2386]  & ~\all_features[2387] ;
  assign new_n14169_ = \all_features[2391]  & (\all_features[2390]  | (new_n12362_ & (\all_features[2386]  | \all_features[2387]  | \all_features[2385] )));
  assign new_n14170_ = \all_features[2390]  & \all_features[2391]  & (\all_features[2388]  | \all_features[2389]  | new_n12361_ | ~new_n14168_);
  assign new_n14171_ = \all_features[2391]  & (\all_features[2389]  | \all_features[2390]  | \all_features[2388] );
  assign new_n14172_ = ~new_n14173_ & ~new_n14177_;
  assign new_n14173_ = ~new_n14174_ & ~new_n12367_;
  assign new_n14174_ = ~new_n12369_ & (new_n12363_ | (~new_n12359_ & (new_n12368_ | (~new_n12355_ & ~new_n14175_))));
  assign new_n14175_ = ~new_n12364_ & (new_n12370_ | (new_n14171_ & (~new_n14167_ | (~new_n14176_ & new_n14169_))));
  assign new_n14176_ = ~\all_features[2389]  & \all_features[2390]  & \all_features[2391]  & (\all_features[2388]  ? new_n14168_ : (new_n12361_ | ~new_n14168_));
  assign new_n14177_ = ~new_n12367_ & ~new_n12369_ & (~new_n12358_ | (~new_n12355_ & ~new_n14178_ & ~new_n12368_));
  assign new_n14178_ = ~new_n12364_ & ~new_n12370_ & (~new_n14171_ | ~new_n14167_ | new_n14179_);
  assign new_n14179_ = new_n14169_ & new_n14170_ & (new_n14180_ | ~\all_features[2389]  | ~\all_features[2390]  | ~\all_features[2391] );
  assign new_n14180_ = ~\all_features[2387]  & ~\all_features[2388]  & (~\all_features[2386]  | new_n12357_);
  assign new_n14181_ = ~new_n14182_ & new_n14206_;
  assign new_n14182_ = new_n14198_ & (~new_n14201_ | (~new_n14183_ & ~new_n14204_ & ~new_n14205_));
  assign new_n14183_ = ~new_n14192_ & ~new_n14194_ & (~new_n14197_ | ~new_n14196_ | new_n14184_);
  assign new_n14184_ = new_n14185_ & new_n14187_ & (new_n14190_ | ~\all_features[1509]  | ~\all_features[1510]  | ~\all_features[1511] );
  assign new_n14185_ = \all_features[1511]  & (\all_features[1510]  | (new_n14186_ & (\all_features[1506]  | \all_features[1507]  | \all_features[1505] )));
  assign new_n14186_ = \all_features[1508]  & \all_features[1509] ;
  assign new_n14187_ = \all_features[1510]  & \all_features[1511]  & (\all_features[1508]  | \all_features[1509]  | new_n14188_ | ~new_n14189_);
  assign new_n14188_ = \all_features[1504]  & \all_features[1505] ;
  assign new_n14189_ = ~\all_features[1506]  & ~\all_features[1507] ;
  assign new_n14190_ = ~\all_features[1507]  & ~\all_features[1508]  & (~\all_features[1506]  | new_n14191_);
  assign new_n14191_ = ~\all_features[1504]  & ~\all_features[1505] ;
  assign new_n14192_ = ~new_n14193_ & ~\all_features[1511] ;
  assign new_n14193_ = \all_features[1509]  & \all_features[1510]  & (\all_features[1508]  | (\all_features[1506]  & \all_features[1507]  & \all_features[1505] ));
  assign new_n14194_ = ~\all_features[1511]  & (~\all_features[1510]  | ~new_n14188_ | ~new_n14186_ | ~new_n14195_);
  assign new_n14195_ = \all_features[1506]  & \all_features[1507] ;
  assign new_n14196_ = \all_features[1511]  & (\all_features[1510]  | (\all_features[1509]  & (\all_features[1508]  | ~new_n14189_ | ~new_n14191_)));
  assign new_n14197_ = \all_features[1511]  & (\all_features[1509]  | \all_features[1510]  | \all_features[1508] );
  assign new_n14198_ = ~new_n14199_ & (\all_features[1507]  | \all_features[1508]  | \all_features[1509]  | \all_features[1510]  | \all_features[1511] );
  assign new_n14199_ = ~\all_features[1509]  & new_n14200_ & ((~\all_features[1506]  & new_n14191_) | ~\all_features[1508]  | ~\all_features[1507] );
  assign new_n14200_ = ~\all_features[1510]  & ~\all_features[1511] ;
  assign new_n14201_ = ~new_n14202_ & ~new_n14203_;
  assign new_n14202_ = new_n14200_ & (~\all_features[1509]  | (~\all_features[1508]  & (~\all_features[1507]  | (~\all_features[1506]  & ~\all_features[1505] ))));
  assign new_n14203_ = new_n14200_ & (~\all_features[1507]  | ~new_n14186_ | (~\all_features[1506]  & ~new_n14188_));
  assign new_n14204_ = ~\all_features[1511]  & (~\all_features[1510]  | (~\all_features[1508]  & ~\all_features[1509]  & ~new_n14195_));
  assign new_n14205_ = ~\all_features[1511]  & (~\all_features[1510]  | (~\all_features[1509]  & (new_n14191_ | ~new_n14195_ | ~\all_features[1508] )));
  assign new_n14206_ = ~new_n14207_ & ~new_n14210_;
  assign new_n14207_ = new_n14198_ & new_n14201_ & (new_n14208_ | new_n14205_ | new_n14192_ | ~new_n14209_);
  assign new_n14208_ = new_n14197_ & new_n14187_ & new_n14196_ & new_n14185_;
  assign new_n14209_ = ~new_n14204_ & ~new_n14194_;
  assign new_n14210_ = new_n14198_ & new_n14209_ & ~new_n14192_ & ~new_n14205_ & ~new_n14202_ & ~new_n14203_;
  assign new_n14211_ = ~new_n14212_ & ~new_n14235_;
  assign new_n14212_ = new_n14233_ & ~new_n14213_ & new_n14229_;
  assign new_n14213_ = ~new_n14228_ & ~new_n14227_ & ~new_n14225_ & ~new_n14214_ & ~new_n14217_;
  assign new_n14214_ = ~\all_features[4375]  & (~\all_features[4374]  | new_n14215_);
  assign new_n14215_ = ~\all_features[4373]  & (new_n14216_ | ~\all_features[4371]  | ~\all_features[4372]  | ~\all_features[4370] );
  assign new_n14216_ = ~\all_features[4368]  & ~\all_features[4369] ;
  assign new_n14217_ = new_n14224_ & new_n14222_ & new_n14218_ & new_n14220_;
  assign new_n14218_ = \all_features[4375]  & (\all_features[4374]  | (\all_features[4373]  & (\all_features[4372]  | ~new_n14219_ | ~new_n14216_)));
  assign new_n14219_ = ~\all_features[4370]  & ~\all_features[4371] ;
  assign new_n14220_ = \all_features[4375]  & (\all_features[4374]  | (new_n14221_ & (\all_features[4370]  | \all_features[4371]  | \all_features[4369] )));
  assign new_n14221_ = \all_features[4372]  & \all_features[4373] ;
  assign new_n14222_ = \all_features[4374]  & \all_features[4375]  & (\all_features[4372]  | \all_features[4373]  | new_n14223_ | ~new_n14219_);
  assign new_n14223_ = \all_features[4368]  & \all_features[4369] ;
  assign new_n14224_ = \all_features[4375]  & (\all_features[4373]  | \all_features[4374]  | \all_features[4372] );
  assign new_n14225_ = ~new_n14226_ & ~\all_features[4375] ;
  assign new_n14226_ = \all_features[4373]  & \all_features[4374]  & (\all_features[4372]  | (\all_features[4370]  & \all_features[4371]  & \all_features[4369] ));
  assign new_n14227_ = ~\all_features[4375]  & (~new_n14221_ | ~\all_features[4370]  | ~\all_features[4371]  | ~\all_features[4374]  | ~new_n14223_);
  assign new_n14228_ = ~\all_features[4375]  & (~\all_features[4374]  | (~\all_features[4373]  & ~\all_features[4372]  & (~\all_features[4371]  | ~\all_features[4370] )));
  assign new_n14229_ = ~new_n14230_ & ~new_n14232_;
  assign new_n14230_ = new_n14231_ & (~\all_features[4371]  | ~new_n14221_ | (~\all_features[4370]  & ~new_n14223_));
  assign new_n14231_ = ~\all_features[4374]  & ~\all_features[4375] ;
  assign new_n14232_ = new_n14231_ & (~\all_features[4373]  | (~\all_features[4372]  & (~\all_features[4371]  | (~\all_features[4370]  & ~\all_features[4369] ))));
  assign new_n14233_ = ~new_n14234_ & (\all_features[4371]  | \all_features[4372]  | \all_features[4373]  | \all_features[4374]  | \all_features[4375] );
  assign new_n14234_ = ~\all_features[4373]  & new_n14231_ & ((~\all_features[4370]  & new_n14216_) | ~\all_features[4372]  | ~\all_features[4371] );
  assign new_n14235_ = new_n14229_ & new_n14236_ & ~new_n14228_ & ~new_n14234_ & ~new_n14214_ & ~new_n14225_;
  assign new_n14236_ = ~new_n14227_ & (\all_features[4371]  | \all_features[4372]  | \all_features[4373]  | \all_features[4374]  | \all_features[4375] );
  assign new_n14237_ = new_n14233_ & (~new_n14229_ | (~new_n14238_ & ~new_n14214_ & ~new_n14228_));
  assign new_n14238_ = ~new_n14225_ & ~new_n14227_ & (~new_n14224_ | ~new_n14218_ | new_n14239_);
  assign new_n14239_ = new_n14220_ & new_n14222_ & (new_n14240_ | ~\all_features[4373]  | ~\all_features[4374]  | ~\all_features[4375] );
  assign new_n14240_ = ~\all_features[4371]  & ~\all_features[4372]  & (~\all_features[4370]  | new_n14216_);
  assign new_n14241_ = ~new_n14242_ & ~new_n14124_ & ~new_n14158_;
  assign new_n14242_ = new_n14273_ & new_n14269_ & new_n14243_ & new_n14264_;
  assign new_n14243_ = ~new_n14244_ & (\all_features[1531]  | \all_features[1532]  | \all_features[1533]  | \all_features[1534]  | \all_features[1535] );
  assign new_n14244_ = ~new_n14258_ & (new_n14260_ | (~new_n14261_ & (new_n14262_ | (~new_n14245_ & ~new_n14263_))));
  assign new_n14245_ = ~new_n14246_ & (new_n14248_ | (new_n14257_ & (~new_n14252_ | (~new_n14256_ & new_n14255_))));
  assign new_n14246_ = ~new_n14247_ & ~\all_features[1535] ;
  assign new_n14247_ = \all_features[1533]  & \all_features[1534]  & (\all_features[1532]  | (\all_features[1530]  & \all_features[1531]  & \all_features[1529] ));
  assign new_n14248_ = ~\all_features[1535]  & (~\all_features[1534]  | ~new_n14249_ | ~new_n14250_ | ~new_n14251_);
  assign new_n14249_ = \all_features[1528]  & \all_features[1529] ;
  assign new_n14250_ = \all_features[1532]  & \all_features[1533] ;
  assign new_n14251_ = \all_features[1530]  & \all_features[1531] ;
  assign new_n14252_ = \all_features[1535]  & (\all_features[1534]  | (\all_features[1533]  & (\all_features[1532]  | ~new_n14254_ | ~new_n14253_)));
  assign new_n14253_ = ~\all_features[1528]  & ~\all_features[1529] ;
  assign new_n14254_ = ~\all_features[1530]  & ~\all_features[1531] ;
  assign new_n14255_ = \all_features[1535]  & (\all_features[1534]  | (new_n14250_ & (\all_features[1530]  | \all_features[1531]  | \all_features[1529] )));
  assign new_n14256_ = ~\all_features[1533]  & \all_features[1534]  & \all_features[1535]  & (\all_features[1532]  ? new_n14254_ : (new_n14249_ | ~new_n14254_));
  assign new_n14257_ = \all_features[1535]  & (\all_features[1533]  | \all_features[1534]  | \all_features[1532] );
  assign new_n14258_ = ~\all_features[1533]  & new_n14259_ & ((~\all_features[1530]  & new_n14253_) | ~\all_features[1532]  | ~\all_features[1531] );
  assign new_n14259_ = ~\all_features[1534]  & ~\all_features[1535] ;
  assign new_n14260_ = new_n14259_ & (~\all_features[1533]  | (~\all_features[1532]  & (~\all_features[1531]  | (~\all_features[1530]  & ~\all_features[1529] ))));
  assign new_n14261_ = new_n14259_ & (~\all_features[1531]  | ~new_n14250_ | (~\all_features[1530]  & ~new_n14249_));
  assign new_n14262_ = ~\all_features[1535]  & (~\all_features[1534]  | (~\all_features[1532]  & ~\all_features[1533]  & ~new_n14251_));
  assign new_n14263_ = ~\all_features[1535]  & (~\all_features[1534]  | (~\all_features[1533]  & (new_n14253_ | ~new_n14251_ | ~\all_features[1532] )));
  assign new_n14264_ = new_n14268_ & ~new_n14261_ & ~new_n14265_ & ~new_n14260_;
  assign new_n14265_ = new_n14266_ & (~new_n14267_ | ~new_n14257_ | ~new_n14252_ | ~new_n14255_);
  assign new_n14266_ = ~new_n14248_ & ~new_n14246_ & ~new_n14262_ & ~new_n14263_;
  assign new_n14267_ = \all_features[1534]  & \all_features[1535]  & (\all_features[1532]  | \all_features[1533]  | new_n14249_ | ~new_n14254_);
  assign new_n14268_ = ~new_n14258_ & (\all_features[1531]  | \all_features[1532]  | \all_features[1533]  | \all_features[1534]  | \all_features[1535] );
  assign new_n14269_ = new_n14268_ & (new_n14261_ | new_n14260_ | (~new_n14270_ & ~new_n14262_ & ~new_n14263_));
  assign new_n14270_ = ~new_n14246_ & ~new_n14248_ & (~new_n14257_ | ~new_n14252_ | new_n14271_);
  assign new_n14271_ = new_n14255_ & new_n14267_ & (new_n14272_ | ~\all_features[1533]  | ~\all_features[1534]  | ~\all_features[1535] );
  assign new_n14272_ = ~\all_features[1531]  & ~\all_features[1532]  & (~\all_features[1530]  | new_n14253_);
  assign new_n14273_ = new_n14274_ & new_n14268_ & ~new_n14260_ & ~new_n14246_;
  assign new_n14274_ = ~new_n14248_ & ~new_n14263_ & ~new_n14261_ & ~new_n14262_;
  assign new_n14275_ = ~new_n14162_ & ~new_n14276_;
  assign new_n14276_ = new_n12717_ & new_n14277_;
  assign new_n14277_ = new_n12688_ & new_n12709_;
  assign new_n14278_ = new_n14279_ & ~new_n11199_ & ~new_n11201_;
  assign new_n14279_ = ~new_n11173_ & (new_n11195_ | (~new_n11194_ & (new_n11192_ | new_n14280_)));
  assign new_n14280_ = ~new_n11190_ & (new_n11186_ | (~new_n11188_ & (new_n11196_ | (~new_n14281_ & ~new_n11198_))));
  assign new_n14281_ = ~new_n14282_ & \all_features[3439]  & (\all_features[3438]  | \all_features[3437]  | \all_features[3436] );
  assign new_n14282_ = \all_features[3439]  & ((~new_n14283_ & ~\all_features[3437]  & \all_features[3438] ) | (~new_n11180_ & (\all_features[3438]  | (~new_n11176_ & \all_features[3437] ))));
  assign new_n14283_ = (\all_features[3436]  & ~new_n11178_) | (~new_n11183_ & ~\all_features[3436]  & new_n11178_);
  assign new_n14284_ = new_n14285_ ^ new_n14432_;
  assign new_n14285_ = new_n14286_ & (~new_n14430_ | (new_n14427_ & (new_n14429_ | new_n14428_)));
  assign new_n14286_ = ~new_n14287_ & new_n14347_ & (~new_n14389_ | (new_n14392_ & new_n14390_) | (new_n14426_ & ~new_n14390_));
  assign new_n14287_ = new_n14288_ & (new_n14293_ ? ~new_n14329_ : ~new_n14336_);
  assign new_n14288_ = new_n14289_ & new_n14290_;
  assign new_n14289_ = ~new_n6532_ | (~new_n6529_ & ~new_n6498_);
  assign new_n14290_ = new_n14291_ & new_n14292_;
  assign new_n14291_ = new_n11204_ & new_n11228_;
  assign new_n14292_ = new_n11233_ & new_n11236_;
  assign new_n14293_ = new_n14294_ & new_n14320_;
  assign new_n14294_ = ~new_n14295_ & ~new_n14317_;
  assign new_n14295_ = ~new_n14316_ & ~new_n14315_ & ~new_n14314_ & ~new_n14296_ & ~new_n14312_;
  assign new_n14296_ = new_n14297_ & (~new_n14310_ | ~new_n14311_ | ~new_n14307_ | ~new_n14309_);
  assign new_n14297_ = ~new_n14304_ & ~new_n14303_ & ~new_n14298_ & ~new_n14301_;
  assign new_n14298_ = ~\all_features[1671]  & (~\all_features[1670]  | (~\all_features[1669]  & (new_n14299_ | ~new_n14300_ | ~\all_features[1668] )));
  assign new_n14299_ = ~\all_features[1664]  & ~\all_features[1665] ;
  assign new_n14300_ = \all_features[1666]  & \all_features[1667] ;
  assign new_n14301_ = ~new_n14302_ & ~\all_features[1671] ;
  assign new_n14302_ = \all_features[1669]  & \all_features[1670]  & (\all_features[1668]  | (\all_features[1666]  & \all_features[1667]  & \all_features[1665] ));
  assign new_n14303_ = ~\all_features[1671]  & (~\all_features[1670]  | (~\all_features[1668]  & ~\all_features[1669]  & ~new_n14300_));
  assign new_n14304_ = ~\all_features[1671]  & (~\all_features[1670]  | ~new_n14305_ | ~new_n14306_ | ~new_n14300_);
  assign new_n14305_ = \all_features[1668]  & \all_features[1669] ;
  assign new_n14306_ = \all_features[1664]  & \all_features[1665] ;
  assign new_n14307_ = \all_features[1671]  & (\all_features[1670]  | (\all_features[1669]  & (\all_features[1668]  | ~new_n14299_ | ~new_n14308_)));
  assign new_n14308_ = ~\all_features[1666]  & ~\all_features[1667] ;
  assign new_n14309_ = \all_features[1671]  & (\all_features[1670]  | (new_n14305_ & (\all_features[1666]  | \all_features[1667]  | \all_features[1665] )));
  assign new_n14310_ = \all_features[1670]  & \all_features[1671]  & (\all_features[1668]  | \all_features[1669]  | new_n14306_ | ~new_n14308_);
  assign new_n14311_ = \all_features[1671]  & (\all_features[1669]  | \all_features[1670]  | \all_features[1668] );
  assign new_n14312_ = new_n14313_ & (~\all_features[1669]  | (~\all_features[1668]  & (~\all_features[1667]  | (~\all_features[1666]  & ~\all_features[1665] ))));
  assign new_n14313_ = ~\all_features[1670]  & ~\all_features[1671] ;
  assign new_n14314_ = ~\all_features[1669]  & new_n14313_ & ((~\all_features[1666]  & new_n14299_) | ~\all_features[1668]  | ~\all_features[1667] );
  assign new_n14315_ = new_n14313_ & (~\all_features[1667]  | ~new_n14305_ | (~\all_features[1666]  & ~new_n14306_));
  assign new_n14316_ = ~\all_features[1671]  & ~\all_features[1670]  & ~\all_features[1669]  & ~\all_features[1667]  & ~\all_features[1668] ;
  assign new_n14317_ = new_n14319_ & new_n14318_ & ~new_n14314_ & ~new_n14304_ & ~new_n14298_ & ~new_n14301_;
  assign new_n14318_ = ~new_n14303_ & ~new_n14316_;
  assign new_n14319_ = ~new_n14312_ & ~new_n14315_;
  assign new_n14320_ = ~new_n14321_ & ~new_n14325_;
  assign new_n14321_ = ~new_n14314_ & ~new_n14316_ & (~new_n14319_ | (~new_n14322_ & ~new_n14298_ & ~new_n14303_));
  assign new_n14322_ = ~new_n14304_ & ~new_n14301_ & (~new_n14311_ | ~new_n14307_ | new_n14323_);
  assign new_n14323_ = new_n14309_ & new_n14310_ & (new_n14324_ | ~\all_features[1669]  | ~\all_features[1670]  | ~\all_features[1671] );
  assign new_n14324_ = ~\all_features[1667]  & ~\all_features[1668]  & (~\all_features[1666]  | new_n14299_);
  assign new_n14325_ = ~new_n14326_ & ~new_n14316_;
  assign new_n14326_ = ~new_n14314_ & (new_n14312_ | (~new_n14315_ & (new_n14303_ | (~new_n14298_ & ~new_n14327_))));
  assign new_n14327_ = ~new_n14301_ & (new_n14304_ | (new_n14311_ & (~new_n14307_ | (~new_n14328_ & new_n14309_))));
  assign new_n14328_ = ~\all_features[1669]  & \all_features[1670]  & \all_features[1671]  & (\all_features[1668]  ? new_n14308_ : (new_n14306_ | ~new_n14308_));
  assign new_n14329_ = new_n14330_ & ~new_n10801_ & ~new_n14331_;
  assign new_n14330_ = ~new_n10778_ & ~new_n10834_;
  assign new_n14331_ = ~new_n10794_ & (new_n10797_ | (~new_n10800_ & (new_n10799_ | (~new_n14332_ & ~new_n10791_))));
  assign new_n14332_ = ~new_n10787_ & (new_n10789_ | (~new_n10792_ & (~new_n14335_ | new_n14333_)));
  assign new_n14333_ = \all_features[4391]  & ((~new_n14334_ & ~\all_features[4389]  & \all_features[4390] ) | (~new_n10784_ & (\all_features[4390]  | (~new_n10781_ & \all_features[4389] ))));
  assign new_n14334_ = (~\all_features[4386]  & ~\all_features[4387]  & ~\all_features[4388]  & (~\all_features[4385]  | ~\all_features[4384] )) | (\all_features[4388]  & (\all_features[4386]  | \all_features[4387] ));
  assign new_n14335_ = \all_features[4391]  & (\all_features[4389]  | \all_features[4390]  | \all_features[4388] );
  assign new_n14336_ = new_n14337_ & new_n14338_;
  assign new_n14337_ = ~new_n13015_ & ~new_n13038_;
  assign new_n14338_ = ~new_n14339_ & ~new_n14343_;
  assign new_n14339_ = new_n13033_ & (~new_n13039_ | (~new_n14340_ & ~new_n13027_ & ~new_n13031_));
  assign new_n14340_ = ~new_n13032_ & ~new_n13025_ & (~new_n13023_ | ~new_n13029_ | new_n14341_);
  assign new_n14341_ = new_n13018_ & new_n13020_ & (new_n14342_ | ~\all_features[2605]  | ~\all_features[2606]  | ~\all_features[2607] );
  assign new_n14342_ = ~\all_features[2603]  & ~\all_features[2604]  & (~\all_features[2602]  | new_n13030_);
  assign new_n14343_ = ~new_n14344_ & (\all_features[2603]  | \all_features[2604]  | \all_features[2605]  | \all_features[2606]  | \all_features[2607] );
  assign new_n14344_ = ~new_n13034_ & (new_n13036_ | (~new_n13037_ & (new_n13027_ | (~new_n13031_ & ~new_n14345_))));
  assign new_n14345_ = ~new_n13025_ & (new_n13032_ | (new_n13023_ & (~new_n13029_ | (~new_n14346_ & new_n13018_))));
  assign new_n14346_ = ~\all_features[2605]  & \all_features[2606]  & \all_features[2607]  & (\all_features[2604]  ? new_n13021_ : (new_n13022_ | ~new_n13021_));
  assign new_n14347_ = (new_n14387_ | ~new_n14386_) & (new_n14388_ | ~new_n14348_);
  assign new_n14348_ = new_n14384_ & ~new_n14289_ & ~new_n14349_;
  assign new_n14349_ = ~new_n14380_ & new_n14350_;
  assign new_n14350_ = ~new_n14376_ & new_n14351_;
  assign new_n14351_ = ~new_n14352_ & ~new_n14374_;
  assign new_n14352_ = new_n14369_ & ~new_n14373_ & ~new_n14353_ & ~new_n14372_;
  assign new_n14353_ = new_n14354_ & (~new_n14367_ | ~new_n14368_ | ~new_n14364_ | ~new_n14366_);
  assign new_n14354_ = ~new_n14361_ & ~new_n14359_ & ~new_n14355_ & ~new_n14357_;
  assign new_n14355_ = ~\all_features[4407]  & (~\all_features[4406]  | (~\all_features[4404]  & ~\all_features[4405]  & ~new_n14356_));
  assign new_n14356_ = \all_features[4402]  & \all_features[4403] ;
  assign new_n14357_ = ~\all_features[4407]  & (~\all_features[4406]  | (~\all_features[4405]  & (new_n14358_ | ~new_n14356_ | ~\all_features[4404] )));
  assign new_n14358_ = ~\all_features[4400]  & ~\all_features[4401] ;
  assign new_n14359_ = ~new_n14360_ & ~\all_features[4407] ;
  assign new_n14360_ = \all_features[4405]  & \all_features[4406]  & (\all_features[4404]  | (\all_features[4402]  & \all_features[4403]  & \all_features[4401] ));
  assign new_n14361_ = ~\all_features[4407]  & (~\all_features[4406]  | ~new_n14362_ | ~new_n14363_ | ~new_n14356_);
  assign new_n14362_ = \all_features[4400]  & \all_features[4401] ;
  assign new_n14363_ = \all_features[4404]  & \all_features[4405] ;
  assign new_n14364_ = \all_features[4407]  & (\all_features[4406]  | (\all_features[4405]  & (\all_features[4404]  | ~new_n14365_ | ~new_n14358_)));
  assign new_n14365_ = ~\all_features[4402]  & ~\all_features[4403] ;
  assign new_n14366_ = \all_features[4407]  & (\all_features[4406]  | (new_n14363_ & (\all_features[4402]  | \all_features[4403]  | \all_features[4401] )));
  assign new_n14367_ = \all_features[4406]  & \all_features[4407]  & (\all_features[4404]  | \all_features[4405]  | new_n14362_ | ~new_n14365_);
  assign new_n14368_ = \all_features[4407]  & (\all_features[4405]  | \all_features[4406]  | \all_features[4404] );
  assign new_n14369_ = ~new_n14370_ & (\all_features[4403]  | \all_features[4404]  | \all_features[4405]  | \all_features[4406]  | \all_features[4407] );
  assign new_n14370_ = ~\all_features[4405]  & new_n14371_ & ((~\all_features[4402]  & new_n14358_) | ~\all_features[4404]  | ~\all_features[4403] );
  assign new_n14371_ = ~\all_features[4406]  & ~\all_features[4407] ;
  assign new_n14372_ = new_n14371_ & (~\all_features[4405]  | (~\all_features[4404]  & (~\all_features[4403]  | (~\all_features[4402]  & ~\all_features[4401] ))));
  assign new_n14373_ = new_n14371_ & (~\all_features[4403]  | ~new_n14363_ | (~\all_features[4402]  & ~new_n14362_));
  assign new_n14374_ = new_n14375_ & new_n14369_ & ~new_n14372_ & ~new_n14359_;
  assign new_n14375_ = ~new_n14361_ & ~new_n14357_ & ~new_n14373_ & ~new_n14355_;
  assign new_n14376_ = new_n14369_ & (new_n14373_ | new_n14372_ | (~new_n14377_ & ~new_n14355_ & ~new_n14357_));
  assign new_n14377_ = ~new_n14359_ & ~new_n14361_ & (~new_n14368_ | ~new_n14364_ | new_n14378_);
  assign new_n14378_ = new_n14366_ & new_n14367_ & (new_n14379_ | ~\all_features[4405]  | ~\all_features[4406]  | ~\all_features[4407] );
  assign new_n14379_ = ~\all_features[4403]  & ~\all_features[4404]  & (~\all_features[4402]  | new_n14358_);
  assign new_n14380_ = ~new_n14381_ & (\all_features[4403]  | \all_features[4404]  | \all_features[4405]  | \all_features[4406]  | \all_features[4407] );
  assign new_n14381_ = ~new_n14370_ & (new_n14372_ | (~new_n14373_ & (new_n14355_ | (~new_n14382_ & ~new_n14357_))));
  assign new_n14382_ = ~new_n14359_ & (new_n14361_ | (new_n14368_ & (~new_n14364_ | (~new_n14383_ & new_n14366_))));
  assign new_n14383_ = ~\all_features[4405]  & \all_features[4406]  & \all_features[4407]  & (\all_features[4404]  ? new_n14365_ : (new_n14362_ | ~new_n14365_));
  assign new_n14384_ = new_n12534_ & new_n14385_;
  assign new_n14385_ = ~new_n9271_ & ~new_n12530_;
  assign new_n14386_ = ~new_n14290_ & new_n14289_;
  assign new_n14387_ = new_n14292_ & ~new_n11203_ & new_n13887_;
  assign new_n14388_ = new_n8693_ & new_n8697_ & new_n8669_;
  assign new_n14389_ = ~new_n14289_ & ~new_n14384_;
  assign new_n14390_ = new_n7581_ & new_n14391_ & new_n7559_;
  assign new_n14391_ = new_n7587_ & new_n7583_;
  assign new_n14392_ = new_n14393_ & new_n14417_;
  assign new_n14393_ = ~new_n14394_ & ~new_n14416_;
  assign new_n14394_ = new_n14395_ & (~new_n14404_ | (new_n14414_ & new_n14415_ & new_n14411_ & new_n14413_));
  assign new_n14395_ = new_n14396_ & ~new_n14400_ & ~new_n14401_;
  assign new_n14396_ = ~new_n14397_ & (\all_features[2995]  | \all_features[2996]  | \all_features[2997]  | \all_features[2998]  | \all_features[2999] );
  assign new_n14397_ = ~\all_features[2997]  & new_n14399_ & ((~\all_features[2994]  & new_n14398_) | ~\all_features[2996]  | ~\all_features[2995] );
  assign new_n14398_ = ~\all_features[2992]  & ~\all_features[2993] ;
  assign new_n14399_ = ~\all_features[2998]  & ~\all_features[2999] ;
  assign new_n14400_ = new_n14399_ & (~\all_features[2997]  | (~\all_features[2996]  & (~\all_features[2995]  | (~\all_features[2994]  & ~\all_features[2993] ))));
  assign new_n14401_ = new_n14399_ & (~\all_features[2995]  | ~new_n14402_ | (~\all_features[2994]  & ~new_n14403_));
  assign new_n14402_ = \all_features[2996]  & \all_features[2997] ;
  assign new_n14403_ = \all_features[2992]  & \all_features[2993] ;
  assign new_n14404_ = ~new_n14410_ & ~new_n14409_ & ~new_n14405_ & ~new_n14407_;
  assign new_n14405_ = ~\all_features[2999]  & (~\all_features[2998]  | (~\all_features[2997]  & (new_n14398_ | ~new_n14406_ | ~\all_features[2996] )));
  assign new_n14406_ = \all_features[2994]  & \all_features[2995] ;
  assign new_n14407_ = ~new_n14408_ & ~\all_features[2999] ;
  assign new_n14408_ = \all_features[2997]  & \all_features[2998]  & (\all_features[2996]  | (\all_features[2994]  & \all_features[2995]  & \all_features[2993] ));
  assign new_n14409_ = ~\all_features[2999]  & (~\all_features[2998]  | ~new_n14402_ | ~new_n14403_ | ~new_n14406_);
  assign new_n14410_ = ~\all_features[2999]  & (~\all_features[2998]  | (~\all_features[2996]  & ~\all_features[2997]  & ~new_n14406_));
  assign new_n14411_ = \all_features[2999]  & (\all_features[2998]  | (\all_features[2997]  & (\all_features[2996]  | ~new_n14398_ | ~new_n14412_)));
  assign new_n14412_ = ~\all_features[2994]  & ~\all_features[2995] ;
  assign new_n14413_ = \all_features[2999]  & (\all_features[2998]  | (new_n14402_ & (\all_features[2994]  | \all_features[2995]  | \all_features[2993] )));
  assign new_n14414_ = \all_features[2998]  & \all_features[2999]  & (\all_features[2996]  | \all_features[2997]  | new_n14403_ | ~new_n14412_);
  assign new_n14415_ = \all_features[2999]  & (\all_features[2997]  | \all_features[2998]  | \all_features[2996] );
  assign new_n14416_ = new_n14395_ & new_n14404_;
  assign new_n14417_ = ~new_n14418_ & ~new_n14422_;
  assign new_n14418_ = ~new_n14419_ & (\all_features[2995]  | \all_features[2996]  | \all_features[2997]  | \all_features[2998]  | \all_features[2999] );
  assign new_n14419_ = ~new_n14397_ & (new_n14400_ | (~new_n14401_ & (new_n14410_ | (~new_n14405_ & ~new_n14420_))));
  assign new_n14420_ = ~new_n14407_ & (new_n14409_ | (new_n14415_ & (~new_n14411_ | (~new_n14421_ & new_n14413_))));
  assign new_n14421_ = ~\all_features[2997]  & \all_features[2998]  & \all_features[2999]  & (\all_features[2996]  ? new_n14412_ : (new_n14403_ | ~new_n14412_));
  assign new_n14422_ = new_n14396_ & (new_n14401_ | new_n14400_ | (~new_n14405_ & ~new_n14410_ & ~new_n14423_));
  assign new_n14423_ = ~new_n14409_ & ~new_n14407_ & (~new_n14415_ | ~new_n14411_ | new_n14424_);
  assign new_n14424_ = new_n14413_ & new_n14414_ & (new_n14425_ | ~\all_features[2997]  | ~\all_features[2998]  | ~\all_features[2999] );
  assign new_n14425_ = ~\all_features[2995]  & ~\all_features[2996]  & (~\all_features[2994]  | new_n14398_);
  assign new_n14426_ = new_n9644_ & new_n9649_;
  assign new_n14427_ = (~new_n14348_ | ~new_n14388_) & (~new_n14387_ | ~new_n14386_);
  assign new_n14428_ = new_n14329_ & new_n14288_ & new_n14293_;
  assign new_n14429_ = new_n14392_ & new_n14389_ & new_n14390_;
  assign new_n14430_ = (new_n14431_ | new_n14289_) & (new_n14293_ | ~new_n14290_ | ~new_n14336_ | ~new_n14289_);
  assign new_n14431_ = (new_n11095_ | ~new_n14349_ | ~new_n14384_) & (new_n14390_ | ~new_n14426_ | new_n14384_);
  assign new_n14432_ = ~new_n14433_ & new_n14611_;
  assign new_n14433_ = ~new_n14434_ & new_n14575_ & new_n14550_ & (new_n14384_ | ~new_n14549_);
  assign new_n14434_ = ~new_n14435_ & ((~new_n14469_ & new_n14539_ & new_n14503_) | (new_n14289_ & ~new_n14503_));
  assign new_n14435_ = ~new_n14465_ & new_n14436_;
  assign new_n14436_ = ~new_n14463_ & ~new_n14437_ & ~new_n14461_;
  assign new_n14437_ = new_n14453_ & (~new_n14456_ | (~new_n14438_ & ~new_n14459_ & ~new_n14460_));
  assign new_n14438_ = ~new_n14447_ & ~new_n14449_ & (~new_n14452_ | ~new_n14451_ | new_n14439_);
  assign new_n14439_ = new_n14440_ & new_n14442_ & (new_n14445_ | ~\all_features[3061]  | ~\all_features[3062]  | ~\all_features[3063] );
  assign new_n14440_ = \all_features[3063]  & (\all_features[3062]  | (new_n14441_ & (\all_features[3058]  | \all_features[3059]  | \all_features[3057] )));
  assign new_n14441_ = \all_features[3060]  & \all_features[3061] ;
  assign new_n14442_ = \all_features[3062]  & \all_features[3063]  & (\all_features[3060]  | \all_features[3061]  | new_n14443_ | ~new_n14444_);
  assign new_n14443_ = \all_features[3056]  & \all_features[3057] ;
  assign new_n14444_ = ~\all_features[3058]  & ~\all_features[3059] ;
  assign new_n14445_ = ~\all_features[3059]  & ~\all_features[3060]  & (~\all_features[3058]  | new_n14446_);
  assign new_n14446_ = ~\all_features[3056]  & ~\all_features[3057] ;
  assign new_n14447_ = ~new_n14448_ & ~\all_features[3063] ;
  assign new_n14448_ = \all_features[3061]  & \all_features[3062]  & (\all_features[3060]  | (\all_features[3058]  & \all_features[3059]  & \all_features[3057] ));
  assign new_n14449_ = ~\all_features[3063]  & (~\all_features[3062]  | ~new_n14450_ | ~new_n14443_ | ~new_n14441_);
  assign new_n14450_ = \all_features[3058]  & \all_features[3059] ;
  assign new_n14451_ = \all_features[3063]  & (\all_features[3062]  | (\all_features[3061]  & (\all_features[3060]  | ~new_n14444_ | ~new_n14446_)));
  assign new_n14452_ = \all_features[3063]  & (\all_features[3061]  | \all_features[3062]  | \all_features[3060] );
  assign new_n14453_ = ~new_n14454_ & (\all_features[3059]  | \all_features[3060]  | \all_features[3061]  | \all_features[3062]  | \all_features[3063] );
  assign new_n14454_ = ~\all_features[3061]  & new_n14455_ & ((~\all_features[3058]  & new_n14446_) | ~\all_features[3060]  | ~\all_features[3059] );
  assign new_n14455_ = ~\all_features[3062]  & ~\all_features[3063] ;
  assign new_n14456_ = ~new_n14457_ & ~new_n14458_;
  assign new_n14457_ = new_n14455_ & (~\all_features[3061]  | (~\all_features[3060]  & (~\all_features[3059]  | (~\all_features[3058]  & ~\all_features[3057] ))));
  assign new_n14458_ = new_n14455_ & (~\all_features[3059]  | ~new_n14441_ | (~\all_features[3058]  & ~new_n14443_));
  assign new_n14459_ = ~\all_features[3063]  & (~\all_features[3062]  | (~\all_features[3061]  & (new_n14446_ | ~new_n14450_ | ~\all_features[3060] )));
  assign new_n14460_ = ~\all_features[3063]  & (~\all_features[3062]  | (~\all_features[3060]  & ~\all_features[3061]  & ~new_n14450_));
  assign new_n14461_ = new_n14462_ & new_n14453_ & ~new_n14458_ & ~new_n14459_ & ~new_n14447_ & ~new_n14457_;
  assign new_n14462_ = ~new_n14449_ & ~new_n14460_;
  assign new_n14463_ = new_n14453_ & new_n14456_ & (new_n14464_ | new_n14447_ | new_n14459_ | ~new_n14462_);
  assign new_n14464_ = new_n14452_ & new_n14442_ & new_n14451_ & new_n14440_;
  assign new_n14465_ = ~new_n14466_ & (\all_features[3059]  | \all_features[3060]  | \all_features[3061]  | \all_features[3062]  | \all_features[3063] );
  assign new_n14466_ = ~new_n14454_ & (new_n14457_ | (~new_n14458_ & (new_n14460_ | (~new_n14459_ & ~new_n14467_))));
  assign new_n14467_ = ~new_n14447_ & (new_n14449_ | (new_n14452_ & (~new_n14451_ | (~new_n14468_ & new_n14440_))));
  assign new_n14468_ = ~\all_features[3061]  & \all_features[3062]  & \all_features[3063]  & (\all_features[3060]  ? new_n14444_ : (new_n14443_ | ~new_n14444_));
  assign new_n14469_ = new_n14470_ & new_n14494_;
  assign new_n14470_ = ~new_n14471_ & ~new_n14493_;
  assign new_n14471_ = new_n14472_ & (~new_n14481_ | (new_n14491_ & new_n14492_ & new_n14488_ & new_n14490_));
  assign new_n14472_ = new_n14473_ & ~new_n14477_ & ~new_n14478_;
  assign new_n14473_ = ~new_n14474_ & (\all_features[2099]  | \all_features[2100]  | \all_features[2101]  | \all_features[2102]  | \all_features[2103] );
  assign new_n14474_ = ~\all_features[2101]  & new_n14476_ & ((~\all_features[2098]  & new_n14475_) | ~\all_features[2100]  | ~\all_features[2099] );
  assign new_n14475_ = ~\all_features[2096]  & ~\all_features[2097] ;
  assign new_n14476_ = ~\all_features[2102]  & ~\all_features[2103] ;
  assign new_n14477_ = new_n14476_ & (~\all_features[2101]  | (~\all_features[2100]  & (~\all_features[2099]  | (~\all_features[2098]  & ~\all_features[2097] ))));
  assign new_n14478_ = new_n14476_ & (~\all_features[2099]  | ~new_n14479_ | (~\all_features[2098]  & ~new_n14480_));
  assign new_n14479_ = \all_features[2100]  & \all_features[2101] ;
  assign new_n14480_ = \all_features[2096]  & \all_features[2097] ;
  assign new_n14481_ = ~new_n14487_ & ~new_n14486_ & ~new_n14482_ & ~new_n14484_;
  assign new_n14482_ = ~\all_features[2103]  & (~\all_features[2102]  | (~\all_features[2101]  & (new_n14475_ | ~new_n14483_ | ~\all_features[2100] )));
  assign new_n14483_ = \all_features[2098]  & \all_features[2099] ;
  assign new_n14484_ = ~new_n14485_ & ~\all_features[2103] ;
  assign new_n14485_ = \all_features[2101]  & \all_features[2102]  & (\all_features[2100]  | (\all_features[2098]  & \all_features[2099]  & \all_features[2097] ));
  assign new_n14486_ = ~\all_features[2103]  & (~\all_features[2102]  | ~new_n14479_ | ~new_n14480_ | ~new_n14483_);
  assign new_n14487_ = ~\all_features[2103]  & (~\all_features[2102]  | (~\all_features[2100]  & ~\all_features[2101]  & ~new_n14483_));
  assign new_n14488_ = \all_features[2103]  & (\all_features[2102]  | (\all_features[2101]  & (\all_features[2100]  | ~new_n14475_ | ~new_n14489_)));
  assign new_n14489_ = ~\all_features[2098]  & ~\all_features[2099] ;
  assign new_n14490_ = \all_features[2103]  & (\all_features[2102]  | (new_n14479_ & (\all_features[2098]  | \all_features[2099]  | \all_features[2097] )));
  assign new_n14491_ = \all_features[2102]  & \all_features[2103]  & (\all_features[2100]  | \all_features[2101]  | new_n14480_ | ~new_n14489_);
  assign new_n14492_ = \all_features[2103]  & (\all_features[2101]  | \all_features[2102]  | \all_features[2100] );
  assign new_n14493_ = new_n14472_ & new_n14481_;
  assign new_n14494_ = ~new_n14495_ & ~new_n14499_;
  assign new_n14495_ = new_n14473_ & (new_n14478_ | new_n14477_ | (~new_n14482_ & ~new_n14487_ & ~new_n14496_));
  assign new_n14496_ = ~new_n14486_ & ~new_n14484_ & (~new_n14492_ | ~new_n14488_ | new_n14497_);
  assign new_n14497_ = new_n14490_ & new_n14491_ & (new_n14498_ | ~\all_features[2101]  | ~\all_features[2102]  | ~\all_features[2103] );
  assign new_n14498_ = ~\all_features[2099]  & ~\all_features[2100]  & (~\all_features[2098]  | new_n14475_);
  assign new_n14499_ = ~new_n14500_ & (\all_features[2099]  | \all_features[2100]  | \all_features[2101]  | \all_features[2102]  | \all_features[2103] );
  assign new_n14500_ = ~new_n14474_ & (new_n14477_ | (~new_n14478_ & (new_n14487_ | (~new_n14482_ & ~new_n14501_))));
  assign new_n14501_ = ~new_n14484_ & (new_n14486_ | (new_n14492_ & (~new_n14488_ | (~new_n14502_ & new_n14490_))));
  assign new_n14502_ = ~\all_features[2101]  & \all_features[2102]  & \all_features[2103]  & (\all_features[2100]  ? new_n14489_ : (new_n14480_ | ~new_n14489_));
  assign new_n14503_ = new_n14504_ & new_n14530_;
  assign new_n14504_ = new_n14505_ & new_n14528_;
  assign new_n14505_ = new_n14523_ & ~new_n14527_ & ~new_n14506_ & ~new_n14526_;
  assign new_n14506_ = ~new_n14521_ & ~new_n14522_ & new_n14514_ & (~new_n14519_ | ~new_n14507_);
  assign new_n14507_ = new_n14513_ & new_n14508_ & new_n14510_;
  assign new_n14508_ = \all_features[4135]  & (\all_features[4134]  | (new_n14509_ & (\all_features[4130]  | \all_features[4131]  | \all_features[4129] )));
  assign new_n14509_ = \all_features[4132]  & \all_features[4133] ;
  assign new_n14510_ = \all_features[4134]  & \all_features[4135]  & (\all_features[4132]  | \all_features[4133]  | new_n14512_ | ~new_n14511_);
  assign new_n14511_ = ~\all_features[4130]  & ~\all_features[4131] ;
  assign new_n14512_ = \all_features[4128]  & \all_features[4129] ;
  assign new_n14513_ = \all_features[4135]  & (\all_features[4133]  | \all_features[4134]  | \all_features[4132] );
  assign new_n14514_ = ~new_n14515_ & ~new_n14517_;
  assign new_n14515_ = ~new_n14516_ & ~\all_features[4135] ;
  assign new_n14516_ = \all_features[4133]  & \all_features[4134]  & (\all_features[4132]  | (\all_features[4130]  & \all_features[4131]  & \all_features[4129] ));
  assign new_n14517_ = ~\all_features[4135]  & (~\all_features[4134]  | (~\all_features[4132]  & ~\all_features[4133]  & ~new_n14518_));
  assign new_n14518_ = \all_features[4130]  & \all_features[4131] ;
  assign new_n14519_ = \all_features[4135]  & (\all_features[4134]  | (\all_features[4133]  & (\all_features[4132]  | ~new_n14520_ | ~new_n14511_)));
  assign new_n14520_ = ~\all_features[4128]  & ~\all_features[4129] ;
  assign new_n14521_ = ~\all_features[4135]  & (~\all_features[4134]  | (~\all_features[4133]  & (new_n14520_ | ~new_n14518_ | ~\all_features[4132] )));
  assign new_n14522_ = ~\all_features[4135]  & (~\all_features[4134]  | ~new_n14509_ | ~new_n14512_ | ~new_n14518_);
  assign new_n14523_ = ~new_n14524_ & (\all_features[4131]  | \all_features[4132]  | \all_features[4133]  | \all_features[4134]  | \all_features[4135] );
  assign new_n14524_ = ~\all_features[4133]  & new_n14525_ & ((~\all_features[4130]  & new_n14520_) | ~\all_features[4132]  | ~\all_features[4131] );
  assign new_n14525_ = ~\all_features[4134]  & ~\all_features[4135] ;
  assign new_n14526_ = new_n14525_ & (~\all_features[4133]  | (~\all_features[4132]  & (~\all_features[4131]  | (~\all_features[4130]  & ~\all_features[4129] ))));
  assign new_n14527_ = new_n14525_ & (~\all_features[4131]  | ~new_n14509_ | (~\all_features[4130]  & ~new_n14512_));
  assign new_n14528_ = new_n14523_ & new_n14514_ & new_n14529_ & ~new_n14521_ & ~new_n14522_;
  assign new_n14529_ = ~new_n14526_ & ~new_n14527_;
  assign new_n14530_ = new_n14531_ & new_n14535_;
  assign new_n14531_ = new_n14523_ & (~new_n14529_ | (~new_n14532_ & ~new_n14517_ & ~new_n14521_));
  assign new_n14532_ = ~new_n14522_ & ~new_n14515_ & (~new_n14513_ | ~new_n14519_ | new_n14533_);
  assign new_n14533_ = new_n14508_ & new_n14510_ & (new_n14534_ | ~\all_features[4133]  | ~\all_features[4134]  | ~\all_features[4135] );
  assign new_n14534_ = ~\all_features[4131]  & ~\all_features[4132]  & (~\all_features[4130]  | new_n14520_);
  assign new_n14535_ = ~new_n14536_ & (\all_features[4131]  | \all_features[4132]  | \all_features[4133]  | \all_features[4134]  | \all_features[4135] );
  assign new_n14536_ = ~new_n14524_ & (new_n14526_ | (~new_n14527_ & (new_n14517_ | (~new_n14521_ & ~new_n14537_))));
  assign new_n14537_ = ~new_n14515_ & (new_n14522_ | (new_n14513_ & (~new_n14519_ | (~new_n14538_ & new_n14508_))));
  assign new_n14538_ = ~\all_features[4133]  & \all_features[4134]  & \all_features[4135]  & (\all_features[4132]  ? new_n14511_ : (new_n14512_ | ~new_n14511_));
  assign new_n14539_ = ~new_n14540_ & new_n6674_;
  assign new_n14540_ = ~new_n14541_ & ~new_n14545_;
  assign new_n14541_ = ~new_n14542_ & (\all_features[2595]  | \all_features[2596]  | \all_features[2597]  | \all_features[2598]  | \all_features[2599] );
  assign new_n14542_ = ~new_n6694_ & (new_n6696_ | (~new_n6697_ & (new_n6687_ | (~new_n6691_ & ~new_n14543_))));
  assign new_n14543_ = ~new_n6685_ & (new_n6692_ | (new_n6683_ & (~new_n6689_ | (~new_n14544_ & new_n6678_))));
  assign new_n14544_ = ~\all_features[2597]  & \all_features[2598]  & \all_features[2599]  & (\all_features[2596]  ? new_n6681_ : (new_n6682_ | ~new_n6681_));
  assign new_n14545_ = new_n6693_ & (~new_n6699_ | (~new_n14546_ & ~new_n6687_ & ~new_n6691_));
  assign new_n14546_ = ~new_n6692_ & ~new_n6685_ & (~new_n6683_ | ~new_n6689_ | new_n14547_);
  assign new_n14547_ = new_n6678_ & new_n6680_ & (new_n14548_ | ~\all_features[2597]  | ~\all_features[2598]  | ~\all_features[2599] );
  assign new_n14548_ = ~\all_features[2595]  & ~\all_features[2596]  & (~\all_features[2594]  | new_n6690_);
  assign new_n14549_ = ~new_n14503_ & ~new_n14289_ & ~new_n14435_;
  assign new_n14550_ = (new_n9209_ | ~new_n11337_ | ~new_n11902_ | ~new_n14435_) & (new_n14293_ | ~new_n14551_);
  assign new_n14551_ = ~new_n11902_ & new_n14435_ & (~new_n14568_ | ~new_n14552_);
  assign new_n14552_ = new_n14553_ & new_n14562_;
  assign new_n14553_ = ~new_n14561_ & ~new_n14559_ & ~new_n14554_ & ~new_n14557_;
  assign new_n14554_ = ~\all_features[559]  & (~\all_features[558]  | (~\all_features[557]  & (new_n14556_ | ~\all_features[556]  | ~new_n14555_)));
  assign new_n14555_ = \all_features[554]  & \all_features[555] ;
  assign new_n14556_ = ~\all_features[552]  & ~\all_features[553] ;
  assign new_n14557_ = ~new_n14558_ & ~\all_features[559] ;
  assign new_n14558_ = \all_features[557]  & \all_features[558]  & (\all_features[556]  | (\all_features[554]  & \all_features[555]  & \all_features[553] ));
  assign new_n14559_ = ~\all_features[559]  & (~new_n14560_ | ~\all_features[552]  | ~\all_features[553]  | ~\all_features[558]  | ~new_n14555_);
  assign new_n14560_ = \all_features[556]  & \all_features[557] ;
  assign new_n14561_ = ~\all_features[559]  & (~\all_features[558]  | (~\all_features[556]  & ~\all_features[557]  & ~new_n14555_));
  assign new_n14562_ = ~new_n14567_ & ~new_n14566_ & ~new_n14563_ & ~new_n14565_;
  assign new_n14563_ = new_n14564_ & (~\all_features[557]  | (~\all_features[556]  & (~\all_features[555]  | (~\all_features[554]  & ~\all_features[553] ))));
  assign new_n14564_ = ~\all_features[558]  & ~\all_features[559] ;
  assign new_n14565_ = new_n14564_ & (~new_n14560_ | ~\all_features[555]  | (~\all_features[554]  & (~\all_features[552]  | ~\all_features[553] )));
  assign new_n14566_ = ~\all_features[557]  & new_n14564_ & ((~\all_features[554]  & new_n14556_) | ~\all_features[556]  | ~\all_features[555] );
  assign new_n14567_ = ~\all_features[559]  & ~\all_features[558]  & ~\all_features[557]  & ~\all_features[555]  & ~\all_features[556] ;
  assign new_n14568_ = new_n14562_ & (~new_n14553_ | (new_n14572_ & new_n14574_ & new_n14569_ & new_n14571_));
  assign new_n14569_ = \all_features[559]  & (\all_features[558]  | (\all_features[557]  & (\all_features[556]  | ~new_n14570_ | ~new_n14556_)));
  assign new_n14570_ = ~\all_features[554]  & ~\all_features[555] ;
  assign new_n14571_ = \all_features[559]  & (\all_features[558]  | (new_n14560_ & (\all_features[554]  | \all_features[555]  | \all_features[553] )));
  assign new_n14572_ = new_n14573_ & (\all_features[556]  | \all_features[557]  | ~new_n14570_ | (\all_features[553]  & \all_features[552] ));
  assign new_n14573_ = \all_features[558]  & \all_features[559] ;
  assign new_n14574_ = \all_features[559]  & (\all_features[557]  | \all_features[558]  | \all_features[556] );
  assign new_n14575_ = (new_n14158_ | ~new_n14577_) & (new_n14578_ | ~new_n14576_);
  assign new_n14576_ = new_n14435_ & ~new_n11337_ & new_n11902_;
  assign new_n14577_ = new_n14503_ & ~new_n14435_ & ~new_n14539_;
  assign new_n14578_ = ~new_n14607_ & (~new_n14609_ | (~new_n14600_ & ~new_n14579_));
  assign new_n14579_ = ~new_n14580_ & (\all_features[1291]  | \all_features[1292]  | \all_features[1293]  | \all_features[1294]  | \all_features[1295] );
  assign new_n14580_ = ~new_n14596_ & (new_n14594_ | (~new_n14598_ & (new_n14599_ | (~new_n14597_ & ~new_n14581_))));
  assign new_n14581_ = ~new_n14582_ & (new_n14584_ | (new_n14593_ & (~new_n14588_ | (~new_n14592_ & new_n14591_))));
  assign new_n14582_ = ~new_n14583_ & ~\all_features[1295] ;
  assign new_n14583_ = \all_features[1293]  & \all_features[1294]  & (\all_features[1292]  | (\all_features[1290]  & \all_features[1291]  & \all_features[1289] ));
  assign new_n14584_ = ~\all_features[1295]  & (~\all_features[1294]  | ~new_n14585_ | ~new_n14586_ | ~new_n14587_);
  assign new_n14585_ = \all_features[1290]  & \all_features[1291] ;
  assign new_n14586_ = \all_features[1288]  & \all_features[1289] ;
  assign new_n14587_ = \all_features[1292]  & \all_features[1293] ;
  assign new_n14588_ = \all_features[1295]  & (\all_features[1294]  | (\all_features[1293]  & (\all_features[1292]  | ~new_n14590_ | ~new_n14589_)));
  assign new_n14589_ = ~\all_features[1288]  & ~\all_features[1289] ;
  assign new_n14590_ = ~\all_features[1290]  & ~\all_features[1291] ;
  assign new_n14591_ = \all_features[1295]  & (\all_features[1294]  | (new_n14587_ & (\all_features[1290]  | \all_features[1291]  | \all_features[1289] )));
  assign new_n14592_ = ~\all_features[1293]  & \all_features[1294]  & \all_features[1295]  & (\all_features[1292]  ? new_n14590_ : (new_n14586_ | ~new_n14590_));
  assign new_n14593_ = \all_features[1295]  & (\all_features[1293]  | \all_features[1294]  | \all_features[1292] );
  assign new_n14594_ = new_n14595_ & (~\all_features[1293]  | (~\all_features[1292]  & (~\all_features[1291]  | (~\all_features[1290]  & ~\all_features[1289] ))));
  assign new_n14595_ = ~\all_features[1294]  & ~\all_features[1295] ;
  assign new_n14596_ = ~\all_features[1293]  & new_n14595_ & ((~\all_features[1290]  & new_n14589_) | ~\all_features[1292]  | ~\all_features[1291] );
  assign new_n14597_ = ~\all_features[1295]  & (~\all_features[1294]  | (~\all_features[1293]  & (new_n14589_ | ~new_n14585_ | ~\all_features[1292] )));
  assign new_n14598_ = new_n14595_ & (~\all_features[1291]  | ~new_n14587_ | (~\all_features[1290]  & ~new_n14586_));
  assign new_n14599_ = ~\all_features[1295]  & (~\all_features[1294]  | (~\all_features[1292]  & ~\all_features[1293]  & ~new_n14585_));
  assign new_n14600_ = new_n14605_ & (~new_n14606_ | (~new_n14601_ & ~new_n14597_ & ~new_n14599_));
  assign new_n14601_ = ~new_n14582_ & ~new_n14584_ & (~new_n14593_ | ~new_n14588_ | new_n14602_);
  assign new_n14602_ = new_n14591_ & new_n14603_ & (new_n14604_ | ~\all_features[1293]  | ~\all_features[1294]  | ~\all_features[1295] );
  assign new_n14603_ = \all_features[1294]  & \all_features[1295]  & (\all_features[1292]  | \all_features[1293]  | new_n14586_ | ~new_n14590_);
  assign new_n14604_ = ~\all_features[1291]  & ~\all_features[1292]  & (~\all_features[1290]  | new_n14589_);
  assign new_n14605_ = ~new_n14596_ & (\all_features[1291]  | \all_features[1292]  | \all_features[1293]  | \all_features[1294]  | \all_features[1295] );
  assign new_n14606_ = ~new_n14594_ & ~new_n14598_;
  assign new_n14607_ = new_n14608_ & new_n14605_ & ~new_n14598_ & ~new_n14597_ & ~new_n14582_ & ~new_n14594_;
  assign new_n14608_ = ~new_n14584_ & ~new_n14599_;
  assign new_n14609_ = new_n14605_ & new_n14606_ & (new_n14610_ | new_n14582_ | new_n14597_ | ~new_n14608_);
  assign new_n14610_ = new_n14593_ & new_n14603_ & new_n14588_ & new_n14591_;
  assign new_n14611_ = new_n14612_ & (~new_n14384_ | ~new_n14549_) & (~new_n14551_ | ~new_n14293_);
  assign new_n14612_ = (~new_n14576_ | ~new_n14578_) & (~new_n14158_ | ~new_n14577_);
  assign new_n14613_ = new_n14614_ & new_n14865_;
  assign new_n14614_ = new_n14615_ & (new_n14786_ | new_n14654_ | (new_n14812_ ? ~new_n14849_ : ~new_n14846_));
  assign new_n14615_ = new_n14616_ & (new_n14654_ | ~new_n14786_ | (new_n14783_ ? ~new_n14785_ : ~new_n13366_));
  assign new_n14616_ = ~new_n14654_ | (new_n14690_ ? (new_n14724_ ? ~new_n14725_ : ~new_n14759_) : new_n14617_);
  assign new_n14617_ = new_n14624_ ? ~new_n14618_ : new_n14626_;
  assign new_n14618_ = ~new_n14619_ & ~new_n14235_;
  assign new_n14619_ = new_n14212_ & new_n14620_ & new_n14237_;
  assign new_n14620_ = ~new_n14621_ & (\all_features[4371]  | \all_features[4372]  | \all_features[4373]  | \all_features[4374]  | \all_features[4375] );
  assign new_n14621_ = ~new_n14234_ & (new_n14232_ | (~new_n14230_ & (new_n14228_ | (~new_n14214_ & ~new_n14622_))));
  assign new_n14622_ = ~new_n14225_ & (new_n14227_ | (new_n14224_ & (~new_n14218_ | (~new_n14623_ & new_n14220_))));
  assign new_n14623_ = ~\all_features[4373]  & \all_features[4374]  & \all_features[4375]  & (\all_features[4372]  ? new_n14219_ : (new_n14223_ | ~new_n14219_));
  assign new_n14624_ = new_n14625_ & new_n13242_;
  assign new_n14625_ = new_n13238_ & new_n13210_;
  assign new_n14626_ = ~new_n14627_ & ~new_n14651_;
  assign new_n14627_ = ~new_n14650_ & ~new_n14649_ & ~new_n14648_ & ~new_n14628_ & ~new_n14646_;
  assign new_n14628_ = new_n14632_ & new_n14636_ & (~new_n14643_ | ~new_n14645_ | ~new_n14629_ | ~new_n14642_);
  assign new_n14629_ = \all_features[4847]  & (\all_features[4846]  | new_n14630_);
  assign new_n14630_ = \all_features[4845]  & (\all_features[4842]  | \all_features[4843]  | \all_features[4844]  | ~new_n14631_);
  assign new_n14631_ = ~\all_features[4840]  & ~\all_features[4841] ;
  assign new_n14632_ = ~new_n14633_ & ~new_n14635_;
  assign new_n14633_ = ~\all_features[4847]  & (~\all_features[4846]  | (~\all_features[4844]  & ~\all_features[4845]  & ~new_n14634_));
  assign new_n14634_ = \all_features[4842]  & \all_features[4843] ;
  assign new_n14635_ = ~\all_features[4847]  & (~\all_features[4846]  | (~\all_features[4845]  & (new_n14631_ | ~new_n14634_ | ~\all_features[4844] )));
  assign new_n14636_ = ~new_n14637_ & ~new_n14640_;
  assign new_n14637_ = ~\all_features[4847]  & (~\all_features[4846]  | ~new_n14638_ | ~new_n14639_ | ~new_n14634_);
  assign new_n14638_ = \all_features[4844]  & \all_features[4845] ;
  assign new_n14639_ = \all_features[4840]  & \all_features[4841] ;
  assign new_n14640_ = ~new_n14641_ & ~\all_features[4847] ;
  assign new_n14641_ = \all_features[4845]  & \all_features[4846]  & (\all_features[4844]  | (\all_features[4842]  & \all_features[4843]  & \all_features[4841] ));
  assign new_n14642_ = \all_features[4847]  & (\all_features[4846]  | (new_n14638_ & (\all_features[4842]  | \all_features[4843]  | \all_features[4841] )));
  assign new_n14643_ = new_n14644_ & (new_n14639_ | \all_features[4842]  | \all_features[4843]  | \all_features[4844]  | \all_features[4845] );
  assign new_n14644_ = \all_features[4846]  & \all_features[4847] ;
  assign new_n14645_ = \all_features[4847]  & (\all_features[4845]  | \all_features[4846]  | \all_features[4844] );
  assign new_n14646_ = new_n14647_ & (~\all_features[4845]  | (~\all_features[4844]  & (~\all_features[4843]  | (~\all_features[4842]  & ~\all_features[4841] ))));
  assign new_n14647_ = ~\all_features[4846]  & ~\all_features[4847] ;
  assign new_n14648_ = ~\all_features[4845]  & new_n14647_ & ((~\all_features[4842]  & new_n14631_) | ~\all_features[4844]  | ~\all_features[4843] );
  assign new_n14649_ = new_n14647_ & (~\all_features[4843]  | ~new_n14638_ | (~\all_features[4842]  & ~new_n14639_));
  assign new_n14650_ = ~\all_features[4847]  & ~\all_features[4846]  & ~\all_features[4845]  & ~\all_features[4843]  & ~\all_features[4844] ;
  assign new_n14651_ = new_n14653_ & new_n14652_ & ~new_n14648_ & ~new_n14640_ & ~new_n14633_ & ~new_n14635_;
  assign new_n14652_ = ~new_n14637_ & ~new_n14650_;
  assign new_n14653_ = ~new_n14646_ & ~new_n14649_;
  assign new_n14654_ = new_n14655_ & new_n14681_;
  assign new_n14655_ = ~new_n14656_ & ~new_n14679_;
  assign new_n14656_ = new_n14674_ & ~new_n14678_ & ~new_n14657_ & ~new_n14677_;
  assign new_n14657_ = ~new_n14672_ & ~new_n14673_ & new_n14665_ & (~new_n14670_ | ~new_n14658_);
  assign new_n14658_ = new_n14664_ & new_n14659_ & new_n14661_;
  assign new_n14659_ = \all_features[2111]  & (\all_features[2110]  | (new_n14660_ & (\all_features[2106]  | \all_features[2107]  | \all_features[2105] )));
  assign new_n14660_ = \all_features[2108]  & \all_features[2109] ;
  assign new_n14661_ = \all_features[2110]  & \all_features[2111]  & (\all_features[2108]  | \all_features[2109]  | new_n14663_ | ~new_n14662_);
  assign new_n14662_ = ~\all_features[2106]  & ~\all_features[2107] ;
  assign new_n14663_ = \all_features[2104]  & \all_features[2105] ;
  assign new_n14664_ = \all_features[2111]  & (\all_features[2109]  | \all_features[2110]  | \all_features[2108] );
  assign new_n14665_ = ~new_n14666_ & ~new_n14668_;
  assign new_n14666_ = ~new_n14667_ & ~\all_features[2111] ;
  assign new_n14667_ = \all_features[2109]  & \all_features[2110]  & (\all_features[2108]  | (\all_features[2106]  & \all_features[2107]  & \all_features[2105] ));
  assign new_n14668_ = ~\all_features[2111]  & (~\all_features[2110]  | (~\all_features[2108]  & ~\all_features[2109]  & ~new_n14669_));
  assign new_n14669_ = \all_features[2106]  & \all_features[2107] ;
  assign new_n14670_ = \all_features[2111]  & (\all_features[2110]  | (\all_features[2109]  & (\all_features[2108]  | ~new_n14671_ | ~new_n14662_)));
  assign new_n14671_ = ~\all_features[2104]  & ~\all_features[2105] ;
  assign new_n14672_ = ~\all_features[2111]  & (~\all_features[2110]  | (~\all_features[2109]  & (new_n14671_ | ~new_n14669_ | ~\all_features[2108] )));
  assign new_n14673_ = ~\all_features[2111]  & (~\all_features[2110]  | ~new_n14660_ | ~new_n14663_ | ~new_n14669_);
  assign new_n14674_ = ~new_n14675_ & (\all_features[2107]  | \all_features[2108]  | \all_features[2109]  | \all_features[2110]  | \all_features[2111] );
  assign new_n14675_ = ~\all_features[2109]  & new_n14676_ & ((~\all_features[2106]  & new_n14671_) | ~\all_features[2108]  | ~\all_features[2107] );
  assign new_n14676_ = ~\all_features[2110]  & ~\all_features[2111] ;
  assign new_n14677_ = new_n14676_ & (~\all_features[2109]  | (~\all_features[2108]  & (~\all_features[2107]  | (~\all_features[2106]  & ~\all_features[2105] ))));
  assign new_n14678_ = new_n14676_ & (~\all_features[2107]  | ~new_n14660_ | (~\all_features[2106]  & ~new_n14663_));
  assign new_n14679_ = new_n14674_ & new_n14665_ & new_n14680_ & ~new_n14672_ & ~new_n14673_;
  assign new_n14680_ = ~new_n14677_ & ~new_n14678_;
  assign new_n14681_ = ~new_n14682_ & ~new_n14686_;
  assign new_n14682_ = ~new_n14683_ & (\all_features[2107]  | \all_features[2108]  | \all_features[2109]  | \all_features[2110]  | \all_features[2111] );
  assign new_n14683_ = ~new_n14675_ & (new_n14677_ | (~new_n14678_ & (new_n14668_ | (~new_n14672_ & ~new_n14684_))));
  assign new_n14684_ = ~new_n14666_ & (new_n14673_ | (new_n14664_ & (~new_n14670_ | (~new_n14685_ & new_n14659_))));
  assign new_n14685_ = ~\all_features[2109]  & \all_features[2110]  & \all_features[2111]  & (\all_features[2108]  ? new_n14662_ : (new_n14663_ | ~new_n14662_));
  assign new_n14686_ = new_n14674_ & (~new_n14680_ | (~new_n14687_ & ~new_n14668_ & ~new_n14672_));
  assign new_n14687_ = ~new_n14673_ & ~new_n14666_ & (~new_n14664_ | ~new_n14670_ | new_n14688_);
  assign new_n14688_ = new_n14659_ & new_n14661_ & (new_n14689_ | ~\all_features[2109]  | ~\all_features[2110]  | ~\all_features[2111] );
  assign new_n14689_ = ~\all_features[2107]  & ~\all_features[2108]  & (~\all_features[2106]  | new_n14671_);
  assign new_n14690_ = new_n14691_ & ~new_n14720_ & ~new_n14723_;
  assign new_n14691_ = ~new_n14692_ & (new_n14714_ | (~new_n14717_ & ~new_n14713_));
  assign new_n14692_ = new_n14712_ & (~new_n14708_ | (~new_n14693_ & ~new_n14715_ & ~new_n14716_));
  assign new_n14693_ = ~new_n14705_ & ~new_n14703_ & (~new_n14707_ | ~new_n14702_ | new_n14694_);
  assign new_n14694_ = new_n14695_ & new_n14697_ & (new_n14700_ | ~\all_features[5013]  | ~\all_features[5014]  | ~\all_features[5015] );
  assign new_n14695_ = \all_features[5015]  & (\all_features[5014]  | (new_n14696_ & (\all_features[5010]  | \all_features[5011]  | \all_features[5009] )));
  assign new_n14696_ = \all_features[5012]  & \all_features[5013] ;
  assign new_n14697_ = \all_features[5014]  & \all_features[5015]  & (\all_features[5012]  | \all_features[5013]  | new_n14698_ | ~new_n14699_);
  assign new_n14698_ = \all_features[5008]  & \all_features[5009] ;
  assign new_n14699_ = ~\all_features[5010]  & ~\all_features[5011] ;
  assign new_n14700_ = ~\all_features[5011]  & ~\all_features[5012]  & (~\all_features[5010]  | new_n14701_);
  assign new_n14701_ = ~\all_features[5008]  & ~\all_features[5009] ;
  assign new_n14702_ = \all_features[5015]  & (\all_features[5014]  | (\all_features[5013]  & (\all_features[5012]  | ~new_n14701_ | ~new_n14699_)));
  assign new_n14703_ = ~\all_features[5015]  & (~\all_features[5014]  | ~new_n14698_ | ~new_n14696_ | ~new_n14704_);
  assign new_n14704_ = \all_features[5010]  & \all_features[5011] ;
  assign new_n14705_ = ~new_n14706_ & ~\all_features[5015] ;
  assign new_n14706_ = \all_features[5013]  & \all_features[5014]  & (\all_features[5012]  | (\all_features[5010]  & \all_features[5011]  & \all_features[5009] ));
  assign new_n14707_ = \all_features[5015]  & (\all_features[5013]  | \all_features[5014]  | \all_features[5012] );
  assign new_n14708_ = ~new_n14709_ & ~new_n14711_;
  assign new_n14709_ = new_n14710_ & (~\all_features[5011]  | ~new_n14696_ | (~\all_features[5010]  & ~new_n14698_));
  assign new_n14710_ = ~\all_features[5014]  & ~\all_features[5015] ;
  assign new_n14711_ = new_n14710_ & (~\all_features[5013]  | (~\all_features[5012]  & (~\all_features[5011]  | (~\all_features[5010]  & ~\all_features[5009] ))));
  assign new_n14712_ = ~new_n14713_ & ~new_n14714_;
  assign new_n14713_ = ~\all_features[5013]  & new_n14710_ & ((~\all_features[5010]  & new_n14701_) | ~\all_features[5012]  | ~\all_features[5011] );
  assign new_n14714_ = ~\all_features[5015]  & ~\all_features[5014]  & ~\all_features[5013]  & ~\all_features[5011]  & ~\all_features[5012] ;
  assign new_n14715_ = ~\all_features[5015]  & (~\all_features[5014]  | (~\all_features[5012]  & ~\all_features[5013]  & ~new_n14704_));
  assign new_n14716_ = ~\all_features[5015]  & (~\all_features[5014]  | (~\all_features[5013]  & (new_n14701_ | ~new_n14704_ | ~\all_features[5012] )));
  assign new_n14717_ = ~new_n14711_ & (new_n14709_ | (~new_n14715_ & (new_n14716_ | (~new_n14705_ & ~new_n14718_))));
  assign new_n14718_ = ~new_n14703_ & (~new_n14707_ | (new_n14702_ & (~new_n14695_ | (~new_n14719_ & new_n14697_))));
  assign new_n14719_ = \all_features[5014]  & \all_features[5015]  & (\all_features[5013]  | (~new_n14699_ & \all_features[5012] ));
  assign new_n14720_ = new_n14708_ & new_n14712_ & (new_n14721_ | new_n14703_ | new_n14716_ | ~new_n14722_);
  assign new_n14721_ = new_n14707_ & new_n14702_ & new_n14695_ & new_n14697_;
  assign new_n14722_ = ~new_n14705_ & ~new_n14715_;
  assign new_n14723_ = new_n14712_ & new_n14708_ & new_n14722_ & ~new_n14703_ & ~new_n14716_;
  assign new_n14724_ = new_n7136_ & new_n13356_;
  assign new_n14725_ = new_n14726_ & (~new_n14755_ | ~new_n14751_);
  assign new_n14726_ = ~new_n14727_ & ~new_n14749_;
  assign new_n14727_ = new_n14744_ & ~new_n14748_ & ~new_n14728_ & ~new_n14747_;
  assign new_n14728_ = new_n14729_ & (~new_n14742_ | ~new_n14743_ | ~new_n14739_ | ~new_n14741_);
  assign new_n14729_ = ~new_n14738_ & ~new_n14735_ & ~new_n14730_ & ~new_n14733_;
  assign new_n14730_ = ~\all_features[4535]  & (~\all_features[4534]  | (~\all_features[4533]  & (new_n14731_ | ~new_n14732_ | ~\all_features[4532] )));
  assign new_n14731_ = ~\all_features[4528]  & ~\all_features[4529] ;
  assign new_n14732_ = \all_features[4530]  & \all_features[4531] ;
  assign new_n14733_ = ~new_n14734_ & ~\all_features[4535] ;
  assign new_n14734_ = \all_features[4533]  & \all_features[4534]  & (\all_features[4532]  | (\all_features[4530]  & \all_features[4531]  & \all_features[4529] ));
  assign new_n14735_ = ~\all_features[4535]  & (~\all_features[4534]  | ~new_n14736_ | ~new_n14737_ | ~new_n14732_);
  assign new_n14736_ = \all_features[4532]  & \all_features[4533] ;
  assign new_n14737_ = \all_features[4528]  & \all_features[4529] ;
  assign new_n14738_ = ~\all_features[4535]  & (~\all_features[4534]  | (~\all_features[4532]  & ~\all_features[4533]  & ~new_n14732_));
  assign new_n14739_ = \all_features[4535]  & (\all_features[4534]  | (\all_features[4533]  & (\all_features[4532]  | ~new_n14731_ | ~new_n14740_)));
  assign new_n14740_ = ~\all_features[4530]  & ~\all_features[4531] ;
  assign new_n14741_ = \all_features[4535]  & (\all_features[4534]  | (new_n14736_ & (\all_features[4530]  | \all_features[4531]  | \all_features[4529] )));
  assign new_n14742_ = \all_features[4534]  & \all_features[4535]  & (\all_features[4532]  | \all_features[4533]  | new_n14737_ | ~new_n14740_);
  assign new_n14743_ = \all_features[4535]  & (\all_features[4533]  | \all_features[4534]  | \all_features[4532] );
  assign new_n14744_ = ~new_n14745_ & (\all_features[4531]  | \all_features[4532]  | \all_features[4533]  | \all_features[4534]  | \all_features[4535] );
  assign new_n14745_ = ~\all_features[4533]  & new_n14746_ & ((~\all_features[4530]  & new_n14731_) | ~\all_features[4532]  | ~\all_features[4531] );
  assign new_n14746_ = ~\all_features[4534]  & ~\all_features[4535] ;
  assign new_n14747_ = new_n14746_ & (~\all_features[4533]  | (~\all_features[4532]  & (~\all_features[4531]  | (~\all_features[4530]  & ~\all_features[4529] ))));
  assign new_n14748_ = new_n14746_ & (~\all_features[4531]  | ~new_n14736_ | (~\all_features[4530]  & ~new_n14737_));
  assign new_n14749_ = new_n14750_ & new_n14744_ & ~new_n14733_ & ~new_n14747_;
  assign new_n14750_ = ~new_n14748_ & ~new_n14738_ & ~new_n14730_ & ~new_n14735_;
  assign new_n14751_ = new_n14744_ & (new_n14748_ | new_n14747_ | (~new_n14730_ & ~new_n14738_ & ~new_n14752_));
  assign new_n14752_ = ~new_n14735_ & ~new_n14733_ & (~new_n14743_ | ~new_n14739_ | new_n14753_);
  assign new_n14753_ = new_n14741_ & new_n14742_ & (new_n14754_ | ~\all_features[4533]  | ~\all_features[4534]  | ~\all_features[4535] );
  assign new_n14754_ = ~\all_features[4531]  & ~\all_features[4532]  & (~\all_features[4530]  | new_n14731_);
  assign new_n14755_ = ~new_n14756_ & (\all_features[4531]  | \all_features[4532]  | \all_features[4533]  | \all_features[4534]  | \all_features[4535] );
  assign new_n14756_ = ~new_n14745_ & (new_n14747_ | (~new_n14748_ & (new_n14738_ | (~new_n14730_ & ~new_n14757_))));
  assign new_n14757_ = ~new_n14733_ & (new_n14735_ | (new_n14743_ & (~new_n14739_ | (~new_n14758_ & new_n14741_))));
  assign new_n14758_ = ~\all_features[4533]  & \all_features[4534]  & \all_features[4535]  & (\all_features[4532]  ? new_n14740_ : (new_n14737_ | ~new_n14740_));
  assign new_n14759_ = ~new_n14760_ & ~new_n14782_;
  assign new_n14760_ = new_n14761_ & (~new_n14770_ | (new_n14780_ & new_n14781_ & new_n14777_ & new_n14779_));
  assign new_n14761_ = new_n14762_ & ~new_n14766_ & ~new_n14767_;
  assign new_n14762_ = ~new_n14763_ & (\all_features[1427]  | \all_features[1428]  | \all_features[1429]  | \all_features[1430]  | \all_features[1431] );
  assign new_n14763_ = ~\all_features[1429]  & new_n14765_ & ((~\all_features[1426]  & new_n14764_) | ~\all_features[1428]  | ~\all_features[1427] );
  assign new_n14764_ = ~\all_features[1424]  & ~\all_features[1425] ;
  assign new_n14765_ = ~\all_features[1430]  & ~\all_features[1431] ;
  assign new_n14766_ = new_n14765_ & (~\all_features[1429]  | (~\all_features[1428]  & (~\all_features[1427]  | (~\all_features[1426]  & ~\all_features[1425] ))));
  assign new_n14767_ = new_n14765_ & (~\all_features[1427]  | ~new_n14768_ | (~\all_features[1426]  & ~new_n14769_));
  assign new_n14768_ = \all_features[1428]  & \all_features[1429] ;
  assign new_n14769_ = \all_features[1424]  & \all_features[1425] ;
  assign new_n14770_ = ~new_n14776_ & ~new_n14775_ & ~new_n14771_ & ~new_n14773_;
  assign new_n14771_ = ~\all_features[1431]  & (~\all_features[1430]  | (~\all_features[1429]  & (new_n14764_ | ~new_n14772_ | ~\all_features[1428] )));
  assign new_n14772_ = \all_features[1426]  & \all_features[1427] ;
  assign new_n14773_ = ~new_n14774_ & ~\all_features[1431] ;
  assign new_n14774_ = \all_features[1429]  & \all_features[1430]  & (\all_features[1428]  | (\all_features[1426]  & \all_features[1427]  & \all_features[1425] ));
  assign new_n14775_ = ~\all_features[1431]  & (~\all_features[1430]  | ~new_n14768_ | ~new_n14769_ | ~new_n14772_);
  assign new_n14776_ = ~\all_features[1431]  & (~\all_features[1430]  | (~\all_features[1428]  & ~\all_features[1429]  & ~new_n14772_));
  assign new_n14777_ = \all_features[1431]  & (\all_features[1430]  | (\all_features[1429]  & (\all_features[1428]  | ~new_n14764_ | ~new_n14778_)));
  assign new_n14778_ = ~\all_features[1426]  & ~\all_features[1427] ;
  assign new_n14779_ = \all_features[1431]  & (\all_features[1430]  | (new_n14768_ & (\all_features[1426]  | \all_features[1427]  | \all_features[1425] )));
  assign new_n14780_ = \all_features[1430]  & \all_features[1431]  & (\all_features[1428]  | \all_features[1429]  | new_n14769_ | ~new_n14778_);
  assign new_n14781_ = \all_features[1431]  & (\all_features[1429]  | \all_features[1430]  | \all_features[1428] );
  assign new_n14782_ = new_n14761_ & new_n14770_;
  assign new_n14783_ = ~new_n14154_ & (~new_n14156_ | new_n14784_);
  assign new_n14784_ = ~new_n14126_ & ~new_n14147_;
  assign new_n14785_ = ~new_n6698_ & (~new_n6675_ | new_n14540_);
  assign new_n14786_ = new_n14787_ & new_n14810_;
  assign new_n14787_ = new_n14805_ & ~new_n14809_ & ~new_n14788_ & ~new_n14808_;
  assign new_n14788_ = ~new_n14803_ & ~new_n14804_ & new_n14796_ & (~new_n14801_ | ~new_n14789_);
  assign new_n14789_ = new_n14795_ & new_n14790_ & new_n14792_;
  assign new_n14790_ = \all_features[4591]  & (\all_features[4590]  | (new_n14791_ & (\all_features[4586]  | \all_features[4587]  | \all_features[4585] )));
  assign new_n14791_ = \all_features[4588]  & \all_features[4589] ;
  assign new_n14792_ = \all_features[4590]  & \all_features[4591]  & (\all_features[4588]  | \all_features[4589]  | new_n14794_ | ~new_n14793_);
  assign new_n14793_ = ~\all_features[4586]  & ~\all_features[4587] ;
  assign new_n14794_ = \all_features[4584]  & \all_features[4585] ;
  assign new_n14795_ = \all_features[4591]  & (\all_features[4589]  | \all_features[4590]  | \all_features[4588] );
  assign new_n14796_ = ~new_n14797_ & ~new_n14799_;
  assign new_n14797_ = ~new_n14798_ & ~\all_features[4591] ;
  assign new_n14798_ = \all_features[4589]  & \all_features[4590]  & (\all_features[4588]  | (\all_features[4586]  & \all_features[4587]  & \all_features[4585] ));
  assign new_n14799_ = ~\all_features[4591]  & (~\all_features[4590]  | (~\all_features[4588]  & ~\all_features[4589]  & ~new_n14800_));
  assign new_n14800_ = \all_features[4586]  & \all_features[4587] ;
  assign new_n14801_ = \all_features[4591]  & (\all_features[4590]  | (\all_features[4589]  & (\all_features[4588]  | ~new_n14802_ | ~new_n14793_)));
  assign new_n14802_ = ~\all_features[4584]  & ~\all_features[4585] ;
  assign new_n14803_ = ~\all_features[4591]  & (~\all_features[4590]  | (~\all_features[4589]  & (new_n14802_ | ~new_n14800_ | ~\all_features[4588] )));
  assign new_n14804_ = ~\all_features[4591]  & (~\all_features[4590]  | ~new_n14791_ | ~new_n14794_ | ~new_n14800_);
  assign new_n14805_ = ~new_n14806_ & (\all_features[4587]  | \all_features[4588]  | \all_features[4589]  | \all_features[4590]  | \all_features[4591] );
  assign new_n14806_ = ~\all_features[4589]  & new_n14807_ & ((~\all_features[4586]  & new_n14802_) | ~\all_features[4588]  | ~\all_features[4587] );
  assign new_n14807_ = ~\all_features[4590]  & ~\all_features[4591] ;
  assign new_n14808_ = new_n14807_ & (~\all_features[4589]  | (~\all_features[4588]  & (~\all_features[4587]  | (~\all_features[4586]  & ~\all_features[4585] ))));
  assign new_n14809_ = new_n14807_ & (~\all_features[4587]  | ~new_n14791_ | (~\all_features[4586]  & ~new_n14794_));
  assign new_n14810_ = new_n14805_ & new_n14796_ & new_n14811_ & ~new_n14803_ & ~new_n14804_;
  assign new_n14811_ = ~new_n14808_ & ~new_n14809_;
  assign new_n14812_ = ~new_n14845_ & (~new_n14843_ | new_n14813_);
  assign new_n14813_ = ~new_n14814_ & ~new_n14834_;
  assign new_n14814_ = ~new_n14833_ & (new_n14828_ | (~new_n14830_ & (new_n14831_ | (~new_n14815_ & ~new_n14832_))));
  assign new_n14815_ = ~new_n14822_ & (new_n14825_ | (~new_n14824_ & (~new_n14827_ | new_n14816_)));
  assign new_n14816_ = \all_features[1439]  & ((~new_n14821_ & ~\all_features[1437]  & \all_features[1438] ) | (~new_n14819_ & (\all_features[1438]  | (~new_n14817_ & \all_features[1437] ))));
  assign new_n14817_ = new_n14818_ & ~\all_features[1436]  & ~\all_features[1434]  & ~\all_features[1435] ;
  assign new_n14818_ = ~\all_features[1432]  & ~\all_features[1433] ;
  assign new_n14819_ = \all_features[1439]  & (\all_features[1438]  | (new_n14820_ & (\all_features[1434]  | \all_features[1435]  | \all_features[1433] )));
  assign new_n14820_ = \all_features[1436]  & \all_features[1437] ;
  assign new_n14821_ = (~\all_features[1434]  & ~\all_features[1435]  & ~\all_features[1436]  & (~\all_features[1433]  | ~\all_features[1432] )) | (\all_features[1436]  & (\all_features[1434]  | \all_features[1435] ));
  assign new_n14822_ = ~\all_features[1439]  & (~\all_features[1438]  | (~\all_features[1437]  & (new_n14818_ | ~new_n14823_ | ~\all_features[1436] )));
  assign new_n14823_ = \all_features[1434]  & \all_features[1435] ;
  assign new_n14824_ = ~\all_features[1439]  & (~new_n14823_ | ~\all_features[1432]  | ~\all_features[1433]  | ~\all_features[1438]  | ~new_n14820_);
  assign new_n14825_ = ~new_n14826_ & ~\all_features[1439] ;
  assign new_n14826_ = \all_features[1437]  & \all_features[1438]  & (\all_features[1436]  | (\all_features[1434]  & \all_features[1435]  & \all_features[1433] ));
  assign new_n14827_ = \all_features[1439]  & (\all_features[1437]  | \all_features[1438]  | \all_features[1436] );
  assign new_n14828_ = ~\all_features[1437]  & new_n14829_ & ((~\all_features[1434]  & new_n14818_) | ~\all_features[1436]  | ~\all_features[1435] );
  assign new_n14829_ = ~\all_features[1438]  & ~\all_features[1439] ;
  assign new_n14830_ = new_n14829_ & (~\all_features[1437]  | (~\all_features[1436]  & (~\all_features[1435]  | (~\all_features[1434]  & ~\all_features[1433] ))));
  assign new_n14831_ = new_n14829_ & (~new_n14820_ | ~\all_features[1435]  | (~\all_features[1434]  & (~\all_features[1432]  | ~\all_features[1433] )));
  assign new_n14832_ = ~\all_features[1439]  & (~\all_features[1438]  | (~\all_features[1436]  & ~\all_features[1437]  & ~new_n14823_));
  assign new_n14833_ = ~\all_features[1439]  & ~\all_features[1438]  & ~\all_features[1437]  & ~\all_features[1435]  & ~\all_features[1436] ;
  assign new_n14834_ = new_n14840_ & (~new_n14842_ | (~new_n14832_ & ~new_n14822_ & (~new_n14841_ | new_n14835_)));
  assign new_n14835_ = new_n14836_ & (~new_n14837_ | (~new_n14839_ & \all_features[1437]  & \all_features[1438]  & \all_features[1439] ));
  assign new_n14836_ = \all_features[1439]  & (\all_features[1438]  | (~new_n14817_ & \all_features[1437] ));
  assign new_n14837_ = \all_features[1439]  & \all_features[1438]  & ~new_n14838_ & new_n14819_;
  assign new_n14838_ = ~\all_features[1434]  & ~\all_features[1435]  & ~\all_features[1436]  & ~\all_features[1437]  & (~\all_features[1433]  | ~\all_features[1432] );
  assign new_n14839_ = ~\all_features[1435]  & ~\all_features[1436]  & (~\all_features[1434]  | new_n14818_);
  assign new_n14840_ = ~new_n14828_ & ~new_n14833_;
  assign new_n14841_ = ~new_n14824_ & ~new_n14825_;
  assign new_n14842_ = ~new_n14830_ & ~new_n14831_;
  assign new_n14843_ = new_n14842_ & ~new_n14844_ & new_n14840_;
  assign new_n14844_ = ~new_n14832_ & ~new_n14822_ & ~new_n14824_ & ~new_n14825_ & (~new_n14837_ | ~new_n14836_);
  assign new_n14845_ = new_n14841_ & new_n14840_ & ~new_n14822_ & ~new_n14832_ & ~new_n14830_ & ~new_n14831_;
  assign new_n14846_ = new_n14847_ & new_n14848_;
  assign new_n14847_ = ~new_n7988_ & ~new_n7991_;
  assign new_n14848_ = ~new_n7959_ & ~new_n7980_;
  assign new_n14849_ = new_n14854_ & new_n14850_ & ~new_n14864_ & ~new_n14863_ & ~new_n14860_ & ~new_n14862_;
  assign new_n14850_ = ~new_n14851_ & (\all_features[4859]  | \all_features[4860]  | \all_features[4861]  | \all_features[4862]  | \all_features[4863] );
  assign new_n14851_ = ~\all_features[4861]  & new_n14852_ & ((~\all_features[4858]  & new_n14853_) | ~\all_features[4860]  | ~\all_features[4859] );
  assign new_n14852_ = ~\all_features[4862]  & ~\all_features[4863] ;
  assign new_n14853_ = ~\all_features[4856]  & ~\all_features[4857] ;
  assign new_n14854_ = ~new_n14855_ & ~new_n14859_;
  assign new_n14855_ = ~\all_features[4863]  & (~\all_features[4862]  | ~new_n14856_ | ~new_n14857_ | ~new_n14858_);
  assign new_n14856_ = \all_features[4858]  & \all_features[4859] ;
  assign new_n14857_ = \all_features[4856]  & \all_features[4857] ;
  assign new_n14858_ = \all_features[4860]  & \all_features[4861] ;
  assign new_n14859_ = ~\all_features[4863]  & (~\all_features[4862]  | (~\all_features[4860]  & ~\all_features[4861]  & ~new_n14856_));
  assign new_n14860_ = ~new_n14861_ & ~\all_features[4863] ;
  assign new_n14861_ = \all_features[4861]  & \all_features[4862]  & (\all_features[4860]  | (\all_features[4858]  & \all_features[4859]  & \all_features[4857] ));
  assign new_n14862_ = new_n14852_ & (~\all_features[4861]  | (~\all_features[4860]  & (~\all_features[4859]  | (~\all_features[4858]  & ~\all_features[4857] ))));
  assign new_n14863_ = ~\all_features[4863]  & (~\all_features[4862]  | (~\all_features[4861]  & (new_n14853_ | ~new_n14856_ | ~\all_features[4860] )));
  assign new_n14864_ = new_n14852_ & (~\all_features[4859]  | ~new_n14858_ | (~\all_features[4858]  & ~new_n14857_));
  assign new_n14865_ = new_n14866_ & (new_n14786_ | new_n14654_ | (new_n14812_ ? new_n14849_ : new_n14846_));
  assign new_n14866_ = ~new_n14867_ & (~new_n14654_ | ((new_n14724_ | new_n14759_ | ~new_n14690_) & (new_n14868_ | new_n14690_)));
  assign new_n14867_ = ~new_n14654_ & new_n14786_ & (new_n14783_ ? ~new_n14785_ : ~new_n13366_);
  assign new_n14868_ = new_n14624_ ? new_n14618_ : ~new_n14626_;
  assign new_n14869_ = new_n14870_ ? (~new_n14613_ ^ new_n15211_) : (new_n14613_ ^ new_n15211_);
  assign new_n14870_ = new_n14871_ ? (new_n15025_ ^ new_n15149_) : (~new_n15025_ ^ new_n15149_);
  assign new_n14871_ = ~new_n14872_ & new_n15019_;
  assign new_n14872_ = new_n14873_ & (new_n15018_ | ~new_n14988_ | ~new_n14987_);
  assign new_n14873_ = ~new_n14917_ & (~new_n14874_ | (~new_n14922_ & new_n14953_) | (~new_n14986_ & ~new_n14953_));
  assign new_n14874_ = ~new_n14875_ & new_n14884_;
  assign new_n14875_ = new_n14876_ & new_n14883_;
  assign new_n14876_ = new_n14877_ & new_n11751_;
  assign new_n14877_ = ~new_n14878_ & (\all_features[4619]  | \all_features[4620]  | ~new_n11731_);
  assign new_n14878_ = ~new_n11730_ & (new_n11736_ | (~new_n11734_ & (new_n11747_ | new_n14879_)));
  assign new_n14879_ = ~new_n11745_ & (new_n11741_ | (~new_n11743_ & (~new_n14882_ | new_n14880_)));
  assign new_n14880_ = \all_features[4623]  & ((~new_n14881_ & ~\all_features[4621]  & \all_features[4622] ) | (~new_n11738_ & (\all_features[4622]  | (~new_n11749_ & \all_features[4621] ))));
  assign new_n14881_ = (~\all_features[4618]  & ~\all_features[4619]  & ~\all_features[4620]  & (~\all_features[4617]  | ~\all_features[4616] )) | (\all_features[4620]  & (\all_features[4618]  | \all_features[4619] ));
  assign new_n14882_ = \all_features[4623]  & (\all_features[4621]  | \all_features[4622]  | \all_features[4620] );
  assign new_n14883_ = new_n11727_ & new_n11750_;
  assign new_n14884_ = ~new_n14915_ & ~new_n14913_ & ~new_n14885_ & ~new_n14906_;
  assign new_n14885_ = ~new_n14886_ & (\all_features[2635]  | \all_features[2636]  | \all_features[2637]  | \all_features[2638]  | \all_features[2639] );
  assign new_n14886_ = ~new_n14900_ & (new_n14902_ | (~new_n14903_ & (new_n14904_ | (~new_n14887_ & ~new_n14905_))));
  assign new_n14887_ = ~new_n14888_ & (new_n14890_ | (new_n14899_ & (~new_n14894_ | (~new_n14898_ & new_n14897_))));
  assign new_n14888_ = ~new_n14889_ & ~\all_features[2639] ;
  assign new_n14889_ = \all_features[2637]  & \all_features[2638]  & (\all_features[2636]  | (\all_features[2634]  & \all_features[2635]  & \all_features[2633] ));
  assign new_n14890_ = ~\all_features[2639]  & (~\all_features[2638]  | ~new_n14891_ | ~new_n14892_ | ~new_n14893_);
  assign new_n14891_ = \all_features[2632]  & \all_features[2633] ;
  assign new_n14892_ = \all_features[2636]  & \all_features[2637] ;
  assign new_n14893_ = \all_features[2634]  & \all_features[2635] ;
  assign new_n14894_ = \all_features[2639]  & (\all_features[2638]  | (\all_features[2637]  & (\all_features[2636]  | ~new_n14896_ | ~new_n14895_)));
  assign new_n14895_ = ~\all_features[2632]  & ~\all_features[2633] ;
  assign new_n14896_ = ~\all_features[2634]  & ~\all_features[2635] ;
  assign new_n14897_ = \all_features[2639]  & (\all_features[2638]  | (new_n14892_ & (\all_features[2634]  | \all_features[2635]  | \all_features[2633] )));
  assign new_n14898_ = ~\all_features[2637]  & \all_features[2638]  & \all_features[2639]  & (\all_features[2636]  ? new_n14896_ : (new_n14891_ | ~new_n14896_));
  assign new_n14899_ = \all_features[2639]  & (\all_features[2637]  | \all_features[2638]  | \all_features[2636] );
  assign new_n14900_ = ~\all_features[2637]  & new_n14901_ & ((~\all_features[2634]  & new_n14895_) | ~\all_features[2636]  | ~\all_features[2635] );
  assign new_n14901_ = ~\all_features[2638]  & ~\all_features[2639] ;
  assign new_n14902_ = new_n14901_ & (~\all_features[2637]  | (~\all_features[2636]  & (~\all_features[2635]  | (~\all_features[2634]  & ~\all_features[2633] ))));
  assign new_n14903_ = new_n14901_ & (~\all_features[2635]  | ~new_n14892_ | (~\all_features[2634]  & ~new_n14891_));
  assign new_n14904_ = ~\all_features[2639]  & (~\all_features[2638]  | (~\all_features[2636]  & ~\all_features[2637]  & ~new_n14893_));
  assign new_n14905_ = ~\all_features[2639]  & (~\all_features[2638]  | (~\all_features[2637]  & (new_n14895_ | ~new_n14893_ | ~\all_features[2636] )));
  assign new_n14906_ = new_n14911_ & (~new_n14912_ | (~new_n14907_ & ~new_n14904_ & ~new_n14905_));
  assign new_n14907_ = ~new_n14888_ & ~new_n14890_ & (~new_n14899_ | ~new_n14894_ | new_n14908_);
  assign new_n14908_ = new_n14897_ & new_n14909_ & (new_n14910_ | ~\all_features[2637]  | ~\all_features[2638]  | ~\all_features[2639] );
  assign new_n14909_ = \all_features[2638]  & \all_features[2639]  & (\all_features[2636]  | \all_features[2637]  | new_n14891_ | ~new_n14896_);
  assign new_n14910_ = ~\all_features[2635]  & ~\all_features[2636]  & (~\all_features[2634]  | new_n14895_);
  assign new_n14911_ = ~new_n14900_ & (\all_features[2635]  | \all_features[2636]  | \all_features[2637]  | \all_features[2638]  | \all_features[2639] );
  assign new_n14912_ = ~new_n14902_ & ~new_n14903_;
  assign new_n14913_ = new_n14914_ & new_n14911_ & ~new_n14888_ & ~new_n14905_ & ~new_n14902_ & ~new_n14903_;
  assign new_n14914_ = ~new_n14904_ & ~new_n14890_;
  assign new_n14915_ = new_n14911_ & new_n14912_ & (new_n14916_ | new_n14905_ | new_n14888_ | ~new_n14914_);
  assign new_n14916_ = new_n14899_ & new_n14909_ & new_n14894_ & new_n14897_;
  assign new_n14917_ = new_n11337_ & new_n14921_ & ~new_n14918_ & ~new_n14884_;
  assign new_n14918_ = ~new_n12798_ & (~new_n14920_ | new_n14919_);
  assign new_n14919_ = ~new_n12229_ & ~new_n12794_;
  assign new_n14920_ = ~new_n12254_ & new_n12257_;
  assign new_n14921_ = ~new_n14264_ & ~new_n14273_;
  assign new_n14922_ = ~new_n14950_ & new_n14923_;
  assign new_n14923_ = ~new_n14924_ & ~new_n14947_;
  assign new_n14924_ = new_n14925_ & (new_n14944_ | new_n14945_ | ~new_n14940_ | (new_n14937_ & new_n14935_));
  assign new_n14925_ = new_n14926_ & new_n14932_;
  assign new_n14926_ = ~new_n14927_ & ~new_n14930_;
  assign new_n14927_ = ~\all_features[2334]  & ~\all_features[2335]  & (~\all_features[2331]  | ~new_n14929_ | (~\all_features[2330]  & ~new_n14928_));
  assign new_n14928_ = \all_features[2328]  & \all_features[2329] ;
  assign new_n14929_ = \all_features[2332]  & \all_features[2333] ;
  assign new_n14930_ = ~\all_features[2335]  & ~new_n14931_ & ~\all_features[2334] ;
  assign new_n14931_ = \all_features[2333]  & (\all_features[2332]  | (\all_features[2331]  & (\all_features[2330]  | \all_features[2329] )));
  assign new_n14932_ = ~new_n14934_ | (\all_features[2331]  & \all_features[2332]  & (\all_features[2330]  | ~new_n14933_));
  assign new_n14933_ = ~\all_features[2328]  & ~\all_features[2329] ;
  assign new_n14934_ = ~\all_features[2335]  & ~\all_features[2333]  & ~\all_features[2334] ;
  assign new_n14935_ = \all_features[2335]  & (\all_features[2334]  | (~new_n14936_ & \all_features[2333] ));
  assign new_n14936_ = new_n14933_ & ~\all_features[2332]  & ~\all_features[2330]  & ~\all_features[2331] ;
  assign new_n14937_ = \all_features[2335]  & \all_features[2334]  & ~new_n14939_ & new_n14938_;
  assign new_n14938_ = \all_features[2335]  & (\all_features[2334]  | (new_n14929_ & (\all_features[2330]  | \all_features[2331]  | \all_features[2329] )));
  assign new_n14939_ = ~\all_features[2333]  & ~\all_features[2332]  & ~\all_features[2331]  & ~new_n14928_ & ~\all_features[2330] ;
  assign new_n14940_ = ~new_n14941_ & ~new_n14943_;
  assign new_n14941_ = ~\all_features[2335]  & (~\all_features[2334]  | (~\all_features[2332]  & ~\all_features[2333]  & ~new_n14942_));
  assign new_n14942_ = \all_features[2330]  & \all_features[2331] ;
  assign new_n14943_ = ~\all_features[2335]  & (~\all_features[2334]  | ~new_n14928_ | ~new_n14929_ | ~new_n14942_);
  assign new_n14944_ = ~\all_features[2335]  & (~\all_features[2334]  | (~\all_features[2333]  & (new_n14933_ | ~new_n14942_ | ~\all_features[2332] )));
  assign new_n14945_ = ~new_n14946_ & ~\all_features[2335] ;
  assign new_n14946_ = \all_features[2333]  & \all_features[2334]  & (\all_features[2332]  | (\all_features[2330]  & \all_features[2331]  & \all_features[2329] ));
  assign new_n14947_ = new_n14949_ & new_n14925_ & new_n14948_;
  assign new_n14948_ = ~new_n14941_ & ~new_n14944_;
  assign new_n14949_ = ~new_n14943_ & ~new_n14945_;
  assign new_n14950_ = new_n14932_ & (~new_n14926_ | (new_n14948_ & (~new_n14949_ | new_n14951_)));
  assign new_n14951_ = new_n14935_ & (~new_n14937_ | (~new_n14952_ & \all_features[2333]  & \all_features[2334]  & \all_features[2335] ));
  assign new_n14952_ = ~\all_features[2331]  & ~\all_features[2332]  & (~\all_features[2330]  | new_n14933_);
  assign new_n14953_ = ~new_n14985_ & new_n14954_;
  assign new_n14954_ = ~new_n14955_ & ~new_n14980_;
  assign new_n14955_ = new_n14977_ & ~new_n14956_ & new_n14973_;
  assign new_n14956_ = new_n14963_ & (~new_n14971_ | ~new_n14972_ | ~new_n14960_ | ~new_n14957_);
  assign new_n14957_ = \all_features[4167]  & (\all_features[4166]  | new_n14958_);
  assign new_n14958_ = \all_features[4165]  & (\all_features[4162]  | \all_features[4163]  | \all_features[4164]  | ~new_n14959_);
  assign new_n14959_ = ~\all_features[4160]  & ~\all_features[4161] ;
  assign new_n14960_ = \all_features[4167]  & ~new_n14961_ & \all_features[4166] ;
  assign new_n14961_ = ~\all_features[4165]  & ~\all_features[4164]  & ~\all_features[4163]  & ~new_n14962_ & ~\all_features[4162] ;
  assign new_n14962_ = \all_features[4160]  & \all_features[4161] ;
  assign new_n14963_ = ~new_n14969_ & ~new_n14967_ & ~new_n14964_ & ~new_n14966_;
  assign new_n14964_ = ~\all_features[4167]  & (~\all_features[4166]  | (~\all_features[4164]  & ~\all_features[4165]  & ~new_n14965_));
  assign new_n14965_ = \all_features[4162]  & \all_features[4163] ;
  assign new_n14966_ = ~\all_features[4167]  & (~\all_features[4166]  | (~\all_features[4165]  & (new_n14959_ | ~\all_features[4164]  | ~new_n14965_)));
  assign new_n14967_ = ~new_n14968_ & ~\all_features[4167] ;
  assign new_n14968_ = \all_features[4165]  & \all_features[4166]  & (\all_features[4164]  | (\all_features[4162]  & \all_features[4163]  & \all_features[4161] ));
  assign new_n14969_ = ~\all_features[4167]  & (~\all_features[4166]  | ~new_n14965_ | ~new_n14962_ | ~new_n14970_);
  assign new_n14970_ = \all_features[4164]  & \all_features[4165] ;
  assign new_n14971_ = \all_features[4167]  & (\all_features[4166]  | (new_n14970_ & (\all_features[4162]  | \all_features[4163]  | \all_features[4161] )));
  assign new_n14972_ = \all_features[4167]  & (\all_features[4165]  | \all_features[4166]  | \all_features[4164] );
  assign new_n14973_ = ~new_n14974_ & ~new_n14976_;
  assign new_n14974_ = new_n14975_ & (~\all_features[4163]  | ~new_n14970_ | (~\all_features[4162]  & ~new_n14962_));
  assign new_n14975_ = ~\all_features[4166]  & ~\all_features[4167] ;
  assign new_n14976_ = new_n14975_ & (~\all_features[4165]  | (~\all_features[4164]  & (~\all_features[4163]  | (~\all_features[4162]  & ~\all_features[4161] ))));
  assign new_n14977_ = ~new_n14978_ & ~new_n14979_;
  assign new_n14978_ = ~\all_features[4165]  & new_n14975_ & ((~\all_features[4162]  & new_n14959_) | ~\all_features[4164]  | ~\all_features[4163] );
  assign new_n14979_ = ~\all_features[4167]  & ~\all_features[4166]  & ~\all_features[4165]  & ~\all_features[4163]  & ~\all_features[4164] ;
  assign new_n14980_ = new_n14977_ & (~new_n14973_ | (new_n14984_ & (new_n14981_ | new_n14967_ | new_n14969_)));
  assign new_n14981_ = new_n14972_ & ~new_n14982_ & new_n14957_;
  assign new_n14982_ = ~new_n14961_ & new_n14971_ & \all_features[4166]  & \all_features[4167]  & (~\all_features[4165]  | new_n14983_);
  assign new_n14983_ = ~\all_features[4163]  & ~\all_features[4164]  & (~\all_features[4162]  | new_n14959_);
  assign new_n14984_ = ~new_n14964_ & ~new_n14966_;
  assign new_n14985_ = new_n14973_ & new_n14984_ & ~new_n14979_ & ~new_n14969_ & ~new_n14967_ & ~new_n14978_;
  assign new_n14986_ = new_n14619_ & new_n14235_;
  assign new_n14987_ = new_n14875_ & new_n14884_;
  assign new_n14988_ = ~new_n14989_ & new_n15017_;
  assign new_n14989_ = ~new_n14990_ & ~new_n15013_;
  assign new_n14990_ = new_n15010_ & ~new_n14991_ & new_n15005_;
  assign new_n14991_ = ~new_n14999_ & ~new_n15001_ & ~new_n15002_ & ~new_n15004_ & (~new_n14995_ | ~new_n14992_);
  assign new_n14992_ = \all_features[791]  & (\all_features[790]  | (~new_n14993_ & \all_features[789] ));
  assign new_n14993_ = new_n14994_ & ~\all_features[788]  & ~\all_features[786]  & ~\all_features[787] ;
  assign new_n14994_ = ~\all_features[784]  & ~\all_features[785] ;
  assign new_n14995_ = \all_features[791]  & \all_features[790]  & ~new_n14998_ & new_n14996_;
  assign new_n14996_ = \all_features[791]  & (\all_features[790]  | (new_n14997_ & (\all_features[786]  | \all_features[787]  | \all_features[785] )));
  assign new_n14997_ = \all_features[788]  & \all_features[789] ;
  assign new_n14998_ = ~\all_features[786]  & ~\all_features[787]  & ~\all_features[788]  & ~\all_features[789]  & (~\all_features[785]  | ~\all_features[784] );
  assign new_n14999_ = ~\all_features[791]  & (~\all_features[790]  | (~\all_features[788]  & ~\all_features[789]  & ~new_n15000_));
  assign new_n15000_ = \all_features[786]  & \all_features[787] ;
  assign new_n15001_ = ~\all_features[791]  & (~\all_features[790]  | (~\all_features[789]  & (new_n14994_ | ~\all_features[788]  | ~new_n15000_)));
  assign new_n15002_ = ~new_n15003_ & ~\all_features[791] ;
  assign new_n15003_ = \all_features[789]  & \all_features[790]  & (\all_features[788]  | (\all_features[786]  & \all_features[787]  & \all_features[785] ));
  assign new_n15004_ = ~\all_features[791]  & (~new_n14997_ | ~\all_features[784]  | ~\all_features[785]  | ~\all_features[790]  | ~new_n15000_);
  assign new_n15005_ = ~new_n15006_ & ~new_n15009_;
  assign new_n15006_ = new_n15007_ & ((~\all_features[786]  & new_n14994_) | ~\all_features[788]  | ~\all_features[787] );
  assign new_n15007_ = ~\all_features[789]  & new_n15008_;
  assign new_n15008_ = ~\all_features[790]  & ~\all_features[791] ;
  assign new_n15009_ = new_n15007_ & ~\all_features[787]  & ~\all_features[788] ;
  assign new_n15010_ = ~new_n15011_ & ~new_n15012_;
  assign new_n15011_ = new_n15008_ & (~new_n14997_ | ~\all_features[787]  | (~\all_features[786]  & (~\all_features[784]  | ~\all_features[785] )));
  assign new_n15012_ = new_n15008_ & (~\all_features[789]  | (~\all_features[788]  & (~\all_features[787]  | (~\all_features[786]  & ~\all_features[785] ))));
  assign new_n15013_ = new_n15005_ & (~new_n15010_ | (new_n15016_ & (new_n15014_ | new_n15002_ | new_n15004_)));
  assign new_n15014_ = new_n14992_ & (~new_n14995_ | (~new_n15015_ & \all_features[789]  & \all_features[790]  & \all_features[791] ));
  assign new_n15015_ = ~\all_features[787]  & ~\all_features[788]  & (~\all_features[786]  | new_n14994_);
  assign new_n15016_ = ~new_n14999_ & ~new_n15001_;
  assign new_n15017_ = new_n15010_ & new_n15016_ & ~new_n15004_ & ~new_n15002_ & ~new_n15006_ & ~new_n15009_;
  assign new_n15018_ = new_n8701_ & (new_n8698_ | ~new_n8668_);
  assign new_n15019_ = ~new_n15020_ & new_n15021_ & (~new_n14987_ | (new_n14988_ & ~new_n15018_) | (~new_n15024_ & new_n15018_));
  assign new_n15020_ = new_n14874_ & (new_n14953_ ? ~new_n14922_ : ~new_n14986_);
  assign new_n15021_ = new_n14884_ | (~new_n14918_ & new_n11337_ & new_n14921_) | (new_n15022_ & ~new_n14921_);
  assign new_n15022_ = new_n15023_ & ~new_n9686_ & ~new_n9679_;
  assign new_n15023_ = ~new_n9682_ & ~new_n9655_;
  assign new_n15024_ = new_n12442_ & (new_n12439_ | ~new_n12409_);
  assign new_n15025_ = ~new_n15026_ & new_n15111_;
  assign new_n15026_ = ~new_n15105_ & new_n15027_;
  assign new_n15027_ = new_n15028_ & (~new_n15085_ | ~new_n15087_ | ~new_n15088_) & (~new_n15084_ | ~new_n15086_);
  assign new_n15028_ = (~new_n15029_ | ~new_n15041_) & (~new_n15038_ | ~new_n15048_) & (new_n15047_ | ~new_n15035_);
  assign new_n15029_ = new_n15033_ & ~new_n15030_ & new_n15031_;
  assign new_n15030_ = ~new_n8022_ & new_n11168_;
  assign new_n15031_ = new_n10726_ & (new_n10703_ | new_n15032_);
  assign new_n15032_ = new_n10729_ & new_n10733_;
  assign new_n15033_ = ~new_n8192_ & new_n15034_;
  assign new_n15034_ = ~new_n8166_ & ~new_n8188_;
  assign new_n15035_ = ~new_n15036_ & ~new_n15030_ & ~new_n15033_;
  assign new_n15036_ = new_n14122_ & new_n15037_ & new_n14119_;
  assign new_n15037_ = new_n14091_ & new_n14115_;
  assign new_n15038_ = ~new_n15039_ & new_n15030_;
  assign new_n15039_ = new_n6805_ & new_n15040_;
  assign new_n15040_ = new_n6838_ & new_n6841_;
  assign new_n15041_ = ~new_n9340_ & (~new_n9314_ | ~new_n15042_);
  assign new_n15042_ = new_n9341_ & new_n15043_;
  assign new_n15043_ = ~new_n9334_ & (new_n9333_ | new_n15044_);
  assign new_n15044_ = ~new_n9329_ & (new_n9331_ | (~new_n9324_ & (new_n9325_ | (~new_n9317_ & ~new_n15045_))));
  assign new_n15045_ = ~new_n9319_ & (~new_n9339_ | (new_n9338_ & (~new_n9335_ | (~new_n15046_ & new_n9336_))));
  assign new_n15046_ = \all_features[2174]  & \all_features[2175]  & (\all_features[2173]  | (~new_n9337_ & \all_features[2172] ));
  assign new_n15047_ = new_n11236_ & (new_n11233_ | ~new_n11203_);
  assign new_n15048_ = ~new_n15049_ & new_n15078_;
  assign new_n15049_ = new_n15050_ & new_n15074_;
  assign new_n15050_ = new_n15065_ & (~new_n15070_ | (~new_n15068_ & ~new_n15051_ & ~new_n15073_));
  assign new_n15051_ = ~new_n15063_ & ~new_n15061_ & (~new_n15064_ | ~new_n15060_ | new_n15052_);
  assign new_n15052_ = new_n15053_ & new_n15055_ & (new_n15058_ | ~\all_features[5501]  | ~\all_features[5502]  | ~\all_features[5503] );
  assign new_n15053_ = \all_features[5503]  & (\all_features[5502]  | (new_n15054_ & (\all_features[5498]  | \all_features[5499]  | \all_features[5497] )));
  assign new_n15054_ = \all_features[5500]  & \all_features[5501] ;
  assign new_n15055_ = \all_features[5502]  & \all_features[5503]  & (\all_features[5500]  | \all_features[5501]  | new_n15057_ | ~new_n15056_);
  assign new_n15056_ = ~\all_features[5498]  & ~\all_features[5499] ;
  assign new_n15057_ = \all_features[5496]  & \all_features[5497] ;
  assign new_n15058_ = ~\all_features[5499]  & ~\all_features[5500]  & (~\all_features[5498]  | new_n15059_);
  assign new_n15059_ = ~\all_features[5496]  & ~\all_features[5497] ;
  assign new_n15060_ = \all_features[5503]  & (\all_features[5502]  | (\all_features[5501]  & (\all_features[5500]  | ~new_n15056_ | ~new_n15059_)));
  assign new_n15061_ = ~new_n15062_ & ~\all_features[5503] ;
  assign new_n15062_ = \all_features[5501]  & \all_features[5502]  & (\all_features[5500]  | (\all_features[5498]  & \all_features[5499]  & \all_features[5497] ));
  assign new_n15063_ = ~\all_features[5503]  & (~new_n15057_ | ~\all_features[5498]  | ~\all_features[5499]  | ~\all_features[5502]  | ~new_n15054_);
  assign new_n15064_ = \all_features[5503]  & (\all_features[5501]  | \all_features[5502]  | \all_features[5500] );
  assign new_n15065_ = ~new_n15066_ & (\all_features[5499]  | \all_features[5500]  | \all_features[5501]  | \all_features[5502]  | \all_features[5503] );
  assign new_n15066_ = ~\all_features[5501]  & new_n15067_ & ((~\all_features[5498]  & new_n15059_) | ~\all_features[5500]  | ~\all_features[5499] );
  assign new_n15067_ = ~\all_features[5502]  & ~\all_features[5503] ;
  assign new_n15068_ = ~\all_features[5503]  & (~\all_features[5502]  | new_n15069_);
  assign new_n15069_ = ~\all_features[5501]  & (new_n15059_ | ~\all_features[5499]  | ~\all_features[5500]  | ~\all_features[5498] );
  assign new_n15070_ = ~new_n15071_ & ~new_n15072_;
  assign new_n15071_ = new_n15067_ & (~\all_features[5501]  | (~\all_features[5500]  & (~\all_features[5499]  | (~\all_features[5498]  & ~\all_features[5497] ))));
  assign new_n15072_ = new_n15067_ & (~\all_features[5499]  | ~new_n15054_ | (~new_n15057_ & ~\all_features[5498] ));
  assign new_n15073_ = ~\all_features[5503]  & (~\all_features[5502]  | (~\all_features[5501]  & ~\all_features[5500]  & (~\all_features[5499]  | ~\all_features[5498] )));
  assign new_n15074_ = ~new_n15075_ & (\all_features[5499]  | \all_features[5500]  | \all_features[5501]  | \all_features[5502]  | \all_features[5503] );
  assign new_n15075_ = ~new_n15066_ & (new_n15071_ | (~new_n15072_ & (new_n15073_ | (~new_n15068_ & ~new_n15076_))));
  assign new_n15076_ = ~new_n15061_ & (new_n15063_ | (new_n15064_ & (~new_n15060_ | (~new_n15077_ & new_n15053_))));
  assign new_n15077_ = ~\all_features[5501]  & \all_features[5502]  & \all_features[5503]  & (\all_features[5500]  ? new_n15056_ : (new_n15057_ | ~new_n15056_));
  assign new_n15078_ = ~new_n15079_ & ~new_n15082_;
  assign new_n15079_ = new_n15070_ & ~new_n15080_ & new_n15065_;
  assign new_n15080_ = ~new_n15073_ & ~new_n15063_ & ~new_n15061_ & ~new_n15068_ & ~new_n15081_;
  assign new_n15081_ = new_n15064_ & new_n15060_ & new_n15053_ & new_n15055_;
  assign new_n15082_ = new_n15065_ & new_n15083_ & ~new_n15061_ & ~new_n15071_;
  assign new_n15083_ = ~new_n15073_ & ~new_n15072_ & ~new_n15068_ & ~new_n15063_;
  assign new_n15084_ = ~new_n15048_ & new_n15038_;
  assign new_n15085_ = new_n15030_ & new_n15039_;
  assign new_n15086_ = ~new_n11820_ & ~new_n11823_;
  assign new_n15087_ = new_n10906_ & (new_n10908_ | new_n10899_);
  assign new_n15088_ = new_n15094_ & new_n15089_ & ~new_n15104_ & ~new_n15103_ & ~new_n15101_ & ~new_n15102_;
  assign new_n15089_ = ~new_n15090_ & ~new_n15093_;
  assign new_n15090_ = ~\all_features[1501]  & new_n15092_ & ((~\all_features[1498]  & new_n15091_) | ~\all_features[1500]  | ~\all_features[1499] );
  assign new_n15091_ = ~\all_features[1496]  & ~\all_features[1497] ;
  assign new_n15092_ = ~\all_features[1502]  & ~\all_features[1503] ;
  assign new_n15093_ = ~\all_features[1503]  & ~\all_features[1502]  & ~\all_features[1501]  & ~\all_features[1499]  & ~\all_features[1500] ;
  assign new_n15094_ = ~new_n15095_ & ~new_n15097_;
  assign new_n15095_ = ~new_n15096_ & ~\all_features[1503] ;
  assign new_n15096_ = \all_features[1501]  & \all_features[1502]  & (\all_features[1500]  | (\all_features[1498]  & \all_features[1499]  & \all_features[1497] ));
  assign new_n15097_ = ~\all_features[1503]  & (~\all_features[1502]  | ~new_n15098_ | ~new_n15099_ | ~new_n15100_);
  assign new_n15098_ = \all_features[1500]  & \all_features[1501] ;
  assign new_n15099_ = \all_features[1496]  & \all_features[1497] ;
  assign new_n15100_ = \all_features[1498]  & \all_features[1499] ;
  assign new_n15101_ = ~\all_features[1503]  & (~\all_features[1502]  | (~\all_features[1500]  & ~\all_features[1501]  & ~new_n15100_));
  assign new_n15102_ = ~\all_features[1503]  & (~\all_features[1502]  | (~\all_features[1501]  & (new_n15091_ | ~new_n15100_ | ~\all_features[1500] )));
  assign new_n15103_ = new_n15092_ & (~\all_features[1499]  | ~new_n15098_ | (~new_n15099_ & ~\all_features[1498] ));
  assign new_n15104_ = new_n15092_ & (~\all_features[1501]  | (~\all_features[1500]  & (~\all_features[1499]  | (~\all_features[1498]  & ~\all_features[1497] ))));
  assign new_n15105_ = ~new_n15030_ & ((~new_n15031_ & ~new_n15106_ & ~new_n14210_ & new_n15033_) | (new_n15036_ & ~new_n15033_));
  assign new_n15106_ = new_n14207_ & new_n15107_ & new_n14182_;
  assign new_n15107_ = ~new_n15108_ & (\all_features[1507]  | \all_features[1508]  | \all_features[1509]  | \all_features[1510]  | \all_features[1511] );
  assign new_n15108_ = ~new_n14199_ & (new_n14202_ | (~new_n14203_ & (new_n14204_ | (~new_n15109_ & ~new_n14205_))));
  assign new_n15109_ = ~new_n14192_ & (new_n14194_ | (new_n14197_ & (~new_n14196_ | (~new_n15110_ & new_n14185_))));
  assign new_n15110_ = ~\all_features[1509]  & \all_features[1510]  & \all_features[1511]  & (\all_features[1508]  ? new_n14189_ : (new_n14188_ | ~new_n14189_));
  assign new_n15111_ = new_n15112_ & (new_n15041_ | ~new_n15029_) & (~new_n15084_ | new_n15086_);
  assign new_n15112_ = (~new_n15047_ | ~new_n15035_) & (~new_n15085_ | (new_n15088_ ? new_n15087_ : new_n15113_));
  assign new_n15113_ = new_n15114_ & new_n15143_;
  assign new_n15114_ = ~new_n15115_ & ~new_n15139_;
  assign new_n15115_ = new_n15130_ & (~new_n15135_ | (~new_n15133_ & ~new_n15116_ & ~new_n15138_));
  assign new_n15116_ = ~new_n15128_ & ~new_n15126_ & (~new_n15129_ | ~new_n15125_ | new_n15117_);
  assign new_n15117_ = new_n15118_ & new_n15120_ & (new_n15123_ | ~\all_features[1861]  | ~\all_features[1862]  | ~\all_features[1863] );
  assign new_n15118_ = \all_features[1863]  & (\all_features[1862]  | (new_n15119_ & (\all_features[1858]  | \all_features[1859]  | \all_features[1857] )));
  assign new_n15119_ = \all_features[1860]  & \all_features[1861] ;
  assign new_n15120_ = \all_features[1862]  & \all_features[1863]  & (\all_features[1860]  | \all_features[1861]  | new_n15122_ | ~new_n15121_);
  assign new_n15121_ = ~\all_features[1858]  & ~\all_features[1859] ;
  assign new_n15122_ = \all_features[1856]  & \all_features[1857] ;
  assign new_n15123_ = ~\all_features[1859]  & ~\all_features[1860]  & (~\all_features[1858]  | new_n15124_);
  assign new_n15124_ = ~\all_features[1856]  & ~\all_features[1857] ;
  assign new_n15125_ = \all_features[1863]  & (\all_features[1862]  | (\all_features[1861]  & (\all_features[1860]  | ~new_n15121_ | ~new_n15124_)));
  assign new_n15126_ = ~new_n15127_ & ~\all_features[1863] ;
  assign new_n15127_ = \all_features[1861]  & \all_features[1862]  & (\all_features[1860]  | (\all_features[1858]  & \all_features[1859]  & \all_features[1857] ));
  assign new_n15128_ = ~\all_features[1863]  & (~new_n15122_ | ~\all_features[1858]  | ~\all_features[1859]  | ~\all_features[1862]  | ~new_n15119_);
  assign new_n15129_ = \all_features[1863]  & (\all_features[1861]  | \all_features[1862]  | \all_features[1860] );
  assign new_n15130_ = ~new_n15131_ & (\all_features[1859]  | \all_features[1860]  | \all_features[1861]  | \all_features[1862]  | \all_features[1863] );
  assign new_n15131_ = ~\all_features[1861]  & new_n15132_ & ((~\all_features[1858]  & new_n15124_) | ~\all_features[1860]  | ~\all_features[1859] );
  assign new_n15132_ = ~\all_features[1862]  & ~\all_features[1863] ;
  assign new_n15133_ = ~\all_features[1863]  & (~\all_features[1862]  | new_n15134_);
  assign new_n15134_ = ~\all_features[1861]  & (new_n15124_ | ~\all_features[1859]  | ~\all_features[1860]  | ~\all_features[1858] );
  assign new_n15135_ = ~new_n15136_ & ~new_n15137_;
  assign new_n15136_ = new_n15132_ & (~\all_features[1861]  | (~\all_features[1860]  & (~\all_features[1859]  | (~\all_features[1858]  & ~\all_features[1857] ))));
  assign new_n15137_ = new_n15132_ & (~\all_features[1859]  | ~new_n15119_ | (~new_n15122_ & ~\all_features[1858] ));
  assign new_n15138_ = ~\all_features[1863]  & (~\all_features[1862]  | (~\all_features[1861]  & ~\all_features[1860]  & (~\all_features[1859]  | ~\all_features[1858] )));
  assign new_n15139_ = ~new_n15140_ & (\all_features[1859]  | \all_features[1860]  | \all_features[1861]  | \all_features[1862]  | \all_features[1863] );
  assign new_n15140_ = ~new_n15131_ & (new_n15136_ | (~new_n15137_ & (new_n15138_ | (~new_n15133_ & ~new_n15141_))));
  assign new_n15141_ = ~new_n15126_ & (new_n15128_ | (new_n15129_ & (~new_n15125_ | (~new_n15142_ & new_n15118_))));
  assign new_n15142_ = ~\all_features[1861]  & \all_features[1862]  & \all_features[1863]  & (\all_features[1860]  ? new_n15121_ : (new_n15122_ | ~new_n15121_));
  assign new_n15143_ = ~new_n15144_ & ~new_n15147_;
  assign new_n15144_ = new_n15135_ & ~new_n15145_ & new_n15130_;
  assign new_n15145_ = ~new_n15138_ & ~new_n15128_ & ~new_n15126_ & ~new_n15133_ & ~new_n15146_;
  assign new_n15146_ = new_n15129_ & new_n15125_ & new_n15118_ & new_n15120_;
  assign new_n15147_ = new_n15130_ & new_n15148_ & ~new_n15126_ & ~new_n15136_;
  assign new_n15148_ = ~new_n15138_ & ~new_n15137_ & ~new_n15133_ & ~new_n15128_;
  assign new_n15149_ = ~new_n15150_ & new_n15209_;
  assign new_n15150_ = new_n15161_ & (~new_n15151_ | (~new_n15208_ & new_n15206_) | (~new_n15207_ & ~new_n15206_));
  assign new_n15151_ = ~new_n15152_ & new_n13202_;
  assign new_n15152_ = new_n11445_ & ~new_n15153_ & ~new_n15157_;
  assign new_n15153_ = ~new_n15154_ & ~new_n11467_;
  assign new_n15154_ = ~new_n11465_ & (new_n11463_ | (~new_n11466_ & (new_n11454_ | (~new_n11449_ & ~new_n15155_))));
  assign new_n15155_ = ~new_n11452_ & (new_n11455_ | (new_n11462_ & (~new_n11458_ | (~new_n15156_ & new_n11460_))));
  assign new_n15156_ = ~\all_features[5037]  & \all_features[5038]  & \all_features[5039]  & (\all_features[5036]  ? new_n11459_ : (new_n11457_ | ~new_n11459_));
  assign new_n15157_ = ~new_n11465_ & ~new_n11467_ & (~new_n11470_ | (~new_n15158_ & ~new_n11449_ & ~new_n11454_));
  assign new_n15158_ = ~new_n11455_ & ~new_n11452_ & (~new_n11462_ | ~new_n11458_ | new_n15159_);
  assign new_n15159_ = new_n11460_ & new_n11461_ & (new_n15160_ | ~\all_features[5037]  | ~\all_features[5038]  | ~\all_features[5039] );
  assign new_n15160_ = ~\all_features[5035]  & ~\all_features[5036]  & (~\all_features[5034]  | new_n11450_);
  assign new_n15161_ = (new_n15162_ | new_n13202_) & (~new_n15152_ | ~new_n13202_ | (new_n15167_ ? new_n15170_ : ~new_n15165_));
  assign new_n15162_ = ~new_n14046_ & (new_n15164_ | ~new_n15163_);
  assign new_n15163_ = ~new_n14047_ & new_n14070_;
  assign new_n15164_ = ~new_n14073_ & ~new_n14077_;
  assign new_n15165_ = new_n6734_ & (new_n6732_ | new_n15166_);
  assign new_n15166_ = new_n6703_ & new_n6723_;
  assign new_n15167_ = new_n15168_ & new_n15169_;
  assign new_n15168_ = ~new_n12077_ & ~new_n12050_;
  assign new_n15169_ = ~new_n12081_ & ~new_n12074_;
  assign new_n15170_ = new_n15171_ & new_n15197_;
  assign new_n15171_ = new_n15172_ & new_n15195_;
  assign new_n15172_ = new_n15190_ & ~new_n15194_ & ~new_n15173_ & ~new_n15193_;
  assign new_n15173_ = ~new_n15188_ & ~new_n15189_ & new_n15181_ & (~new_n15186_ | ~new_n15174_);
  assign new_n15174_ = new_n15180_ & new_n15175_ & new_n15177_;
  assign new_n15175_ = \all_features[4647]  & (\all_features[4646]  | (new_n15176_ & (\all_features[4642]  | \all_features[4643]  | \all_features[4641] )));
  assign new_n15176_ = \all_features[4644]  & \all_features[4645] ;
  assign new_n15177_ = \all_features[4646]  & \all_features[4647]  & (\all_features[4644]  | \all_features[4645]  | new_n15179_ | ~new_n15178_);
  assign new_n15178_ = ~\all_features[4642]  & ~\all_features[4643] ;
  assign new_n15179_ = \all_features[4640]  & \all_features[4641] ;
  assign new_n15180_ = \all_features[4647]  & (\all_features[4645]  | \all_features[4646]  | \all_features[4644] );
  assign new_n15181_ = ~new_n15182_ & ~new_n15184_;
  assign new_n15182_ = ~new_n15183_ & ~\all_features[4647] ;
  assign new_n15183_ = \all_features[4645]  & \all_features[4646]  & (\all_features[4644]  | (\all_features[4642]  & \all_features[4643]  & \all_features[4641] ));
  assign new_n15184_ = ~\all_features[4647]  & (~\all_features[4646]  | (~\all_features[4644]  & ~\all_features[4645]  & ~new_n15185_));
  assign new_n15185_ = \all_features[4642]  & \all_features[4643] ;
  assign new_n15186_ = \all_features[4647]  & (\all_features[4646]  | (\all_features[4645]  & (\all_features[4644]  | ~new_n15187_ | ~new_n15178_)));
  assign new_n15187_ = ~\all_features[4640]  & ~\all_features[4641] ;
  assign new_n15188_ = ~\all_features[4647]  & (~\all_features[4646]  | (~\all_features[4645]  & (new_n15187_ | ~new_n15185_ | ~\all_features[4644] )));
  assign new_n15189_ = ~\all_features[4647]  & (~\all_features[4646]  | ~new_n15176_ | ~new_n15179_ | ~new_n15185_);
  assign new_n15190_ = ~new_n15191_ & (\all_features[4643]  | \all_features[4644]  | \all_features[4645]  | \all_features[4646]  | \all_features[4647] );
  assign new_n15191_ = ~\all_features[4645]  & new_n15192_ & ((~\all_features[4642]  & new_n15187_) | ~\all_features[4644]  | ~\all_features[4643] );
  assign new_n15192_ = ~\all_features[4646]  & ~\all_features[4647] ;
  assign new_n15193_ = new_n15192_ & (~\all_features[4645]  | (~\all_features[4644]  & (~\all_features[4643]  | (~\all_features[4642]  & ~\all_features[4641] ))));
  assign new_n15194_ = new_n15192_ & (~\all_features[4643]  | ~new_n15176_ | (~\all_features[4642]  & ~new_n15179_));
  assign new_n15195_ = new_n15190_ & new_n15181_ & new_n15196_ & ~new_n15188_ & ~new_n15189_;
  assign new_n15196_ = ~new_n15193_ & ~new_n15194_;
  assign new_n15197_ = new_n15198_ & new_n15202_;
  assign new_n15198_ = new_n15190_ & (~new_n15196_ | (~new_n15199_ & ~new_n15184_ & ~new_n15188_));
  assign new_n15199_ = ~new_n15189_ & ~new_n15182_ & (~new_n15180_ | ~new_n15186_ | new_n15200_);
  assign new_n15200_ = new_n15175_ & new_n15177_ & (new_n15201_ | ~\all_features[4645]  | ~\all_features[4646]  | ~\all_features[4647] );
  assign new_n15201_ = ~\all_features[4643]  & ~\all_features[4644]  & (~\all_features[4642]  | new_n15187_);
  assign new_n15202_ = ~new_n15203_ & (\all_features[4643]  | \all_features[4644]  | \all_features[4645]  | \all_features[4646]  | \all_features[4647] );
  assign new_n15203_ = ~new_n15191_ & (new_n15193_ | (~new_n15194_ & (new_n15184_ | (~new_n15188_ & ~new_n15204_))));
  assign new_n15204_ = ~new_n15182_ & (new_n15189_ | (new_n15180_ & (~new_n15186_ | (~new_n15205_ & new_n15175_))));
  assign new_n15205_ = ~\all_features[4645]  & \all_features[4646]  & \all_features[4647]  & (\all_features[4644]  ? new_n15178_ : (new_n15179_ | ~new_n15178_));
  assign new_n15206_ = new_n12721_ & (new_n12718_ | ~new_n12687_);
  assign new_n15207_ = ~new_n11236_ & (~new_n11233_ | ~new_n14291_);
  assign new_n15208_ = ~new_n8388_ & (~new_n8357_ | ~new_n8385_);
  assign new_n15209_ = new_n15210_ & (~new_n15151_ | (new_n15208_ & new_n15206_) | (new_n15207_ & ~new_n15206_));
  assign new_n15210_ = (~new_n15162_ | new_n13202_) & (new_n15165_ | new_n15167_ | ~new_n15152_ | ~new_n13202_);
  assign new_n15211_ = ~new_n15212_ & new_n15349_;
  assign new_n15212_ = (new_n15320_ & new_n15329_ & new_n15332_) | (~new_n15332_ & (new_n15331_ ? new_n15213_ : new_n15281_));
  assign new_n15213_ = (new_n15214_ & new_n15264_) ? new_n15247_ : new_n15265_;
  assign new_n15214_ = new_n15215_ & new_n15244_;
  assign new_n15215_ = new_n15216_ & new_n15237_;
  assign new_n15216_ = ~new_n15217_ & (\all_features[1707]  | \all_features[1708]  | \all_features[1709]  | \all_features[1710]  | \all_features[1711] );
  assign new_n15217_ = ~new_n15233_ & (new_n15231_ | (~new_n15235_ & (new_n15236_ | (~new_n15234_ & ~new_n15218_))));
  assign new_n15218_ = ~new_n15219_ & (new_n15221_ | (new_n15230_ & (~new_n15225_ | (~new_n15229_ & new_n15228_))));
  assign new_n15219_ = ~new_n15220_ & ~\all_features[1711] ;
  assign new_n15220_ = \all_features[1709]  & \all_features[1710]  & (\all_features[1708]  | (\all_features[1706]  & \all_features[1707]  & \all_features[1705] ));
  assign new_n15221_ = ~\all_features[1711]  & (~\all_features[1710]  | ~new_n15222_ | ~new_n15223_ | ~new_n15224_);
  assign new_n15222_ = \all_features[1706]  & \all_features[1707] ;
  assign new_n15223_ = \all_features[1704]  & \all_features[1705] ;
  assign new_n15224_ = \all_features[1708]  & \all_features[1709] ;
  assign new_n15225_ = \all_features[1711]  & (\all_features[1710]  | (\all_features[1709]  & (\all_features[1708]  | ~new_n15227_ | ~new_n15226_)));
  assign new_n15226_ = ~\all_features[1704]  & ~\all_features[1705] ;
  assign new_n15227_ = ~\all_features[1706]  & ~\all_features[1707] ;
  assign new_n15228_ = \all_features[1711]  & (\all_features[1710]  | (new_n15224_ & (\all_features[1706]  | \all_features[1707]  | \all_features[1705] )));
  assign new_n15229_ = ~\all_features[1709]  & \all_features[1710]  & \all_features[1711]  & (\all_features[1708]  ? new_n15227_ : (new_n15223_ | ~new_n15227_));
  assign new_n15230_ = \all_features[1711]  & (\all_features[1709]  | \all_features[1710]  | \all_features[1708] );
  assign new_n15231_ = new_n15232_ & (~\all_features[1709]  | (~\all_features[1708]  & (~\all_features[1707]  | (~\all_features[1706]  & ~\all_features[1705] ))));
  assign new_n15232_ = ~\all_features[1710]  & ~\all_features[1711] ;
  assign new_n15233_ = ~\all_features[1709]  & new_n15232_ & ((~\all_features[1706]  & new_n15226_) | ~\all_features[1708]  | ~\all_features[1707] );
  assign new_n15234_ = ~\all_features[1711]  & (~\all_features[1710]  | (~\all_features[1709]  & (new_n15226_ | ~new_n15222_ | ~\all_features[1708] )));
  assign new_n15235_ = new_n15232_ & (~\all_features[1707]  | ~new_n15224_ | (~\all_features[1706]  & ~new_n15223_));
  assign new_n15236_ = ~\all_features[1711]  & (~\all_features[1710]  | (~\all_features[1708]  & ~\all_features[1709]  & ~new_n15222_));
  assign new_n15237_ = new_n15242_ & (~new_n15243_ | (~new_n15238_ & ~new_n15234_ & ~new_n15236_));
  assign new_n15238_ = ~new_n15219_ & ~new_n15221_ & (~new_n15230_ | ~new_n15225_ | new_n15239_);
  assign new_n15239_ = new_n15228_ & new_n15240_ & (new_n15241_ | ~\all_features[1709]  | ~\all_features[1710]  | ~\all_features[1711] );
  assign new_n15240_ = \all_features[1710]  & \all_features[1711]  & (\all_features[1708]  | \all_features[1709]  | new_n15223_ | ~new_n15227_);
  assign new_n15241_ = ~\all_features[1707]  & ~\all_features[1708]  & (~\all_features[1706]  | new_n15226_);
  assign new_n15242_ = ~new_n15233_ & (\all_features[1707]  | \all_features[1708]  | \all_features[1709]  | \all_features[1710]  | \all_features[1711] );
  assign new_n15243_ = ~new_n15231_ & ~new_n15235_;
  assign new_n15244_ = new_n15242_ & new_n15243_ & (new_n15246_ | new_n15219_ | new_n15234_ | ~new_n15245_);
  assign new_n15245_ = ~new_n15221_ & ~new_n15236_;
  assign new_n15246_ = new_n15230_ & new_n15240_ & new_n15225_ & new_n15228_;
  assign new_n15247_ = new_n15259_ & new_n15251_ & ~new_n15263_ & ~new_n15262_ & ~new_n15248_ & ~new_n15257_;
  assign new_n15248_ = ~\all_features[1231]  & (~\all_features[1230]  | new_n15249_);
  assign new_n15249_ = ~\all_features[1229]  & (new_n15250_ | ~\all_features[1227]  | ~\all_features[1228]  | ~\all_features[1226] );
  assign new_n15250_ = ~\all_features[1224]  & ~\all_features[1225] ;
  assign new_n15251_ = ~new_n15252_ & ~new_n15256_;
  assign new_n15252_ = new_n15253_ & (~\all_features[1227]  | ~new_n15255_ | (~\all_features[1226]  & ~new_n15254_));
  assign new_n15253_ = ~\all_features[1230]  & ~\all_features[1231] ;
  assign new_n15254_ = \all_features[1224]  & \all_features[1225] ;
  assign new_n15255_ = \all_features[1228]  & \all_features[1229] ;
  assign new_n15256_ = new_n15253_ & (~\all_features[1229]  | (~\all_features[1228]  & (~\all_features[1227]  | (~\all_features[1226]  & ~\all_features[1225] ))));
  assign new_n15257_ = ~new_n15258_ & ~\all_features[1231] ;
  assign new_n15258_ = \all_features[1229]  & \all_features[1230]  & (\all_features[1228]  | (\all_features[1226]  & \all_features[1227]  & \all_features[1225] ));
  assign new_n15259_ = ~new_n15260_ & ~new_n15261_;
  assign new_n15260_ = ~\all_features[1231]  & ~\all_features[1230]  & ~\all_features[1229]  & ~\all_features[1227]  & ~\all_features[1228] ;
  assign new_n15261_ = ~\all_features[1231]  & (~\all_features[1230]  | (~\all_features[1229]  & ~\all_features[1228]  & (~\all_features[1227]  | ~\all_features[1226] )));
  assign new_n15262_ = ~\all_features[1229]  & new_n15253_ & ((~\all_features[1226]  & new_n15250_) | ~\all_features[1228]  | ~\all_features[1227] );
  assign new_n15263_ = ~\all_features[1231]  & (~new_n15255_ | ~\all_features[1226]  | ~\all_features[1227]  | ~\all_features[1230]  | ~new_n15254_);
  assign new_n15264_ = new_n15245_ & new_n15242_ & ~new_n15235_ & ~new_n15234_ & ~new_n15219_ & ~new_n15231_;
  assign new_n15265_ = new_n15271_ & new_n15266_ & ~new_n15280_ & ~new_n15279_ & ~new_n15275_ & ~new_n15277_;
  assign new_n15266_ = ~new_n15267_ & ~new_n15269_;
  assign new_n15267_ = new_n15268_ & ~\all_features[1045]  & ~\all_features[1043]  & ~\all_features[1044] ;
  assign new_n15268_ = ~\all_features[1046]  & ~\all_features[1047] ;
  assign new_n15269_ = ~\all_features[1047]  & (~\all_features[1046]  | (~\all_features[1044]  & ~\all_features[1045]  & ~new_n15270_));
  assign new_n15270_ = \all_features[1042]  & \all_features[1043] ;
  assign new_n15271_ = ~new_n15272_ & ~new_n15274_;
  assign new_n15272_ = new_n15268_ & (~new_n15273_ | ~\all_features[1043]  | (~\all_features[1042]  & (~\all_features[1040]  | ~\all_features[1041] )));
  assign new_n15273_ = \all_features[1044]  & \all_features[1045] ;
  assign new_n15274_ = new_n15268_ & (~\all_features[1045]  | (~\all_features[1044]  & (~\all_features[1043]  | (~\all_features[1042]  & ~\all_features[1041] ))));
  assign new_n15275_ = ~new_n15276_ & ~\all_features[1047] ;
  assign new_n15276_ = \all_features[1045]  & \all_features[1046]  & (\all_features[1044]  | (\all_features[1042]  & \all_features[1043]  & \all_features[1041] ));
  assign new_n15277_ = ~\all_features[1045]  & new_n15268_ & ((~\all_features[1042]  & new_n15278_) | ~\all_features[1044]  | ~\all_features[1043] );
  assign new_n15278_ = ~\all_features[1040]  & ~\all_features[1041] ;
  assign new_n15279_ = ~\all_features[1047]  & (~new_n15273_ | ~\all_features[1040]  | ~\all_features[1041]  | ~\all_features[1046]  | ~new_n15270_);
  assign new_n15280_ = ~\all_features[1047]  & (~\all_features[1046]  | (~\all_features[1045]  & (new_n15278_ | ~\all_features[1044]  | ~new_n15270_)));
  assign new_n15281_ = ~new_n15282_ & ~new_n15318_;
  assign new_n15282_ = new_n15283_ & new_n15311_;
  assign new_n15283_ = ~new_n15284_ & ~new_n15308_;
  assign new_n15284_ = ~new_n15307_ & ~new_n15306_ & ~new_n15305_ & ~new_n15285_ & ~new_n15303_;
  assign new_n15285_ = new_n15289_ & new_n15293_ & (~new_n15300_ | ~new_n15302_ | ~new_n15286_ | ~new_n15299_);
  assign new_n15286_ = \all_features[1471]  & (\all_features[1470]  | new_n15287_);
  assign new_n15287_ = \all_features[1469]  & (\all_features[1466]  | \all_features[1467]  | \all_features[1468]  | ~new_n15288_);
  assign new_n15288_ = ~\all_features[1464]  & ~\all_features[1465] ;
  assign new_n15289_ = ~new_n15290_ & ~new_n15292_;
  assign new_n15290_ = ~\all_features[1471]  & (~\all_features[1470]  | (~\all_features[1468]  & ~\all_features[1469]  & ~new_n15291_));
  assign new_n15291_ = \all_features[1466]  & \all_features[1467] ;
  assign new_n15292_ = ~\all_features[1471]  & (~\all_features[1470]  | (~\all_features[1469]  & (new_n15288_ | ~new_n15291_ | ~\all_features[1468] )));
  assign new_n15293_ = ~new_n15294_ & ~new_n15297_;
  assign new_n15294_ = ~\all_features[1471]  & (~\all_features[1470]  | ~new_n15295_ | ~new_n15296_ | ~new_n15291_);
  assign new_n15295_ = \all_features[1468]  & \all_features[1469] ;
  assign new_n15296_ = \all_features[1464]  & \all_features[1465] ;
  assign new_n15297_ = ~new_n15298_ & ~\all_features[1471] ;
  assign new_n15298_ = \all_features[1469]  & \all_features[1470]  & (\all_features[1468]  | (\all_features[1466]  & \all_features[1467]  & \all_features[1465] ));
  assign new_n15299_ = \all_features[1471]  & (\all_features[1470]  | (new_n15295_ & (\all_features[1466]  | \all_features[1467]  | \all_features[1465] )));
  assign new_n15300_ = new_n15301_ & (new_n15296_ | \all_features[1466]  | \all_features[1467]  | \all_features[1468]  | \all_features[1469] );
  assign new_n15301_ = \all_features[1470]  & \all_features[1471] ;
  assign new_n15302_ = \all_features[1471]  & (\all_features[1469]  | \all_features[1470]  | \all_features[1468] );
  assign new_n15303_ = new_n15304_ & (~\all_features[1469]  | (~\all_features[1468]  & (~\all_features[1467]  | (~\all_features[1466]  & ~\all_features[1465] ))));
  assign new_n15304_ = ~\all_features[1470]  & ~\all_features[1471] ;
  assign new_n15305_ = ~\all_features[1469]  & new_n15304_ & ((~\all_features[1466]  & new_n15288_) | ~\all_features[1468]  | ~\all_features[1467] );
  assign new_n15306_ = new_n15304_ & (~\all_features[1467]  | ~new_n15295_ | (~\all_features[1466]  & ~new_n15296_));
  assign new_n15307_ = ~\all_features[1471]  & ~\all_features[1470]  & ~\all_features[1469]  & ~\all_features[1467]  & ~\all_features[1468] ;
  assign new_n15308_ = new_n15310_ & new_n15309_ & ~new_n15305_ & ~new_n15297_ & ~new_n15290_ & ~new_n15292_;
  assign new_n15309_ = ~new_n15294_ & ~new_n15307_;
  assign new_n15310_ = ~new_n15303_ & ~new_n15306_;
  assign new_n15311_ = ~new_n15315_ & (new_n15307_ | (~new_n15305_ & ~new_n15312_));
  assign new_n15312_ = ~new_n15303_ & (new_n15306_ | (~new_n15290_ & (new_n15292_ | (~new_n15297_ & ~new_n15313_))));
  assign new_n15313_ = ~new_n15294_ & (~new_n15302_ | (new_n15286_ & (~new_n15299_ | (~new_n15314_ & new_n15300_))));
  assign new_n15314_ = new_n15301_ & (\all_features[1469]  | (\all_features[1468]  & (\all_features[1467]  | \all_features[1466] )));
  assign new_n15315_ = ~new_n15305_ & ~new_n15307_ & (~new_n15310_ | (~new_n15316_ & new_n15289_));
  assign new_n15316_ = new_n15293_ & ((~new_n15317_ & new_n15300_ & new_n15299_) | ~new_n15302_ | ~new_n15286_);
  assign new_n15317_ = new_n15301_ & \all_features[1469]  & ((~new_n15288_ & \all_features[1466] ) | \all_features[1468]  | \all_features[1467] );
  assign new_n15318_ = new_n8482_ & new_n15319_;
  assign new_n15319_ = new_n7899_ & new_n7902_;
  assign new_n15320_ = new_n15321_ & new_n15328_;
  assign new_n15321_ = ~new_n15322_ & ~new_n10972_;
  assign new_n15322_ = (new_n15323_ | (new_n10965_ & (~\all_features[1899]  | ~\all_features[1900]  | (~\all_features[1898]  & new_n10953_)))) & (~new_n10965_ | \all_features[1899]  | \all_features[1900] );
  assign new_n15323_ = ~new_n10969_ & (new_n10968_ | (~new_n10963_ & ~new_n15324_));
  assign new_n15324_ = ~new_n10958_ & (new_n10960_ | (~new_n10962_ & (~new_n15327_ | new_n15325_)));
  assign new_n15325_ = \all_features[1903]  & ((~new_n15326_ & ~\all_features[1901]  & \all_features[1902] ) | (~new_n10955_ & (\all_features[1902]  | (~new_n10952_ & \all_features[1901] ))));
  assign new_n15326_ = (~\all_features[1898]  & ~\all_features[1899]  & ~\all_features[1900]  & (~\all_features[1897]  | ~\all_features[1896] )) | (\all_features[1900]  & (\all_features[1898]  | \all_features[1899] ));
  assign new_n15327_ = \all_features[1903]  & (\all_features[1901]  | \all_features[1902]  | \all_features[1900] );
  assign new_n15328_ = ~new_n10949_ & ~new_n10970_;
  assign new_n15329_ = new_n12409_ & new_n15330_;
  assign new_n15330_ = ~new_n12439_ & ~new_n12442_;
  assign new_n15331_ = ~new_n12595_ & (~new_n12588_ | ~new_n12592_ | ~new_n12564_);
  assign new_n15332_ = new_n15344_ & new_n15336_ & ~new_n15348_ & ~new_n15347_ & ~new_n15333_ & ~new_n15342_;
  assign new_n15333_ = ~\all_features[5679]  & (~\all_features[5678]  | new_n15334_);
  assign new_n15334_ = ~\all_features[5677]  & (new_n15335_ | ~\all_features[5675]  | ~\all_features[5676]  | ~\all_features[5674] );
  assign new_n15335_ = ~\all_features[5672]  & ~\all_features[5673] ;
  assign new_n15336_ = ~new_n15337_ & ~new_n15341_;
  assign new_n15337_ = new_n15338_ & (~\all_features[5675]  | ~new_n15340_ | (~\all_features[5674]  & ~new_n15339_));
  assign new_n15338_ = ~\all_features[5678]  & ~\all_features[5679] ;
  assign new_n15339_ = \all_features[5672]  & \all_features[5673] ;
  assign new_n15340_ = \all_features[5676]  & \all_features[5677] ;
  assign new_n15341_ = new_n15338_ & (~\all_features[5677]  | (~\all_features[5676]  & (~\all_features[5675]  | (~\all_features[5674]  & ~\all_features[5673] ))));
  assign new_n15342_ = ~new_n15343_ & ~\all_features[5679] ;
  assign new_n15343_ = \all_features[5677]  & \all_features[5678]  & (\all_features[5676]  | (\all_features[5674]  & \all_features[5675]  & \all_features[5673] ));
  assign new_n15344_ = ~new_n15345_ & ~new_n15346_;
  assign new_n15345_ = ~\all_features[5679]  & ~\all_features[5678]  & ~\all_features[5677]  & ~\all_features[5675]  & ~\all_features[5676] ;
  assign new_n15346_ = ~\all_features[5679]  & (~\all_features[5678]  | (~\all_features[5677]  & ~\all_features[5676]  & (~\all_features[5675]  | ~\all_features[5674] )));
  assign new_n15347_ = ~\all_features[5677]  & new_n15338_ & ((~\all_features[5674]  & new_n15335_) | ~\all_features[5676]  | ~\all_features[5675] );
  assign new_n15348_ = ~\all_features[5679]  & (~new_n15340_ | ~\all_features[5674]  | ~\all_features[5675]  | ~\all_features[5678]  | ~new_n15339_);
  assign new_n15349_ = new_n15332_ | (new_n15331_ ? ~new_n15213_ : ~new_n15281_);
  assign new_n15350_ = (~new_n15364_ | new_n13202_) & (new_n15351_ | ~new_n15365_ | ~new_n13202_);
  assign new_n15351_ = ~new_n7957_ & (new_n15088_ | (new_n15352_ & new_n15362_));
  assign new_n15352_ = new_n15089_ & (new_n15103_ | new_n15104_ | (new_n15361_ & (new_n15353_ | ~new_n15094_)));
  assign new_n15353_ = new_n15354_ & (~new_n15357_ | (~new_n15360_ & \all_features[1501]  & \all_features[1502]  & \all_features[1503] ));
  assign new_n15354_ = \all_features[1503]  & (\all_features[1502]  | (~new_n15355_ & \all_features[1501] ));
  assign new_n15355_ = new_n15091_ & ~\all_features[1500]  & new_n15356_;
  assign new_n15356_ = ~\all_features[1498]  & ~\all_features[1499] ;
  assign new_n15357_ = \all_features[1503]  & \all_features[1502]  & ~new_n15359_ & new_n15358_;
  assign new_n15358_ = \all_features[1503]  & (\all_features[1502]  | (new_n15098_ & (\all_features[1498]  | \all_features[1499]  | \all_features[1497] )));
  assign new_n15359_ = new_n15356_ & ~\all_features[1501]  & ~new_n15099_ & ~\all_features[1500] ;
  assign new_n15360_ = ~\all_features[1499]  & ~\all_features[1500]  & (~\all_features[1498]  | new_n15091_);
  assign new_n15361_ = ~new_n15101_ & ~new_n15102_;
  assign new_n15362_ = new_n15089_ & ~new_n15104_ & ~new_n15363_ & ~new_n15103_;
  assign new_n15363_ = ~new_n15095_ & ~new_n15097_ & ~new_n15101_ & ~new_n15102_ & (~new_n15357_ | ~new_n15354_);
  assign new_n15364_ = new_n12197_ & new_n12226_;
  assign new_n15365_ = ~new_n15399_ & (~new_n15396_ | new_n15366_);
  assign new_n15366_ = ~new_n15367_ & (new_n15386_ | (~new_n15392_ & ~new_n15384_));
  assign new_n15367_ = new_n15383_ & (~new_n15387_ | (~new_n15368_ & ~new_n15390_ & ~new_n15391_));
  assign new_n15368_ = ~new_n15380_ & ~new_n15378_ & (~new_n15382_ | new_n15372_ | ~new_n15369_);
  assign new_n15369_ = \all_features[5695]  & (\all_features[5694]  | new_n15370_);
  assign new_n15370_ = \all_features[5693]  & (\all_features[5690]  | \all_features[5691]  | \all_features[5692]  | ~new_n15371_);
  assign new_n15371_ = ~\all_features[5688]  & ~\all_features[5689] ;
  assign new_n15372_ = ~new_n15375_ & new_n15373_ & \all_features[5694]  & \all_features[5695]  & (~\all_features[5693]  | new_n15377_);
  assign new_n15373_ = \all_features[5695]  & (\all_features[5694]  | (new_n15374_ & (\all_features[5690]  | \all_features[5691]  | \all_features[5689] )));
  assign new_n15374_ = \all_features[5692]  & \all_features[5693] ;
  assign new_n15375_ = ~\all_features[5693]  & ~\all_features[5692]  & ~\all_features[5691]  & ~new_n15376_ & ~\all_features[5690] ;
  assign new_n15376_ = \all_features[5688]  & \all_features[5689] ;
  assign new_n15377_ = ~\all_features[5691]  & ~\all_features[5692]  & (~\all_features[5690]  | new_n15371_);
  assign new_n15378_ = ~new_n15379_ & ~\all_features[5695] ;
  assign new_n15379_ = \all_features[5693]  & \all_features[5694]  & (\all_features[5692]  | (\all_features[5690]  & \all_features[5691]  & \all_features[5689] ));
  assign new_n15380_ = ~\all_features[5695]  & (~\all_features[5694]  | ~new_n15381_ | ~new_n15376_ | ~new_n15374_);
  assign new_n15381_ = \all_features[5690]  & \all_features[5691] ;
  assign new_n15382_ = \all_features[5695]  & (\all_features[5693]  | \all_features[5694]  | \all_features[5692] );
  assign new_n15383_ = ~new_n15384_ & ~new_n15386_;
  assign new_n15384_ = ~\all_features[5693]  & new_n15385_ & ((~\all_features[5690]  & new_n15371_) | ~\all_features[5692]  | ~\all_features[5691] );
  assign new_n15385_ = ~\all_features[5694]  & ~\all_features[5695] ;
  assign new_n15386_ = ~\all_features[5695]  & ~\all_features[5694]  & ~\all_features[5693]  & ~\all_features[5691]  & ~\all_features[5692] ;
  assign new_n15387_ = ~new_n15388_ & ~new_n15389_;
  assign new_n15388_ = new_n15385_ & (~\all_features[5693]  | (~\all_features[5692]  & (~\all_features[5691]  | (~\all_features[5690]  & ~\all_features[5689] ))));
  assign new_n15389_ = new_n15385_ & (~\all_features[5691]  | ~new_n15374_ | (~\all_features[5690]  & ~new_n15376_));
  assign new_n15390_ = ~\all_features[5695]  & (~\all_features[5694]  | (~\all_features[5693]  & (new_n15371_ | ~new_n15381_ | ~\all_features[5692] )));
  assign new_n15391_ = ~\all_features[5695]  & (~\all_features[5694]  | (~\all_features[5692]  & ~\all_features[5693]  & ~new_n15381_));
  assign new_n15392_ = ~new_n15388_ & (new_n15389_ | (~new_n15391_ & (new_n15390_ | (~new_n15378_ & ~new_n15393_))));
  assign new_n15393_ = ~new_n15380_ & (~new_n15382_ | (new_n15369_ & (~new_n15373_ | (~new_n15395_ & new_n15394_))));
  assign new_n15394_ = \all_features[5695]  & ~new_n15375_ & \all_features[5694] ;
  assign new_n15395_ = \all_features[5694]  & \all_features[5695]  & (\all_features[5693]  | (\all_features[5692]  & (\all_features[5691]  | \all_features[5690] )));
  assign new_n15396_ = new_n15383_ & new_n15387_ & (new_n15397_ | new_n15378_ | new_n15390_ | ~new_n15398_);
  assign new_n15397_ = new_n15382_ & new_n15373_ & new_n15369_ & new_n15394_;
  assign new_n15398_ = ~new_n15380_ & ~new_n15391_;
  assign new_n15399_ = new_n15398_ & new_n15383_ & ~new_n15389_ & ~new_n15390_ & ~new_n15378_ & ~new_n15388_;
  assign new_n15400_ = new_n15401_ ? (~new_n15908_ ^ new_n16062_) : (new_n15908_ ^ new_n16062_);
  assign new_n15401_ = new_n15402_ ? (new_n15708_ ^ new_n15907_) : (~new_n15708_ ^ new_n15907_);
  assign new_n15402_ = new_n15403_ ? (new_n15544_ ^ new_n15666_) : (~new_n15544_ ^ new_n15666_);
  assign new_n15403_ = ~new_n15404_ & new_n15541_;
  assign new_n15404_ = new_n15405_ & ~new_n15532_ & new_n15482_;
  assign new_n15405_ = (~new_n15481_ | ~new_n15442_) & (~new_n15406_ | (new_n9689_ ? new_n14504_ : ~new_n15479_));
  assign new_n15406_ = ~new_n13405_ & new_n15407_;
  assign new_n15407_ = new_n15441_ & (new_n15437_ | ~new_n15408_);
  assign new_n15408_ = ~new_n15409_ & ~new_n15433_;
  assign new_n15409_ = ~new_n15431_ & ~new_n15430_ & (~new_n15424_ | (~new_n15410_ & ~new_n15428_ & ~new_n15432_));
  assign new_n15410_ = ~new_n15419_ & ~new_n15420_ & (~new_n15423_ | ~new_n15422_ | new_n15411_);
  assign new_n15411_ = new_n15412_ & new_n15414_ & (new_n15417_ | ~\all_features[1253]  | ~\all_features[1254]  | ~\all_features[1255] );
  assign new_n15412_ = \all_features[1255]  & (\all_features[1254]  | (new_n15413_ & (\all_features[1250]  | \all_features[1251]  | \all_features[1249] )));
  assign new_n15413_ = \all_features[1252]  & \all_features[1253] ;
  assign new_n15414_ = \all_features[1254]  & \all_features[1255]  & (\all_features[1252]  | \all_features[1253]  | new_n15415_ | ~new_n15416_);
  assign new_n15415_ = \all_features[1248]  & \all_features[1249] ;
  assign new_n15416_ = ~\all_features[1250]  & ~\all_features[1251] ;
  assign new_n15417_ = ~\all_features[1251]  & ~\all_features[1252]  & (~\all_features[1250]  | new_n15418_);
  assign new_n15418_ = ~\all_features[1248]  & ~\all_features[1249] ;
  assign new_n15419_ = ~\all_features[1255]  & (~new_n15413_ | ~\all_features[1250]  | ~\all_features[1251]  | ~\all_features[1254]  | ~new_n15415_);
  assign new_n15420_ = ~new_n15421_ & ~\all_features[1255] ;
  assign new_n15421_ = \all_features[1253]  & \all_features[1254]  & (\all_features[1252]  | (\all_features[1250]  & \all_features[1251]  & \all_features[1249] ));
  assign new_n15422_ = \all_features[1255]  & (\all_features[1254]  | (\all_features[1253]  & (\all_features[1252]  | ~new_n15416_ | ~new_n15418_)));
  assign new_n15423_ = \all_features[1255]  & (\all_features[1253]  | \all_features[1254]  | \all_features[1252] );
  assign new_n15424_ = ~new_n15425_ & ~new_n15427_;
  assign new_n15425_ = new_n15426_ & (~\all_features[1251]  | ~new_n15413_ | (~\all_features[1250]  & ~new_n15415_));
  assign new_n15426_ = ~\all_features[1254]  & ~\all_features[1255] ;
  assign new_n15427_ = new_n15426_ & (~\all_features[1253]  | (~\all_features[1252]  & (~\all_features[1251]  | (~\all_features[1250]  & ~\all_features[1249] ))));
  assign new_n15428_ = ~\all_features[1255]  & (~\all_features[1254]  | new_n15429_);
  assign new_n15429_ = ~\all_features[1253]  & (new_n15418_ | ~\all_features[1251]  | ~\all_features[1252]  | ~\all_features[1250] );
  assign new_n15430_ = ~\all_features[1253]  & new_n15426_ & ((~\all_features[1250]  & new_n15418_) | ~\all_features[1252]  | ~\all_features[1251] );
  assign new_n15431_ = ~\all_features[1255]  & ~\all_features[1254]  & ~\all_features[1253]  & ~\all_features[1251]  & ~\all_features[1252] ;
  assign new_n15432_ = ~\all_features[1255]  & (~\all_features[1254]  | (~\all_features[1253]  & ~\all_features[1252]  & (~\all_features[1251]  | ~\all_features[1250] )));
  assign new_n15433_ = ~new_n15434_ & ~new_n15431_;
  assign new_n15434_ = ~new_n15430_ & (new_n15427_ | (~new_n15425_ & (new_n15432_ | (~new_n15428_ & ~new_n15435_))));
  assign new_n15435_ = ~new_n15420_ & (new_n15419_ | (new_n15423_ & (~new_n15422_ | (~new_n15436_ & new_n15412_))));
  assign new_n15436_ = ~\all_features[1253]  & \all_features[1254]  & \all_features[1255]  & (\all_features[1252]  ? new_n15416_ : (new_n15415_ | ~new_n15416_));
  assign new_n15437_ = ~new_n15431_ & ~new_n15430_ & ~new_n15427_ & ~new_n15438_ & ~new_n15425_;
  assign new_n15438_ = ~new_n15428_ & ~new_n15419_ & new_n15439_ & (~new_n15422_ | ~new_n15440_);
  assign new_n15439_ = ~new_n15420_ & ~new_n15432_;
  assign new_n15440_ = new_n15423_ & new_n15412_ & new_n15414_;
  assign new_n15441_ = new_n15424_ & new_n15439_ & ~new_n15431_ & ~new_n15419_ & ~new_n15428_ & ~new_n15430_;
  assign new_n15442_ = new_n15478_ & ~new_n15443_ & new_n13405_;
  assign new_n15443_ = ~new_n15477_ & (~new_n15473_ | ~new_n15444_);
  assign new_n15444_ = new_n15445_ & new_n15469_;
  assign new_n15445_ = ~new_n15467_ & ~new_n15466_ & (~new_n15460_ | (~new_n15446_ & ~new_n15464_ & ~new_n15468_));
  assign new_n15446_ = ~new_n15455_ & ~new_n15456_ & (~new_n15459_ | ~new_n15458_ | new_n15447_);
  assign new_n15447_ = new_n15448_ & new_n15450_ & (new_n15453_ | ~\all_features[3469]  | ~\all_features[3470]  | ~\all_features[3471] );
  assign new_n15448_ = \all_features[3471]  & (\all_features[3470]  | (new_n15449_ & (\all_features[3466]  | \all_features[3467]  | \all_features[3465] )));
  assign new_n15449_ = \all_features[3468]  & \all_features[3469] ;
  assign new_n15450_ = \all_features[3470]  & \all_features[3471]  & (\all_features[3468]  | \all_features[3469]  | new_n15451_ | ~new_n15452_);
  assign new_n15451_ = \all_features[3464]  & \all_features[3465] ;
  assign new_n15452_ = ~\all_features[3466]  & ~\all_features[3467] ;
  assign new_n15453_ = ~\all_features[3467]  & ~\all_features[3468]  & (~\all_features[3466]  | new_n15454_);
  assign new_n15454_ = ~\all_features[3464]  & ~\all_features[3465] ;
  assign new_n15455_ = ~\all_features[3471]  & (~new_n15449_ | ~\all_features[3466]  | ~\all_features[3467]  | ~\all_features[3470]  | ~new_n15451_);
  assign new_n15456_ = ~new_n15457_ & ~\all_features[3471] ;
  assign new_n15457_ = \all_features[3469]  & \all_features[3470]  & (\all_features[3468]  | (\all_features[3466]  & \all_features[3467]  & \all_features[3465] ));
  assign new_n15458_ = \all_features[3471]  & (\all_features[3470]  | (\all_features[3469]  & (\all_features[3468]  | ~new_n15452_ | ~new_n15454_)));
  assign new_n15459_ = \all_features[3471]  & (\all_features[3469]  | \all_features[3470]  | \all_features[3468] );
  assign new_n15460_ = ~new_n15461_ & ~new_n15463_;
  assign new_n15461_ = new_n15462_ & (~\all_features[3467]  | ~new_n15449_ | (~\all_features[3466]  & ~new_n15451_));
  assign new_n15462_ = ~\all_features[3470]  & ~\all_features[3471] ;
  assign new_n15463_ = new_n15462_ & (~\all_features[3469]  | (~\all_features[3468]  & (~\all_features[3467]  | (~\all_features[3466]  & ~\all_features[3465] ))));
  assign new_n15464_ = ~\all_features[3471]  & (~\all_features[3470]  | new_n15465_);
  assign new_n15465_ = ~\all_features[3469]  & (new_n15454_ | ~\all_features[3467]  | ~\all_features[3468]  | ~\all_features[3466] );
  assign new_n15466_ = ~\all_features[3469]  & new_n15462_ & ((~\all_features[3466]  & new_n15454_) | ~\all_features[3468]  | ~\all_features[3467] );
  assign new_n15467_ = ~\all_features[3471]  & ~\all_features[3470]  & ~\all_features[3469]  & ~\all_features[3467]  & ~\all_features[3468] ;
  assign new_n15468_ = ~\all_features[3471]  & (~\all_features[3470]  | (~\all_features[3469]  & ~\all_features[3468]  & (~\all_features[3467]  | ~\all_features[3466] )));
  assign new_n15469_ = ~new_n15470_ & ~new_n15467_;
  assign new_n15470_ = ~new_n15466_ & (new_n15463_ | (~new_n15461_ & (new_n15468_ | (~new_n15464_ & ~new_n15471_))));
  assign new_n15471_ = ~new_n15456_ & (new_n15455_ | (new_n15459_ & (~new_n15458_ | (~new_n15472_ & new_n15448_))));
  assign new_n15472_ = ~\all_features[3469]  & \all_features[3470]  & \all_features[3471]  & (\all_features[3468]  ? new_n15452_ : (new_n15451_ | ~new_n15452_));
  assign new_n15473_ = ~new_n15467_ & ~new_n15466_ & ~new_n15463_ & ~new_n15474_ & ~new_n15461_;
  assign new_n15474_ = ~new_n15464_ & ~new_n15455_ & new_n15475_ & (~new_n15458_ | ~new_n15476_);
  assign new_n15475_ = ~new_n15456_ & ~new_n15468_;
  assign new_n15476_ = new_n15459_ & new_n15448_ & new_n15450_;
  assign new_n15477_ = new_n15460_ & new_n15475_ & ~new_n15467_ & ~new_n15455_ & ~new_n15464_ & ~new_n15466_;
  assign new_n15478_ = ~new_n9379_ & (~new_n9376_ | ~new_n9347_);
  assign new_n15479_ = new_n8668_ & new_n15480_;
  assign new_n15480_ = ~new_n8698_ & ~new_n8701_;
  assign new_n15481_ = ~new_n10972_ & new_n15328_;
  assign new_n15482_ = (~new_n15492_ | ~new_n15483_) & (~new_n15491_ | (new_n15531_ ? ~new_n15496_ : ~new_n15494_));
  assign new_n15483_ = new_n13405_ & ~new_n15478_ & new_n15484_;
  assign new_n15484_ = new_n11120_ & (new_n11097_ | ~new_n15485_);
  assign new_n15485_ = ~new_n15486_ & ~new_n11123_;
  assign new_n15486_ = (new_n15487_ | (new_n11107_ & (~\all_features[3723]  | ~\all_features[3724]  | (~\all_features[3722]  & new_n11106_)))) & (~new_n11107_ | \all_features[3723]  | \all_features[3724] );
  assign new_n15487_ = ~new_n11103_ & (new_n11100_ | (~new_n11114_ & (new_n11117_ | (~new_n15488_ & ~new_n11118_))));
  assign new_n15488_ = ~new_n11116_ & (~\all_features[3727]  | new_n15489_ | (~\all_features[3724]  & ~\all_features[3725]  & ~\all_features[3726] ));
  assign new_n15489_ = \all_features[3727]  & ((~new_n15490_ & ~\all_features[3725]  & \all_features[3726] ) | (~new_n11111_ & (\all_features[3726]  | (~new_n11109_ & \all_features[3725] ))));
  assign new_n15490_ = (\all_features[3724]  & (\all_features[3722]  | \all_features[3723] )) | (~new_n11101_ & ~\all_features[3722]  & ~\all_features[3723]  & ~\all_features[3724] );
  assign new_n15491_ = ~new_n13405_ & ~new_n15407_;
  assign new_n15492_ = new_n15444_ & new_n15493_;
  assign new_n15493_ = new_n15473_ & new_n15477_;
  assign new_n15494_ = new_n15034_ & new_n15495_;
  assign new_n15495_ = ~new_n8192_ & ~new_n8196_;
  assign new_n15496_ = new_n15497_ & new_n15527_;
  assign new_n15497_ = ~new_n15498_ & ~new_n15518_;
  assign new_n15498_ = ~new_n15517_ & (new_n15512_ | (~new_n15514_ & (new_n15515_ | (~new_n15499_ & ~new_n15516_))));
  assign new_n15499_ = ~new_n15506_ & (new_n15509_ | (~new_n15508_ & (~new_n15511_ | new_n15500_)));
  assign new_n15500_ = \all_features[2375]  & ((~new_n15505_ & ~\all_features[2373]  & \all_features[2374] ) | (~new_n15503_ & (\all_features[2374]  | (~new_n15501_ & \all_features[2373] ))));
  assign new_n15501_ = new_n15502_ & ~\all_features[2372]  & ~\all_features[2370]  & ~\all_features[2371] ;
  assign new_n15502_ = ~\all_features[2368]  & ~\all_features[2369] ;
  assign new_n15503_ = \all_features[2375]  & (\all_features[2374]  | (new_n15504_ & (\all_features[2370]  | \all_features[2371]  | \all_features[2369] )));
  assign new_n15504_ = \all_features[2372]  & \all_features[2373] ;
  assign new_n15505_ = (~\all_features[2370]  & ~\all_features[2371]  & ~\all_features[2372]  & (~\all_features[2369]  | ~\all_features[2368] )) | (\all_features[2372]  & (\all_features[2370]  | \all_features[2371] ));
  assign new_n15506_ = ~\all_features[2375]  & (~\all_features[2374]  | (~\all_features[2373]  & (new_n15502_ | ~new_n15507_ | ~\all_features[2372] )));
  assign new_n15507_ = \all_features[2370]  & \all_features[2371] ;
  assign new_n15508_ = ~\all_features[2375]  & (~new_n15507_ | ~\all_features[2368]  | ~\all_features[2369]  | ~\all_features[2374]  | ~new_n15504_);
  assign new_n15509_ = ~new_n15510_ & ~\all_features[2375] ;
  assign new_n15510_ = \all_features[2373]  & \all_features[2374]  & (\all_features[2372]  | (\all_features[2370]  & \all_features[2371]  & \all_features[2369] ));
  assign new_n15511_ = \all_features[2375]  & (\all_features[2373]  | \all_features[2374]  | \all_features[2372] );
  assign new_n15512_ = ~\all_features[2373]  & new_n15513_ & ((~\all_features[2370]  & new_n15502_) | ~\all_features[2372]  | ~\all_features[2371] );
  assign new_n15513_ = ~\all_features[2374]  & ~\all_features[2375] ;
  assign new_n15514_ = new_n15513_ & (~\all_features[2373]  | (~\all_features[2372]  & (~\all_features[2371]  | (~\all_features[2370]  & ~\all_features[2369] ))));
  assign new_n15515_ = new_n15513_ & (~new_n15504_ | ~\all_features[2371]  | (~\all_features[2370]  & (~\all_features[2368]  | ~\all_features[2369] )));
  assign new_n15516_ = ~\all_features[2375]  & (~\all_features[2374]  | (~\all_features[2372]  & ~\all_features[2373]  & ~new_n15507_));
  assign new_n15517_ = ~\all_features[2375]  & ~\all_features[2374]  & ~\all_features[2373]  & ~\all_features[2371]  & ~\all_features[2372] ;
  assign new_n15518_ = new_n15524_ & (~new_n15526_ | (~new_n15516_ & ~new_n15506_ & (~new_n15525_ | new_n15519_)));
  assign new_n15519_ = new_n15520_ & (~new_n15521_ | (~new_n15523_ & \all_features[2373]  & \all_features[2374]  & \all_features[2375] ));
  assign new_n15520_ = \all_features[2375]  & (\all_features[2374]  | (~new_n15501_ & \all_features[2373] ));
  assign new_n15521_ = \all_features[2375]  & \all_features[2374]  & ~new_n15522_ & new_n15503_;
  assign new_n15522_ = ~\all_features[2370]  & ~\all_features[2371]  & ~\all_features[2372]  & ~\all_features[2373]  & (~\all_features[2369]  | ~\all_features[2368] );
  assign new_n15523_ = ~\all_features[2371]  & ~\all_features[2372]  & (~\all_features[2370]  | new_n15502_);
  assign new_n15524_ = ~new_n15512_ & ~new_n15517_;
  assign new_n15525_ = ~new_n15508_ & ~new_n15509_;
  assign new_n15526_ = ~new_n15514_ & ~new_n15515_;
  assign new_n15527_ = ~new_n15528_ & ~new_n15530_;
  assign new_n15528_ = new_n15526_ & ~new_n15529_ & new_n15524_;
  assign new_n15529_ = ~new_n15516_ & ~new_n15506_ & ~new_n15508_ & ~new_n15509_ & (~new_n15521_ | ~new_n15520_);
  assign new_n15530_ = new_n15525_ & new_n15524_ & ~new_n15506_ & ~new_n15516_ & ~new_n15514_ & ~new_n15515_;
  assign new_n15531_ = ~new_n15088_ & ~new_n15352_ & ~new_n15362_;
  assign new_n15532_ = new_n13405_ & ((~new_n15484_ & ~new_n15478_) | (~new_n15533_ & new_n15443_ & new_n15478_));
  assign new_n15533_ = new_n15534_ & (\all_features[5719]  | (~new_n15540_ & \all_features[5717]  & \all_features[5718] ));
  assign new_n15534_ = \all_features[5719]  | (\all_features[5718]  & new_n15535_ & (\all_features[5717]  | (\all_features[5716]  & new_n15537_)));
  assign new_n15535_ = \all_features[5718]  & \all_features[5713]  & new_n15536_ & \all_features[5712] ;
  assign new_n15536_ = \all_features[5717]  & \all_features[5716]  & \all_features[5714]  & \all_features[5715] ;
  assign new_n15537_ = \all_features[5714]  & \all_features[5715]  & (\all_features[5713]  | \all_features[5712] );
  assign new_n15540_ = ~\all_features[5716]  & (~\all_features[5714]  | ~\all_features[5715]  | ~\all_features[5713] );
  assign new_n15541_ = new_n15542_ & (new_n15492_ | ~new_n15483_) & (~new_n15442_ | new_n15481_);
  assign new_n15542_ = new_n13405_ | (new_n15407_ ? (new_n9689_ ? ~new_n14504_ : new_n15479_) : ~new_n15543_);
  assign new_n15543_ = new_n15531_ ? ~new_n15496_ : ~new_n15494_;
  assign new_n15544_ = new_n15545_ & (~new_n15631_ | ~new_n15629_);
  assign new_n15545_ = ~new_n15546_ & new_n15590_ & (new_n12946_ | new_n14654_ | ~new_n15597_);
  assign new_n15546_ = ~new_n15553_ & (new_n15547_ | (~new_n15588_ & ~new_n12946_ & new_n14654_));
  assign new_n15547_ = new_n15548_ & new_n15551_;
  assign new_n15548_ = ~new_n15549_ & new_n12946_;
  assign new_n15549_ = ~new_n11413_ & new_n15550_;
  assign new_n15550_ = ~new_n11444_ & ~new_n11433_ & ~new_n11442_;
  assign new_n15551_ = new_n15552_ & new_n14528_;
  assign new_n15552_ = new_n14505_ & new_n14531_;
  assign new_n15553_ = new_n15554_ & new_n15587_;
  assign new_n15554_ = new_n15555_ & new_n15584_;
  assign new_n15555_ = new_n15556_ & new_n15577_;
  assign new_n15556_ = ~new_n15557_ & (\all_features[4155]  | \all_features[4156]  | \all_features[4157]  | \all_features[4158]  | \all_features[4159] );
  assign new_n15557_ = ~new_n15573_ & (new_n15571_ | (~new_n15575_ & (new_n15576_ | (~new_n15574_ & ~new_n15558_))));
  assign new_n15558_ = ~new_n15559_ & (new_n15561_ | (new_n15570_ & (~new_n15565_ | (~new_n15569_ & new_n15568_))));
  assign new_n15559_ = ~new_n15560_ & ~\all_features[4159] ;
  assign new_n15560_ = \all_features[4157]  & \all_features[4158]  & (\all_features[4156]  | (\all_features[4154]  & \all_features[4155]  & \all_features[4153] ));
  assign new_n15561_ = ~\all_features[4159]  & (~\all_features[4158]  | ~new_n15562_ | ~new_n15563_ | ~new_n15564_);
  assign new_n15562_ = \all_features[4154]  & \all_features[4155] ;
  assign new_n15563_ = \all_features[4152]  & \all_features[4153] ;
  assign new_n15564_ = \all_features[4156]  & \all_features[4157] ;
  assign new_n15565_ = \all_features[4159]  & (\all_features[4158]  | (\all_features[4157]  & (\all_features[4156]  | ~new_n15567_ | ~new_n15566_)));
  assign new_n15566_ = ~\all_features[4152]  & ~\all_features[4153] ;
  assign new_n15567_ = ~\all_features[4154]  & ~\all_features[4155] ;
  assign new_n15568_ = \all_features[4159]  & (\all_features[4158]  | (new_n15564_ & (\all_features[4154]  | \all_features[4155]  | \all_features[4153] )));
  assign new_n15569_ = ~\all_features[4157]  & \all_features[4158]  & \all_features[4159]  & (\all_features[4156]  ? new_n15567_ : (new_n15563_ | ~new_n15567_));
  assign new_n15570_ = \all_features[4159]  & (\all_features[4157]  | \all_features[4158]  | \all_features[4156] );
  assign new_n15571_ = new_n15572_ & (~\all_features[4157]  | (~\all_features[4156]  & (~\all_features[4155]  | (~\all_features[4154]  & ~\all_features[4153] ))));
  assign new_n15572_ = ~\all_features[4158]  & ~\all_features[4159] ;
  assign new_n15573_ = ~\all_features[4157]  & new_n15572_ & ((~\all_features[4154]  & new_n15566_) | ~\all_features[4156]  | ~\all_features[4155] );
  assign new_n15574_ = ~\all_features[4159]  & (~\all_features[4158]  | (~\all_features[4157]  & (new_n15566_ | ~new_n15562_ | ~\all_features[4156] )));
  assign new_n15575_ = new_n15572_ & (~\all_features[4155]  | ~new_n15564_ | (~\all_features[4154]  & ~new_n15563_));
  assign new_n15576_ = ~\all_features[4159]  & (~\all_features[4158]  | (~\all_features[4156]  & ~\all_features[4157]  & ~new_n15562_));
  assign new_n15577_ = new_n15582_ & (~new_n15583_ | (~new_n15578_ & ~new_n15574_ & ~new_n15576_));
  assign new_n15578_ = ~new_n15559_ & ~new_n15561_ & (~new_n15570_ | ~new_n15565_ | new_n15579_);
  assign new_n15579_ = new_n15568_ & new_n15580_ & (new_n15581_ | ~\all_features[4157]  | ~\all_features[4158]  | ~\all_features[4159] );
  assign new_n15580_ = \all_features[4158]  & \all_features[4159]  & (\all_features[4156]  | \all_features[4157]  | new_n15563_ | ~new_n15567_);
  assign new_n15581_ = ~\all_features[4155]  & ~\all_features[4156]  & (~\all_features[4154]  | new_n15566_);
  assign new_n15582_ = ~new_n15573_ & (\all_features[4155]  | \all_features[4156]  | \all_features[4157]  | \all_features[4158]  | \all_features[4159] );
  assign new_n15583_ = ~new_n15571_ & ~new_n15575_;
  assign new_n15584_ = new_n15582_ & new_n15583_ & (new_n15586_ | new_n15559_ | new_n15574_ | ~new_n15585_);
  assign new_n15585_ = ~new_n15561_ & ~new_n15576_;
  assign new_n15586_ = new_n15570_ & new_n15580_ & new_n15565_ & new_n15568_;
  assign new_n15587_ = new_n15585_ & new_n15582_ & ~new_n15575_ & ~new_n15574_ & ~new_n15559_ & ~new_n15571_;
  assign new_n15588_ = new_n14813_ & new_n15589_;
  assign new_n15589_ = ~new_n14843_ & ~new_n14845_;
  assign new_n15590_ = ~new_n15591_ | (new_n15592_ ? new_n15594_ : new_n15595_);
  assign new_n15591_ = new_n15549_ & new_n12946_;
  assign new_n15592_ = ~new_n15593_ & new_n8806_;
  assign new_n15593_ = new_n8778_ & new_n8802_;
  assign new_n15594_ = ~new_n13095_ & (~new_n13067_ | new_n13517_);
  assign new_n15595_ = ~new_n10389_ & new_n15596_;
  assign new_n15596_ = ~new_n8391_ & ~new_n10395_;
  assign new_n15597_ = new_n15598_ & (~new_n11857_ | ~new_n11854_);
  assign new_n15598_ = ~new_n15628_ & new_n15599_;
  assign new_n15599_ = ~new_n15600_ & ~new_n15623_;
  assign new_n15600_ = ~new_n15622_ & ~new_n15621_ & ~new_n15620_ & ~new_n15601_ & ~new_n15618_;
  assign new_n15601_ = ~new_n15602_ & ~new_n15616_ & new_n15605_ & (~new_n15617_ | ~new_n15609_);
  assign new_n15602_ = ~\all_features[5071]  & (~\all_features[5070]  | new_n15603_);
  assign new_n15603_ = ~\all_features[5069]  & (new_n15604_ | ~\all_features[5067]  | ~\all_features[5068]  | ~\all_features[5066] );
  assign new_n15604_ = ~\all_features[5064]  & ~\all_features[5065] ;
  assign new_n15605_ = ~new_n15606_ & ~new_n15608_;
  assign new_n15606_ = ~new_n15607_ & ~\all_features[5071] ;
  assign new_n15607_ = \all_features[5069]  & \all_features[5070]  & (\all_features[5068]  | (\all_features[5066]  & \all_features[5067]  & \all_features[5065] ));
  assign new_n15608_ = ~\all_features[5071]  & (~\all_features[5070]  | (~\all_features[5069]  & ~\all_features[5068]  & (~\all_features[5067]  | ~\all_features[5066] )));
  assign new_n15609_ = new_n15615_ & new_n15610_ & new_n15612_;
  assign new_n15610_ = \all_features[5071]  & (\all_features[5070]  | (new_n15611_ & (\all_features[5066]  | \all_features[5067]  | \all_features[5065] )));
  assign new_n15611_ = \all_features[5068]  & \all_features[5069] ;
  assign new_n15612_ = \all_features[5070]  & \all_features[5071]  & (\all_features[5068]  | \all_features[5069]  | new_n15613_ | ~new_n15614_);
  assign new_n15613_ = \all_features[5064]  & \all_features[5065] ;
  assign new_n15614_ = ~\all_features[5066]  & ~\all_features[5067] ;
  assign new_n15615_ = \all_features[5071]  & (\all_features[5069]  | \all_features[5070]  | \all_features[5068] );
  assign new_n15616_ = ~\all_features[5071]  & (~new_n15611_ | ~\all_features[5066]  | ~\all_features[5067]  | ~\all_features[5070]  | ~new_n15613_);
  assign new_n15617_ = \all_features[5071]  & (\all_features[5070]  | (\all_features[5069]  & (\all_features[5068]  | ~new_n15614_ | ~new_n15604_)));
  assign new_n15618_ = new_n15619_ & (~\all_features[5067]  | ~new_n15611_ | (~\all_features[5066]  & ~new_n15613_));
  assign new_n15619_ = ~\all_features[5070]  & ~\all_features[5071] ;
  assign new_n15620_ = new_n15619_ & (~\all_features[5069]  | (~\all_features[5068]  & (~\all_features[5067]  | (~\all_features[5066]  & ~\all_features[5065] ))));
  assign new_n15621_ = ~\all_features[5069]  & new_n15619_ & ((~\all_features[5066]  & new_n15604_) | ~\all_features[5068]  | ~\all_features[5067] );
  assign new_n15622_ = ~\all_features[5071]  & ~\all_features[5070]  & ~\all_features[5069]  & ~\all_features[5067]  & ~\all_features[5068] ;
  assign new_n15623_ = ~new_n15622_ & ~new_n15621_ & (~new_n15627_ | (~new_n15624_ & ~new_n15602_ & ~new_n15608_));
  assign new_n15624_ = ~new_n15616_ & ~new_n15606_ & (~new_n15615_ | ~new_n15617_ | new_n15625_);
  assign new_n15625_ = new_n15610_ & new_n15612_ & (new_n15626_ | ~\all_features[5069]  | ~\all_features[5070]  | ~\all_features[5071] );
  assign new_n15626_ = ~\all_features[5067]  & ~\all_features[5068]  & (~\all_features[5066]  | new_n15604_);
  assign new_n15627_ = ~new_n15618_ & ~new_n15620_;
  assign new_n15628_ = new_n15627_ & new_n15605_ & ~new_n15622_ & ~new_n15616_ & ~new_n15602_ & ~new_n15621_;
  assign new_n15629_ = new_n15630_ & (~new_n15591_ | (~new_n15594_ & new_n15592_) | (~new_n15595_ & ~new_n15592_));
  assign new_n15630_ = (~new_n15553_ | (~new_n15547_ & (new_n12946_ | ~new_n14654_))) & (new_n12946_ | (new_n14654_ ? ~new_n15588_ : new_n15597_));
  assign new_n15631_ = ~new_n15551_ & ~new_n15664_ & new_n15548_ & (~new_n15632_ | (~new_n15656_ & ~new_n15660_));
  assign new_n15632_ = new_n15653_ & ~new_n15633_ & new_n15649_;
  assign new_n15633_ = new_n15634_ & (~new_n15647_ | ~new_n15648_ | ~new_n15644_ | ~new_n15646_);
  assign new_n15634_ = ~new_n15643_ & ~new_n15640_ & ~new_n15635_ & ~new_n15638_;
  assign new_n15635_ = ~\all_features[4447]  & (~\all_features[4446]  | (~\all_features[4445]  & (new_n15636_ | ~new_n15637_ | ~\all_features[4444] )));
  assign new_n15636_ = ~\all_features[4440]  & ~\all_features[4441] ;
  assign new_n15637_ = \all_features[4442]  & \all_features[4443] ;
  assign new_n15638_ = ~new_n15639_ & ~\all_features[4447] ;
  assign new_n15639_ = \all_features[4445]  & \all_features[4446]  & (\all_features[4444]  | (\all_features[4442]  & \all_features[4443]  & \all_features[4441] ));
  assign new_n15640_ = ~\all_features[4447]  & (~\all_features[4446]  | ~new_n15641_ | ~new_n15642_ | ~new_n15637_);
  assign new_n15641_ = \all_features[4444]  & \all_features[4445] ;
  assign new_n15642_ = \all_features[4440]  & \all_features[4441] ;
  assign new_n15643_ = ~\all_features[4447]  & (~\all_features[4446]  | (~\all_features[4444]  & ~\all_features[4445]  & ~new_n15637_));
  assign new_n15644_ = \all_features[4447]  & (\all_features[4446]  | (\all_features[4445]  & (\all_features[4444]  | ~new_n15636_ | ~new_n15645_)));
  assign new_n15645_ = ~\all_features[4442]  & ~\all_features[4443] ;
  assign new_n15646_ = \all_features[4447]  & (\all_features[4446]  | (new_n15641_ & (\all_features[4442]  | \all_features[4443]  | \all_features[4441] )));
  assign new_n15647_ = \all_features[4446]  & \all_features[4447]  & (\all_features[4444]  | \all_features[4445]  | new_n15642_ | ~new_n15645_);
  assign new_n15648_ = \all_features[4447]  & (\all_features[4445]  | \all_features[4446]  | \all_features[4444] );
  assign new_n15649_ = ~new_n15650_ & ~new_n15652_;
  assign new_n15650_ = ~\all_features[4445]  & new_n15651_ & ((~\all_features[4442]  & new_n15636_) | ~\all_features[4444]  | ~\all_features[4443] );
  assign new_n15651_ = ~\all_features[4446]  & ~\all_features[4447] ;
  assign new_n15652_ = ~\all_features[4447]  & ~\all_features[4446]  & ~\all_features[4445]  & ~\all_features[4443]  & ~\all_features[4444] ;
  assign new_n15653_ = ~new_n15654_ & ~new_n15655_;
  assign new_n15654_ = new_n15651_ & (~\all_features[4445]  | (~\all_features[4444]  & (~\all_features[4443]  | (~\all_features[4442]  & ~\all_features[4441] ))));
  assign new_n15655_ = new_n15651_ & (~\all_features[4443]  | ~new_n15641_ | (~\all_features[4442]  & ~new_n15642_));
  assign new_n15656_ = new_n15649_ & (~new_n15653_ | (~new_n15657_ & ~new_n15635_ & ~new_n15643_));
  assign new_n15657_ = ~new_n15640_ & ~new_n15638_ & (~new_n15648_ | ~new_n15644_ | new_n15658_);
  assign new_n15658_ = new_n15646_ & new_n15647_ & (new_n15659_ | ~\all_features[4445]  | ~\all_features[4446]  | ~\all_features[4447] );
  assign new_n15659_ = ~\all_features[4443]  & ~\all_features[4444]  & (~\all_features[4442]  | new_n15636_);
  assign new_n15660_ = ~new_n15661_ & ~new_n15652_;
  assign new_n15661_ = ~new_n15650_ & (new_n15654_ | (~new_n15655_ & (new_n15643_ | (~new_n15635_ & ~new_n15662_))));
  assign new_n15662_ = ~new_n15638_ & (new_n15640_ | (new_n15648_ & (~new_n15644_ | (~new_n15663_ & new_n15646_))));
  assign new_n15663_ = ~\all_features[4445]  & \all_features[4446]  & \all_features[4447]  & (\all_features[4444]  ? new_n15645_ : (new_n15642_ | ~new_n15645_));
  assign new_n15664_ = new_n15665_ & ~new_n15655_ & ~new_n15650_ & ~new_n15635_ & ~new_n15643_;
  assign new_n15665_ = ~new_n15652_ & ~new_n15654_ & ~new_n15638_ & ~new_n15640_;
  assign new_n15666_ = (new_n15670_ | new_n9689_ | new_n15707_) & (new_n15667_ | (~new_n9689_ & (new_n15674_ | new_n14330_ | ~new_n15707_)));
  assign new_n15667_ = ~new_n15669_ & new_n9689_ & (new_n14154_ | new_n15668_);
  assign new_n15668_ = ~new_n10970_ & (~new_n10949_ | new_n15321_);
  assign new_n15669_ = ~new_n14160_ & new_n10999_;
  assign new_n15670_ = new_n15671_ ? ~new_n15673_ : new_n7408_;
  assign new_n15671_ = new_n8099_ & new_n15672_;
  assign new_n15672_ = new_n8129_ & new_n8132_;
  assign new_n15673_ = ~new_n9129_ & (~new_n9131_ | new_n12448_);
  assign new_n15674_ = ~new_n15703_ & new_n15675_;
  assign new_n15675_ = ~new_n15676_ & ~new_n15702_;
  assign new_n15676_ = new_n15689_ & (~new_n15677_ | (new_n15700_ & new_n15701_ & new_n15697_ & new_n15698_));
  assign new_n15677_ = new_n15678_ & new_n15685_;
  assign new_n15678_ = ~new_n15679_ & ~new_n15681_;
  assign new_n15679_ = ~new_n15680_ & ~\all_features[2151] ;
  assign new_n15680_ = \all_features[2149]  & \all_features[2150]  & (\all_features[2148]  | (\all_features[2146]  & \all_features[2147]  & \all_features[2145] ));
  assign new_n15681_ = ~\all_features[2151]  & (~\all_features[2150]  | ~new_n15682_ | ~new_n15683_ | ~new_n15684_);
  assign new_n15682_ = \all_features[2148]  & \all_features[2149] ;
  assign new_n15683_ = \all_features[2144]  & \all_features[2145] ;
  assign new_n15684_ = \all_features[2146]  & \all_features[2147] ;
  assign new_n15685_ = ~new_n15686_ & ~new_n15687_;
  assign new_n15686_ = ~\all_features[2151]  & (~\all_features[2150]  | (~\all_features[2148]  & ~\all_features[2149]  & ~new_n15684_));
  assign new_n15687_ = ~\all_features[2151]  & (~\all_features[2150]  | (~\all_features[2149]  & (new_n15688_ | ~new_n15684_ | ~\all_features[2148] )));
  assign new_n15688_ = ~\all_features[2144]  & ~\all_features[2145] ;
  assign new_n15689_ = new_n15690_ & new_n15694_;
  assign new_n15690_ = ~new_n15691_ & ~new_n15693_;
  assign new_n15691_ = new_n15692_ & (~\all_features[2149]  | (~\all_features[2148]  & (~\all_features[2147]  | (~\all_features[2146]  & ~\all_features[2145] ))));
  assign new_n15692_ = ~\all_features[2150]  & ~\all_features[2151] ;
  assign new_n15693_ = new_n15692_ & (~\all_features[2147]  | ~new_n15682_ | (~\all_features[2146]  & ~new_n15683_));
  assign new_n15694_ = ~new_n15695_ & ~new_n15696_;
  assign new_n15695_ = ~\all_features[2149]  & new_n15692_ & ((~\all_features[2146]  & new_n15688_) | ~\all_features[2148]  | ~\all_features[2147] );
  assign new_n15696_ = ~\all_features[2151]  & ~\all_features[2150]  & ~\all_features[2149]  & ~\all_features[2147]  & ~\all_features[2148] ;
  assign new_n15697_ = \all_features[2151]  & (\all_features[2150]  | (new_n15682_ & (\all_features[2146]  | \all_features[2147]  | \all_features[2145] )));
  assign new_n15698_ = \all_features[2150]  & \all_features[2151]  & (\all_features[2148]  | \all_features[2149]  | new_n15683_ | ~new_n15699_);
  assign new_n15699_ = ~\all_features[2146]  & ~\all_features[2147] ;
  assign new_n15700_ = \all_features[2151]  & (\all_features[2150]  | (\all_features[2149]  & (\all_features[2148]  | ~new_n15699_ | ~new_n15688_)));
  assign new_n15701_ = \all_features[2151]  & (\all_features[2149]  | \all_features[2150]  | \all_features[2148] );
  assign new_n15702_ = new_n15677_ & new_n15689_;
  assign new_n15703_ = new_n15694_ & (~new_n15690_ | (~new_n15704_ & new_n15685_));
  assign new_n15704_ = new_n15678_ & ((~new_n15705_ & new_n15698_ & new_n15697_) | ~new_n15701_ | ~new_n15700_);
  assign new_n15705_ = \all_features[2151]  & \all_features[2150]  & ~new_n15706_ & \all_features[2149] ;
  assign new_n15706_ = ~\all_features[2147]  & ~\all_features[2148]  & (~\all_features[2146]  | new_n15688_);
  assign new_n15707_ = ~new_n6566_ & (~new_n6563_ | ~new_n6556_);
  assign new_n15708_ = new_n15709_ ? (new_n15759_ ^ new_n15865_) : (~new_n15759_ ^ new_n15865_);
  assign new_n15709_ = ~new_n15710_ & new_n15758_;
  assign new_n15710_ = new_n15711_ & (new_n14461_ | ((new_n15755_ | ~new_n15752_) & (new_n15757_ | new_n11750_ | new_n15752_)));
  assign new_n15711_ = new_n15712_ & (new_n14461_ | ~new_n11750_ | ~new_n9686_ | new_n15752_) & (~new_n15754_ | ~new_n15752_);
  assign new_n15712_ = ~new_n14461_ | (new_n15751_ ? ~new_n15715_ : ~new_n15713_);
  assign new_n15713_ = ~new_n15714_ & new_n12486_;
  assign new_n15714_ = ~new_n12455_ & ~new_n12476_;
  assign new_n15715_ = new_n15716_ & new_n15747_;
  assign new_n15716_ = new_n15745_ & new_n15717_ & new_n15743_;
  assign new_n15717_ = ~new_n15741_ & ~new_n15742_ & (~new_n15734_ | (~new_n15718_ & new_n15738_));
  assign new_n15718_ = new_n15719_ & ((~new_n15726_ & new_n15730_ & new_n15729_) | ~new_n15733_ | ~new_n15732_);
  assign new_n15719_ = ~new_n15720_ & ~new_n15724_;
  assign new_n15720_ = ~\all_features[2167]  & (~\all_features[2166]  | ~new_n15721_ | ~new_n15722_ | ~new_n15723_);
  assign new_n15721_ = \all_features[2160]  & \all_features[2161] ;
  assign new_n15722_ = \all_features[2164]  & \all_features[2165] ;
  assign new_n15723_ = \all_features[2162]  & \all_features[2163] ;
  assign new_n15724_ = ~new_n15725_ & ~\all_features[2167] ;
  assign new_n15725_ = \all_features[2165]  & \all_features[2166]  & (\all_features[2164]  | (\all_features[2162]  & \all_features[2163]  & \all_features[2161] ));
  assign new_n15726_ = \all_features[2167]  & \all_features[2166]  & ~new_n15727_ & \all_features[2165] ;
  assign new_n15727_ = ~\all_features[2163]  & ~\all_features[2164]  & (~\all_features[2162]  | new_n15728_);
  assign new_n15728_ = ~\all_features[2160]  & ~\all_features[2161] ;
  assign new_n15729_ = \all_features[2167]  & (\all_features[2166]  | (new_n15722_ & (\all_features[2162]  | \all_features[2163]  | \all_features[2161] )));
  assign new_n15730_ = \all_features[2166]  & \all_features[2167]  & (\all_features[2164]  | \all_features[2165]  | new_n15721_ | ~new_n15731_);
  assign new_n15731_ = ~\all_features[2162]  & ~\all_features[2163] ;
  assign new_n15732_ = \all_features[2167]  & (\all_features[2166]  | (\all_features[2165]  & (\all_features[2164]  | ~new_n15731_ | ~new_n15728_)));
  assign new_n15733_ = \all_features[2167]  & (\all_features[2165]  | \all_features[2166]  | \all_features[2164] );
  assign new_n15734_ = ~new_n15735_ & ~new_n15737_;
  assign new_n15735_ = new_n15736_ & (~\all_features[2165]  | (~\all_features[2164]  & (~\all_features[2163]  | (~\all_features[2162]  & ~\all_features[2161] ))));
  assign new_n15736_ = ~\all_features[2166]  & ~\all_features[2167] ;
  assign new_n15737_ = new_n15736_ & (~\all_features[2163]  | ~new_n15722_ | (~\all_features[2162]  & ~new_n15721_));
  assign new_n15738_ = ~new_n15739_ & ~new_n15740_;
  assign new_n15739_ = ~\all_features[2167]  & (~\all_features[2166]  | (~\all_features[2165]  & (new_n15728_ | ~new_n15723_ | ~\all_features[2164] )));
  assign new_n15740_ = ~\all_features[2167]  & (~\all_features[2166]  | (~\all_features[2164]  & ~\all_features[2165]  & ~new_n15723_));
  assign new_n15741_ = ~\all_features[2165]  & new_n15736_ & ((~\all_features[2162]  & new_n15728_) | ~\all_features[2164]  | ~\all_features[2163] );
  assign new_n15742_ = ~\all_features[2167]  & ~\all_features[2166]  & ~\all_features[2165]  & ~\all_features[2163]  & ~\all_features[2164] ;
  assign new_n15743_ = ~new_n15742_ & ~new_n15741_ & ~new_n15737_ & ~new_n15744_ & ~new_n15735_;
  assign new_n15744_ = new_n15738_ & new_n15719_ & (~new_n15732_ | ~new_n15733_ | ~new_n15729_ | ~new_n15730_);
  assign new_n15745_ = new_n15746_ & new_n15734_ & ~new_n15741_ & ~new_n15724_ & ~new_n15739_ & ~new_n15740_;
  assign new_n15746_ = ~new_n15720_ & ~new_n15742_;
  assign new_n15747_ = ~new_n15748_ & ~new_n15742_;
  assign new_n15748_ = ~new_n15741_ & (new_n15735_ | (~new_n15737_ & (new_n15740_ | (~new_n15739_ & ~new_n15749_))));
  assign new_n15749_ = ~new_n15724_ & (new_n15720_ | (new_n15733_ & (~new_n15732_ | (~new_n15750_ & new_n15729_))));
  assign new_n15750_ = ~\all_features[2165]  & \all_features[2166]  & \all_features[2167]  & (\all_features[2164]  ? new_n15731_ : (new_n15721_ | ~new_n15731_));
  assign new_n15751_ = new_n14921_ & ~new_n14243_ & ~new_n14269_;
  assign new_n15752_ = ~new_n8391_ & (~new_n10395_ | new_n15753_);
  assign new_n15753_ = ~new_n10381_ & ~new_n10389_;
  assign new_n15754_ = ~new_n14461_ & new_n10999_ & new_n15755_ & (new_n10977_ | new_n15756_);
  assign new_n15755_ = new_n15600_ & new_n15628_;
  assign new_n15756_ = new_n13320_ & new_n13324_;
  assign new_n15757_ = new_n6391_ & new_n8390_;
  assign new_n15758_ = (~new_n15751_ | new_n15715_ | ~new_n14461_) & (new_n15752_ | new_n11750_ | ~new_n15757_ | new_n14461_);
  assign new_n15759_ = ~new_n15829_ & (new_n15830_ | (new_n15760_ & (new_n15821_ | new_n15752_ | new_n13982_)));
  assign new_n15760_ = new_n13982_ ? new_n15761_ : (~new_n15821_ | (new_n15828_ & new_n14540_));
  assign new_n15761_ = (~new_n8891_ & (~new_n15819_ | ~new_n15797_)) | (new_n15788_ & new_n15762_ & new_n8891_);
  assign new_n15762_ = new_n15763_ & new_n15786_;
  assign new_n15763_ = new_n15781_ & ~new_n15785_ & ~new_n15764_ & ~new_n15784_;
  assign new_n15764_ = ~new_n15779_ & ~new_n15780_ & new_n15772_ & (~new_n15777_ | ~new_n15765_);
  assign new_n15765_ = new_n15771_ & new_n15766_ & new_n15768_;
  assign new_n15766_ = \all_features[3495]  & (\all_features[3494]  | (new_n15767_ & (\all_features[3490]  | \all_features[3491]  | \all_features[3489] )));
  assign new_n15767_ = \all_features[3492]  & \all_features[3493] ;
  assign new_n15768_ = \all_features[3494]  & \all_features[3495]  & (\all_features[3492]  | \all_features[3493]  | new_n15770_ | ~new_n15769_);
  assign new_n15769_ = ~\all_features[3490]  & ~\all_features[3491] ;
  assign new_n15770_ = \all_features[3488]  & \all_features[3489] ;
  assign new_n15771_ = \all_features[3495]  & (\all_features[3493]  | \all_features[3494]  | \all_features[3492] );
  assign new_n15772_ = ~new_n15773_ & ~new_n15775_;
  assign new_n15773_ = ~new_n15774_ & ~\all_features[3495] ;
  assign new_n15774_ = \all_features[3493]  & \all_features[3494]  & (\all_features[3492]  | (\all_features[3490]  & \all_features[3491]  & \all_features[3489] ));
  assign new_n15775_ = ~\all_features[3495]  & (~\all_features[3494]  | (~\all_features[3492]  & ~\all_features[3493]  & ~new_n15776_));
  assign new_n15776_ = \all_features[3490]  & \all_features[3491] ;
  assign new_n15777_ = \all_features[3495]  & (\all_features[3494]  | (\all_features[3493]  & (\all_features[3492]  | ~new_n15778_ | ~new_n15769_)));
  assign new_n15778_ = ~\all_features[3488]  & ~\all_features[3489] ;
  assign new_n15779_ = ~\all_features[3495]  & (~\all_features[3494]  | (~\all_features[3493]  & (new_n15778_ | ~new_n15776_ | ~\all_features[3492] )));
  assign new_n15780_ = ~\all_features[3495]  & (~\all_features[3494]  | ~new_n15767_ | ~new_n15770_ | ~new_n15776_);
  assign new_n15781_ = ~new_n15782_ & (\all_features[3491]  | \all_features[3492]  | \all_features[3493]  | \all_features[3494]  | \all_features[3495] );
  assign new_n15782_ = ~\all_features[3493]  & new_n15783_ & ((~\all_features[3490]  & new_n15778_) | ~\all_features[3492]  | ~\all_features[3491] );
  assign new_n15783_ = ~\all_features[3494]  & ~\all_features[3495] ;
  assign new_n15784_ = new_n15783_ & (~\all_features[3493]  | (~\all_features[3492]  & (~\all_features[3491]  | (~\all_features[3490]  & ~\all_features[3489] ))));
  assign new_n15785_ = new_n15783_ & (~\all_features[3491]  | ~new_n15767_ | (~\all_features[3490]  & ~new_n15770_));
  assign new_n15786_ = new_n15781_ & new_n15772_ & new_n15787_ & ~new_n15779_ & ~new_n15780_;
  assign new_n15787_ = ~new_n15784_ & ~new_n15785_;
  assign new_n15788_ = new_n15789_ & new_n15793_;
  assign new_n15789_ = ~new_n15790_ & (\all_features[3491]  | \all_features[3492]  | \all_features[3493]  | \all_features[3494]  | \all_features[3495] );
  assign new_n15790_ = ~new_n15782_ & (new_n15784_ | (~new_n15785_ & (new_n15775_ | (~new_n15779_ & ~new_n15791_))));
  assign new_n15791_ = ~new_n15773_ & (new_n15780_ | (new_n15771_ & (~new_n15777_ | (~new_n15792_ & new_n15766_))));
  assign new_n15792_ = ~\all_features[3493]  & \all_features[3494]  & \all_features[3495]  & (\all_features[3492]  ? new_n15769_ : (new_n15770_ | ~new_n15769_));
  assign new_n15793_ = new_n15781_ & (~new_n15787_ | (~new_n15794_ & ~new_n15775_ & ~new_n15779_));
  assign new_n15794_ = ~new_n15780_ & ~new_n15773_ & (~new_n15771_ | ~new_n15777_ | new_n15795_);
  assign new_n15795_ = new_n15766_ & new_n15768_ & (new_n15796_ | ~\all_features[3493]  | ~\all_features[3494]  | ~\all_features[3495] );
  assign new_n15796_ = ~\all_features[3491]  & ~\all_features[3492]  & (~\all_features[3490]  | new_n15778_);
  assign new_n15797_ = new_n15814_ & ~new_n15818_ & ~new_n15798_ & ~new_n15817_;
  assign new_n15798_ = new_n15799_ & (~new_n15812_ | ~new_n15813_ | ~new_n15809_ | ~new_n15811_);
  assign new_n15799_ = ~new_n15806_ & ~new_n15805_ & ~new_n15800_ & ~new_n15803_;
  assign new_n15800_ = ~\all_features[991]  & (~\all_features[990]  | (~\all_features[989]  & (new_n15801_ | ~new_n15802_ | ~\all_features[988] )));
  assign new_n15801_ = ~\all_features[984]  & ~\all_features[985] ;
  assign new_n15802_ = \all_features[986]  & \all_features[987] ;
  assign new_n15803_ = ~new_n15804_ & ~\all_features[991] ;
  assign new_n15804_ = \all_features[989]  & \all_features[990]  & (\all_features[988]  | (\all_features[986]  & \all_features[987]  & \all_features[985] ));
  assign new_n15805_ = ~\all_features[991]  & (~\all_features[990]  | (~\all_features[988]  & ~\all_features[989]  & ~new_n15802_));
  assign new_n15806_ = ~\all_features[991]  & (~\all_features[990]  | ~new_n15807_ | ~new_n15808_ | ~new_n15802_);
  assign new_n15807_ = \all_features[988]  & \all_features[989] ;
  assign new_n15808_ = \all_features[984]  & \all_features[985] ;
  assign new_n15809_ = \all_features[991]  & (\all_features[990]  | (\all_features[989]  & (\all_features[988]  | ~new_n15801_ | ~new_n15810_)));
  assign new_n15810_ = ~\all_features[986]  & ~\all_features[987] ;
  assign new_n15811_ = \all_features[991]  & (\all_features[990]  | (new_n15807_ & (\all_features[986]  | \all_features[987]  | \all_features[985] )));
  assign new_n15812_ = \all_features[990]  & \all_features[991]  & (\all_features[988]  | \all_features[989]  | new_n15808_ | ~new_n15810_);
  assign new_n15813_ = \all_features[991]  & (\all_features[989]  | \all_features[990]  | \all_features[988] );
  assign new_n15814_ = ~new_n15815_ & (\all_features[987]  | \all_features[988]  | \all_features[989]  | \all_features[990]  | \all_features[991] );
  assign new_n15815_ = ~\all_features[989]  & new_n15816_ & ((~\all_features[986]  & new_n15801_) | ~\all_features[988]  | ~\all_features[987] );
  assign new_n15816_ = ~\all_features[990]  & ~\all_features[991] ;
  assign new_n15817_ = new_n15816_ & (~\all_features[989]  | (~\all_features[988]  & (~\all_features[987]  | (~\all_features[986]  & ~\all_features[985] ))));
  assign new_n15818_ = new_n15816_ & (~\all_features[987]  | ~new_n15807_ | (~\all_features[986]  & ~new_n15808_));
  assign new_n15819_ = new_n15820_ & new_n15814_ & ~new_n15803_ & ~new_n15817_;
  assign new_n15820_ = ~new_n15818_ & ~new_n15806_ & ~new_n15800_ & ~new_n15805_;
  assign new_n15821_ = new_n15017_ & (new_n14990_ | new_n15822_);
  assign new_n15822_ = new_n15823_ & new_n15013_;
  assign new_n15823_ = ~new_n15009_ & (new_n15006_ | (~new_n15012_ & (new_n15011_ | (~new_n14999_ & ~new_n15824_))));
  assign new_n15824_ = ~new_n15001_ & (new_n15002_ | (~new_n15004_ & (~new_n15827_ | new_n15825_)));
  assign new_n15825_ = \all_features[791]  & ((~new_n15826_ & ~\all_features[789]  & \all_features[790] ) | (~new_n14996_ & (\all_features[790]  | (~new_n14993_ & \all_features[789] ))));
  assign new_n15826_ = (~\all_features[786]  & ~\all_features[787]  & ~\all_features[788]  & (~\all_features[785]  | ~\all_features[784] )) | (\all_features[788]  & (\all_features[786]  | \all_features[787] ));
  assign new_n15827_ = \all_features[791]  & (\all_features[789]  | \all_features[790]  | \all_features[788] );
  assign new_n15828_ = ~new_n6675_ & ~new_n6698_;
  assign new_n15829_ = new_n15864_ & ~new_n11260_ & new_n15830_;
  assign new_n15830_ = new_n15860_ & (new_n15862_ | ~new_n15831_);
  assign new_n15831_ = ~new_n15832_ & ~new_n15853_;
  assign new_n15832_ = ~new_n15833_ & (\all_features[2531]  | \all_features[2532]  | \all_features[2533]  | \all_features[2534]  | \all_features[2535] );
  assign new_n15833_ = ~new_n15849_ & (new_n15847_ | (~new_n15851_ & (new_n15852_ | (~new_n15850_ & ~new_n15834_))));
  assign new_n15834_ = ~new_n15835_ & (new_n15837_ | (new_n15846_ & (~new_n15841_ | (~new_n15845_ & new_n15844_))));
  assign new_n15835_ = ~new_n15836_ & ~\all_features[2535] ;
  assign new_n15836_ = \all_features[2533]  & \all_features[2534]  & (\all_features[2532]  | (\all_features[2530]  & \all_features[2531]  & \all_features[2529] ));
  assign new_n15837_ = ~\all_features[2535]  & (~\all_features[2534]  | ~new_n15838_ | ~new_n15839_ | ~new_n15840_);
  assign new_n15838_ = \all_features[2530]  & \all_features[2531] ;
  assign new_n15839_ = \all_features[2528]  & \all_features[2529] ;
  assign new_n15840_ = \all_features[2532]  & \all_features[2533] ;
  assign new_n15841_ = \all_features[2535]  & (\all_features[2534]  | (\all_features[2533]  & (\all_features[2532]  | ~new_n15843_ | ~new_n15842_)));
  assign new_n15842_ = ~\all_features[2528]  & ~\all_features[2529] ;
  assign new_n15843_ = ~\all_features[2530]  & ~\all_features[2531] ;
  assign new_n15844_ = \all_features[2535]  & (\all_features[2534]  | (new_n15840_ & (\all_features[2530]  | \all_features[2531]  | \all_features[2529] )));
  assign new_n15845_ = ~\all_features[2533]  & \all_features[2534]  & \all_features[2535]  & (\all_features[2532]  ? new_n15843_ : (new_n15839_ | ~new_n15843_));
  assign new_n15846_ = \all_features[2535]  & (\all_features[2533]  | \all_features[2534]  | \all_features[2532] );
  assign new_n15847_ = new_n15848_ & (~\all_features[2533]  | (~\all_features[2532]  & (~\all_features[2531]  | (~\all_features[2530]  & ~\all_features[2529] ))));
  assign new_n15848_ = ~\all_features[2534]  & ~\all_features[2535] ;
  assign new_n15849_ = ~\all_features[2533]  & new_n15848_ & ((~\all_features[2530]  & new_n15842_) | ~\all_features[2532]  | ~\all_features[2531] );
  assign new_n15850_ = ~\all_features[2535]  & (~\all_features[2534]  | (~\all_features[2533]  & (new_n15842_ | ~new_n15838_ | ~\all_features[2532] )));
  assign new_n15851_ = new_n15848_ & (~\all_features[2531]  | ~new_n15840_ | (~\all_features[2530]  & ~new_n15839_));
  assign new_n15852_ = ~\all_features[2535]  & (~\all_features[2534]  | (~\all_features[2532]  & ~\all_features[2533]  & ~new_n15838_));
  assign new_n15853_ = new_n15858_ & (~new_n15859_ | (~new_n15854_ & ~new_n15850_ & ~new_n15852_));
  assign new_n15854_ = ~new_n15835_ & ~new_n15837_ & (~new_n15846_ | ~new_n15841_ | new_n15855_);
  assign new_n15855_ = new_n15844_ & new_n15856_ & (new_n15857_ | ~\all_features[2533]  | ~\all_features[2534]  | ~\all_features[2535] );
  assign new_n15856_ = \all_features[2534]  & \all_features[2535]  & (\all_features[2532]  | \all_features[2533]  | new_n15839_ | ~new_n15843_);
  assign new_n15857_ = ~\all_features[2531]  & ~\all_features[2532]  & (~\all_features[2530]  | new_n15842_);
  assign new_n15858_ = ~new_n15849_ & (\all_features[2531]  | \all_features[2532]  | \all_features[2533]  | \all_features[2534]  | \all_features[2535] );
  assign new_n15859_ = ~new_n15847_ & ~new_n15851_;
  assign new_n15860_ = new_n15861_ & new_n15858_ & ~new_n15851_ & ~new_n15850_ & ~new_n15835_ & ~new_n15847_;
  assign new_n15861_ = ~new_n15837_ & ~new_n15852_;
  assign new_n15862_ = new_n15858_ & new_n15859_ & (new_n15863_ | new_n15835_ | new_n15850_ | ~new_n15861_);
  assign new_n15863_ = new_n15846_ & new_n15856_ & new_n15841_ & new_n15844_;
  assign new_n15864_ = ~new_n11267_ & ~new_n11269_;
  assign new_n15865_ = ~new_n15829_ & (new_n15830_ | ((new_n10645_ | ~new_n15874_ | new_n11622_) & (new_n15866_ | ~new_n11622_)));
  assign new_n15866_ = new_n15873_ ? new_n13318_ : new_n15867_;
  assign new_n15867_ = new_n8929_ & new_n15868_;
  assign new_n15868_ = ~new_n8957_ & ~new_n15869_;
  assign new_n15869_ = ~new_n8950_ & (new_n8949_ | new_n15870_);
  assign new_n15870_ = ~new_n8945_ & (new_n8947_ | (~new_n8940_ & (new_n8941_ | (~new_n8933_ & ~new_n15871_))));
  assign new_n15871_ = ~new_n8935_ & (~new_n8955_ | (new_n8954_ & (~new_n8951_ | (~new_n15872_ & new_n8952_))));
  assign new_n15872_ = \all_features[1198]  & \all_features[1199]  & (\all_features[1197]  | (~new_n8953_ & \all_features[1196] ));
  assign new_n15873_ = new_n6605_ & new_n6627_;
  assign new_n15874_ = new_n15906_ & new_n15904_ & new_n15875_ & new_n15895_;
  assign new_n15875_ = ~new_n15894_ & (new_n15889_ | (~new_n15891_ & (new_n15892_ | (~new_n15876_ & ~new_n15893_))));
  assign new_n15876_ = ~new_n15883_ & (new_n15885_ | (~new_n15887_ & (~new_n15888_ | new_n15877_)));
  assign new_n15877_ = \all_features[1239]  & ((~new_n15882_ & ~\all_features[1237]  & \all_features[1238] ) | (~new_n15880_ & (\all_features[1238]  | (~new_n15878_ & \all_features[1237] ))));
  assign new_n15878_ = new_n15879_ & ~\all_features[1236]  & ~\all_features[1234]  & ~\all_features[1235] ;
  assign new_n15879_ = ~\all_features[1232]  & ~\all_features[1233] ;
  assign new_n15880_ = \all_features[1239]  & (\all_features[1238]  | (new_n15881_ & (\all_features[1234]  | \all_features[1235]  | \all_features[1233] )));
  assign new_n15881_ = \all_features[1236]  & \all_features[1237] ;
  assign new_n15882_ = (~\all_features[1234]  & ~\all_features[1235]  & ~\all_features[1236]  & (~\all_features[1233]  | ~\all_features[1232] )) | (\all_features[1236]  & (\all_features[1234]  | \all_features[1235] ));
  assign new_n15883_ = ~\all_features[1239]  & (~\all_features[1238]  | (~\all_features[1237]  & (new_n15879_ | ~new_n15884_ | ~\all_features[1236] )));
  assign new_n15884_ = \all_features[1234]  & \all_features[1235] ;
  assign new_n15885_ = ~new_n15886_ & ~\all_features[1239] ;
  assign new_n15886_ = \all_features[1237]  & \all_features[1238]  & (\all_features[1236]  | (\all_features[1234]  & \all_features[1235]  & \all_features[1233] ));
  assign new_n15887_ = ~\all_features[1239]  & (~new_n15884_ | ~\all_features[1232]  | ~\all_features[1233]  | ~\all_features[1238]  | ~new_n15881_);
  assign new_n15888_ = \all_features[1239]  & (\all_features[1237]  | \all_features[1238]  | \all_features[1236] );
  assign new_n15889_ = ~\all_features[1237]  & new_n15890_ & ((~\all_features[1234]  & new_n15879_) | ~\all_features[1236]  | ~\all_features[1235] );
  assign new_n15890_ = ~\all_features[1238]  & ~\all_features[1239] ;
  assign new_n15891_ = new_n15890_ & (~\all_features[1237]  | (~\all_features[1236]  & (~\all_features[1235]  | (~\all_features[1234]  & ~\all_features[1233] ))));
  assign new_n15892_ = new_n15890_ & (~new_n15881_ | ~\all_features[1235]  | (~\all_features[1234]  & (~\all_features[1232]  | ~\all_features[1233] )));
  assign new_n15893_ = ~\all_features[1239]  & (~\all_features[1238]  | (~\all_features[1236]  & ~\all_features[1237]  & ~new_n15884_));
  assign new_n15894_ = ~\all_features[1239]  & ~\all_features[1238]  & ~\all_features[1237]  & ~\all_features[1235]  & ~\all_features[1236] ;
  assign new_n15895_ = new_n15901_ & (~new_n15902_ | (new_n15903_ & (new_n15896_ | new_n15885_ | new_n15887_)));
  assign new_n15896_ = new_n15897_ & (~new_n15898_ | (~new_n15900_ & \all_features[1237]  & \all_features[1238]  & \all_features[1239] ));
  assign new_n15897_ = \all_features[1239]  & (\all_features[1238]  | (~new_n15878_ & \all_features[1237] ));
  assign new_n15898_ = \all_features[1239]  & \all_features[1238]  & ~new_n15899_ & new_n15880_;
  assign new_n15899_ = ~\all_features[1234]  & ~\all_features[1235]  & ~\all_features[1236]  & ~\all_features[1237]  & (~\all_features[1233]  | ~\all_features[1232] );
  assign new_n15900_ = ~\all_features[1235]  & ~\all_features[1236]  & (~\all_features[1234]  | new_n15879_);
  assign new_n15901_ = ~new_n15889_ & ~new_n15894_;
  assign new_n15902_ = ~new_n15891_ & ~new_n15892_;
  assign new_n15903_ = ~new_n15893_ & ~new_n15883_;
  assign new_n15904_ = new_n15902_ & ~new_n15905_ & new_n15901_;
  assign new_n15905_ = ~new_n15893_ & ~new_n15883_ & ~new_n15885_ & ~new_n15887_ & (~new_n15898_ | ~new_n15897_);
  assign new_n15906_ = new_n15903_ & new_n15902_ & ~new_n15894_ & ~new_n15887_ & ~new_n15889_ & ~new_n15885_;
  assign new_n15907_ = new_n15404_ & new_n15541_;
  assign new_n15908_ = new_n16059_ & (~new_n14124_ | ~new_n15917_ | ~new_n15909_ | ~new_n15912_);
  assign new_n15909_ = new_n15910_ & (~new_n16024_ | (~new_n16026_ & new_n16025_) | (~new_n16028_ & ~new_n16025_));
  assign new_n15910_ = ~new_n15911_ & new_n15955_ & (~new_n15954_ | (~new_n15919_ & new_n15991_));
  assign new_n15911_ = new_n15912_ & (new_n14124_ ? ~new_n15917_ : ~new_n15918_);
  assign new_n15912_ = new_n15913_ & new_n15915_;
  assign new_n15913_ = ~new_n15914_ & ~new_n9867_;
  assign new_n15914_ = new_n9836_ & new_n9864_;
  assign new_n15915_ = ~new_n11094_ & new_n15916_;
  assign new_n15916_ = ~new_n11083_ & ~new_n11092_;
  assign new_n15917_ = ~new_n7798_ & (~new_n7772_ | ~new_n7799_);
  assign new_n15918_ = ~new_n15587_ & ~new_n15584_;
  assign new_n15919_ = new_n15920_ & new_n15953_;
  assign new_n15920_ = new_n15921_ & new_n15951_;
  assign new_n15921_ = new_n15922_ & new_n15942_;
  assign new_n15922_ = ~new_n15941_ & (new_n15940_ | (~new_n15939_ & (new_n15937_ | (~new_n15936_ & ~new_n15923_))));
  assign new_n15923_ = ~new_n15930_ & (new_n15932_ | (~new_n15934_ & (~new_n15935_ | new_n15924_)));
  assign new_n15924_ = \all_features[5295]  & ((~new_n15929_ & ~\all_features[5293]  & \all_features[5294] ) | (~new_n15927_ & (\all_features[5294]  | (~new_n15925_ & \all_features[5293] ))));
  assign new_n15925_ = new_n15926_ & ~\all_features[5292]  & ~\all_features[5290]  & ~\all_features[5291] ;
  assign new_n15926_ = ~\all_features[5288]  & ~\all_features[5289] ;
  assign new_n15927_ = \all_features[5295]  & (\all_features[5294]  | (new_n15928_ & (\all_features[5290]  | \all_features[5291]  | \all_features[5289] )));
  assign new_n15928_ = \all_features[5292]  & \all_features[5293] ;
  assign new_n15929_ = (~\all_features[5290]  & ~\all_features[5291]  & ~\all_features[5292]  & (~\all_features[5289]  | ~\all_features[5288] )) | (\all_features[5292]  & (\all_features[5290]  | \all_features[5291] ));
  assign new_n15930_ = ~\all_features[5295]  & (~\all_features[5294]  | (~\all_features[5293]  & (new_n15926_ | ~\all_features[5292]  | ~new_n15931_)));
  assign new_n15931_ = \all_features[5290]  & \all_features[5291] ;
  assign new_n15932_ = ~new_n15933_ & ~\all_features[5295] ;
  assign new_n15933_ = \all_features[5293]  & \all_features[5294]  & (\all_features[5292]  | (\all_features[5290]  & \all_features[5291]  & \all_features[5289] ));
  assign new_n15934_ = ~\all_features[5295]  & (~new_n15928_ | ~\all_features[5288]  | ~\all_features[5289]  | ~\all_features[5294]  | ~new_n15931_);
  assign new_n15935_ = \all_features[5295]  & (\all_features[5293]  | \all_features[5294]  | \all_features[5292] );
  assign new_n15936_ = ~\all_features[5295]  & (~\all_features[5294]  | (~\all_features[5292]  & ~\all_features[5293]  & ~new_n15931_));
  assign new_n15937_ = new_n15938_ & (~new_n15928_ | ~\all_features[5291]  | (~\all_features[5290]  & (~\all_features[5288]  | ~\all_features[5289] )));
  assign new_n15938_ = ~\all_features[5294]  & ~\all_features[5295] ;
  assign new_n15939_ = new_n15938_ & (~\all_features[5293]  | (~\all_features[5292]  & (~\all_features[5291]  | (~\all_features[5290]  & ~\all_features[5289] ))));
  assign new_n15940_ = ~\all_features[5293]  & new_n15938_ & ((~\all_features[5290]  & new_n15926_) | ~\all_features[5292]  | ~\all_features[5291] );
  assign new_n15941_ = ~\all_features[5295]  & ~\all_features[5294]  & ~\all_features[5293]  & ~\all_features[5291]  & ~\all_features[5292] ;
  assign new_n15942_ = new_n15950_ & (~new_n15949_ | (new_n15948_ & (new_n15943_ | new_n15932_ | new_n15934_)));
  assign new_n15943_ = new_n15944_ & (~new_n15945_ | (~new_n15947_ & \all_features[5293]  & \all_features[5294]  & \all_features[5295] ));
  assign new_n15944_ = \all_features[5295]  & (\all_features[5294]  | (~new_n15925_ & \all_features[5293] ));
  assign new_n15945_ = \all_features[5295]  & \all_features[5294]  & ~new_n15946_ & new_n15927_;
  assign new_n15946_ = ~\all_features[5290]  & ~\all_features[5291]  & ~\all_features[5292]  & ~\all_features[5293]  & (~\all_features[5289]  | ~\all_features[5288] );
  assign new_n15947_ = ~\all_features[5291]  & ~\all_features[5292]  & (~\all_features[5290]  | new_n15926_);
  assign new_n15948_ = ~new_n15930_ & ~new_n15936_;
  assign new_n15949_ = ~new_n15937_ & ~new_n15939_;
  assign new_n15950_ = ~new_n15940_ & ~new_n15941_;
  assign new_n15951_ = new_n15950_ & ~new_n15952_ & new_n15949_;
  assign new_n15952_ = ~new_n15930_ & ~new_n15936_ & ~new_n15932_ & ~new_n15934_ & (~new_n15945_ | ~new_n15944_);
  assign new_n15953_ = new_n15949_ & new_n15948_ & new_n15950_ & ~new_n15932_ & ~new_n15934_;
  assign new_n15954_ = ~new_n15913_ & new_n12152_;
  assign new_n15955_ = ~new_n15913_ | ((new_n14124_ | ~new_n15918_ | ~new_n15915_) & (new_n10099_ | ~new_n15956_ | new_n15915_));
  assign new_n15956_ = new_n15990_ & (new_n15986_ | ~new_n15957_);
  assign new_n15957_ = ~new_n15958_ & ~new_n15982_;
  assign new_n15958_ = ~new_n15980_ & ~new_n15979_ & (~new_n15973_ | (~new_n15959_ & ~new_n15977_ & ~new_n15981_));
  assign new_n15959_ = ~new_n15968_ & ~new_n15969_ & (~new_n15972_ | ~new_n15971_ | new_n15960_);
  assign new_n15960_ = new_n15961_ & new_n15963_ & (new_n15966_ | ~\all_features[2341]  | ~\all_features[2342]  | ~\all_features[2343] );
  assign new_n15961_ = \all_features[2343]  & (\all_features[2342]  | (new_n15962_ & (\all_features[2338]  | \all_features[2339]  | \all_features[2337] )));
  assign new_n15962_ = \all_features[2340]  & \all_features[2341] ;
  assign new_n15963_ = \all_features[2342]  & \all_features[2343]  & (\all_features[2340]  | \all_features[2341]  | new_n15964_ | ~new_n15965_);
  assign new_n15964_ = \all_features[2336]  & \all_features[2337] ;
  assign new_n15965_ = ~\all_features[2338]  & ~\all_features[2339] ;
  assign new_n15966_ = ~\all_features[2339]  & ~\all_features[2340]  & (~\all_features[2338]  | new_n15967_);
  assign new_n15967_ = ~\all_features[2336]  & ~\all_features[2337] ;
  assign new_n15968_ = ~\all_features[2343]  & (~new_n15962_ | ~\all_features[2338]  | ~\all_features[2339]  | ~\all_features[2342]  | ~new_n15964_);
  assign new_n15969_ = ~new_n15970_ & ~\all_features[2343] ;
  assign new_n15970_ = \all_features[2341]  & \all_features[2342]  & (\all_features[2340]  | (\all_features[2338]  & \all_features[2339]  & \all_features[2337] ));
  assign new_n15971_ = \all_features[2343]  & (\all_features[2342]  | (\all_features[2341]  & (\all_features[2340]  | ~new_n15965_ | ~new_n15967_)));
  assign new_n15972_ = \all_features[2343]  & (\all_features[2341]  | \all_features[2342]  | \all_features[2340] );
  assign new_n15973_ = ~new_n15974_ & ~new_n15976_;
  assign new_n15974_ = new_n15975_ & (~\all_features[2339]  | ~new_n15962_ | (~\all_features[2338]  & ~new_n15964_));
  assign new_n15975_ = ~\all_features[2342]  & ~\all_features[2343] ;
  assign new_n15976_ = new_n15975_ & (~\all_features[2341]  | (~\all_features[2340]  & (~\all_features[2339]  | (~\all_features[2338]  & ~\all_features[2337] ))));
  assign new_n15977_ = ~\all_features[2343]  & (~\all_features[2342]  | new_n15978_);
  assign new_n15978_ = ~\all_features[2341]  & (new_n15967_ | ~\all_features[2339]  | ~\all_features[2340]  | ~\all_features[2338] );
  assign new_n15979_ = ~\all_features[2341]  & new_n15975_ & ((~\all_features[2338]  & new_n15967_) | ~\all_features[2340]  | ~\all_features[2339] );
  assign new_n15980_ = ~\all_features[2343]  & ~\all_features[2342]  & ~\all_features[2341]  & ~\all_features[2339]  & ~\all_features[2340] ;
  assign new_n15981_ = ~\all_features[2343]  & (~\all_features[2342]  | (~\all_features[2341]  & ~\all_features[2340]  & (~\all_features[2339]  | ~\all_features[2338] )));
  assign new_n15982_ = ~new_n15983_ & ~new_n15980_;
  assign new_n15983_ = ~new_n15979_ & (new_n15976_ | (~new_n15974_ & (new_n15981_ | (~new_n15977_ & ~new_n15984_))));
  assign new_n15984_ = ~new_n15969_ & (new_n15968_ | (new_n15972_ & (~new_n15971_ | (~new_n15985_ & new_n15961_))));
  assign new_n15985_ = ~\all_features[2341]  & \all_features[2342]  & \all_features[2343]  & (\all_features[2340]  ? new_n15965_ : (new_n15964_ | ~new_n15965_));
  assign new_n15986_ = ~new_n15980_ & ~new_n15979_ & ~new_n15976_ & ~new_n15987_ & ~new_n15974_;
  assign new_n15987_ = ~new_n15977_ & ~new_n15968_ & new_n15988_ & (~new_n15971_ | ~new_n15989_);
  assign new_n15988_ = ~new_n15969_ & ~new_n15981_;
  assign new_n15989_ = new_n15972_ & new_n15961_ & new_n15963_;
  assign new_n15990_ = new_n15973_ & new_n15988_ & ~new_n15980_ & ~new_n15968_ & ~new_n15977_ & ~new_n15979_;
  assign new_n15991_ = ~new_n16023_ & new_n15992_;
  assign new_n15992_ = ~new_n15993_ & ~new_n16018_;
  assign new_n15993_ = new_n16015_ & ~new_n15994_ & new_n16011_;
  assign new_n15994_ = new_n16001_ & (~new_n16009_ | ~new_n16010_ | ~new_n15998_ | ~new_n15995_);
  assign new_n15995_ = \all_features[4663]  & (\all_features[4662]  | new_n15996_);
  assign new_n15996_ = \all_features[4661]  & (\all_features[4658]  | \all_features[4659]  | \all_features[4660]  | ~new_n15997_);
  assign new_n15997_ = ~\all_features[4656]  & ~\all_features[4657] ;
  assign new_n15998_ = \all_features[4663]  & ~new_n15999_ & \all_features[4662] ;
  assign new_n15999_ = ~\all_features[4661]  & ~\all_features[4660]  & ~\all_features[4659]  & ~new_n16000_ & ~\all_features[4658] ;
  assign new_n16000_ = \all_features[4656]  & \all_features[4657] ;
  assign new_n16001_ = ~new_n16007_ & ~new_n16005_ & ~new_n16002_ & ~new_n16004_;
  assign new_n16002_ = ~\all_features[4663]  & (~\all_features[4662]  | (~\all_features[4660]  & ~\all_features[4661]  & ~new_n16003_));
  assign new_n16003_ = \all_features[4658]  & \all_features[4659] ;
  assign new_n16004_ = ~\all_features[4663]  & (~\all_features[4662]  | (~\all_features[4661]  & (new_n15997_ | ~\all_features[4660]  | ~new_n16003_)));
  assign new_n16005_ = ~new_n16006_ & ~\all_features[4663] ;
  assign new_n16006_ = \all_features[4661]  & \all_features[4662]  & (\all_features[4660]  | (\all_features[4658]  & \all_features[4659]  & \all_features[4657] ));
  assign new_n16007_ = ~\all_features[4663]  & (~\all_features[4662]  | ~new_n16003_ | ~new_n16000_ | ~new_n16008_);
  assign new_n16008_ = \all_features[4660]  & \all_features[4661] ;
  assign new_n16009_ = \all_features[4663]  & (\all_features[4662]  | (new_n16008_ & (\all_features[4658]  | \all_features[4659]  | \all_features[4657] )));
  assign new_n16010_ = \all_features[4663]  & (\all_features[4661]  | \all_features[4662]  | \all_features[4660] );
  assign new_n16011_ = ~new_n16012_ & ~new_n16014_;
  assign new_n16012_ = new_n16013_ & (~\all_features[4659]  | ~new_n16008_ | (~\all_features[4658]  & ~new_n16000_));
  assign new_n16013_ = ~\all_features[4662]  & ~\all_features[4663] ;
  assign new_n16014_ = new_n16013_ & (~\all_features[4661]  | (~\all_features[4660]  & (~\all_features[4659]  | (~\all_features[4658]  & ~\all_features[4657] ))));
  assign new_n16015_ = ~new_n16016_ & ~new_n16017_;
  assign new_n16016_ = ~\all_features[4661]  & new_n16013_ & ((~\all_features[4658]  & new_n15997_) | ~\all_features[4660]  | ~\all_features[4659] );
  assign new_n16017_ = ~\all_features[4663]  & ~\all_features[4662]  & ~\all_features[4661]  & ~\all_features[4659]  & ~\all_features[4660] ;
  assign new_n16018_ = new_n16015_ & (~new_n16011_ | (new_n16022_ & (new_n16019_ | new_n16005_ | new_n16007_)));
  assign new_n16019_ = new_n16010_ & ~new_n16020_ & new_n15995_;
  assign new_n16020_ = ~new_n15999_ & new_n16009_ & \all_features[4662]  & \all_features[4663]  & (~\all_features[4661]  | new_n16021_);
  assign new_n16021_ = ~\all_features[4659]  & ~\all_features[4660]  & (~\all_features[4658]  | new_n15997_);
  assign new_n16022_ = ~new_n16002_ & ~new_n16004_;
  assign new_n16023_ = new_n16011_ & new_n16022_ & ~new_n16017_ & ~new_n16007_ & ~new_n16005_ & ~new_n16016_;
  assign new_n16024_ = ~new_n15913_ & ~new_n12152_;
  assign new_n16025_ = new_n15587_ & (new_n15584_ | new_n15555_);
  assign new_n16026_ = new_n16027_ & ~new_n15743_ & ~new_n15745_;
  assign new_n16027_ = ~new_n15717_ & ~new_n15747_;
  assign new_n16028_ = new_n16029_ & new_n16058_;
  assign new_n16029_ = new_n16030_ & new_n16054_;
  assign new_n16030_ = new_n16031_ & (~new_n16045_ | (new_n16041_ & new_n16052_ & new_n16053_));
  assign new_n16031_ = new_n16032_ & ~new_n16037_ & ~new_n16038_;
  assign new_n16032_ = ~new_n16033_ & ~new_n16036_;
  assign new_n16033_ = ~\all_features[2549]  & new_n16035_ & ((~\all_features[2546]  & new_n16034_) | ~\all_features[2548]  | ~\all_features[2547] );
  assign new_n16034_ = ~\all_features[2544]  & ~\all_features[2545] ;
  assign new_n16035_ = ~\all_features[2550]  & ~\all_features[2551] ;
  assign new_n16036_ = ~\all_features[2551]  & ~\all_features[2550]  & ~\all_features[2549]  & ~\all_features[2547]  & ~\all_features[2548] ;
  assign new_n16037_ = new_n16035_ & (~\all_features[2549]  | (~\all_features[2548]  & (~\all_features[2547]  | (~\all_features[2546]  & ~\all_features[2545] ))));
  assign new_n16038_ = new_n16035_ & (~\all_features[2547]  | ~new_n16040_ | (~\all_features[2546]  & ~new_n16039_));
  assign new_n16039_ = \all_features[2544]  & \all_features[2545] ;
  assign new_n16040_ = \all_features[2548]  & \all_features[2549] ;
  assign new_n16041_ = new_n16042_ & new_n16044_;
  assign new_n16042_ = \all_features[2551]  & (\all_features[2550]  | (\all_features[2549]  & (\all_features[2548]  | ~new_n16034_ | ~new_n16043_)));
  assign new_n16043_ = ~\all_features[2546]  & ~\all_features[2547] ;
  assign new_n16044_ = \all_features[2551]  & (\all_features[2549]  | \all_features[2550]  | \all_features[2548] );
  assign new_n16045_ = ~new_n16051_ & ~new_n16050_ & ~new_n16046_ & ~new_n16048_;
  assign new_n16046_ = ~\all_features[2551]  & (~\all_features[2550]  | (~\all_features[2549]  & (new_n16034_ | ~new_n16047_ | ~\all_features[2548] )));
  assign new_n16047_ = \all_features[2546]  & \all_features[2547] ;
  assign new_n16048_ = ~new_n16049_ & ~\all_features[2551] ;
  assign new_n16049_ = \all_features[2549]  & \all_features[2550]  & (\all_features[2548]  | (\all_features[2546]  & \all_features[2547]  & \all_features[2545] ));
  assign new_n16050_ = ~\all_features[2551]  & (~\all_features[2550]  | ~new_n16039_ | ~new_n16040_ | ~new_n16047_);
  assign new_n16051_ = ~\all_features[2551]  & (~\all_features[2550]  | (~\all_features[2548]  & ~\all_features[2549]  & ~new_n16047_));
  assign new_n16052_ = \all_features[2550]  & \all_features[2551]  & (\all_features[2548]  | \all_features[2549]  | new_n16039_ | ~new_n16043_);
  assign new_n16053_ = \all_features[2551]  & (\all_features[2550]  | (new_n16040_ & (\all_features[2546]  | \all_features[2547]  | \all_features[2545] )));
  assign new_n16054_ = new_n16032_ & (new_n16038_ | new_n16037_ | (~new_n16046_ & ~new_n16051_ & ~new_n16055_));
  assign new_n16055_ = ~new_n16048_ & ~new_n16050_ & (~new_n16041_ | (~new_n16056_ & new_n16052_ & new_n16053_));
  assign new_n16056_ = \all_features[2551]  & \all_features[2550]  & ~new_n16057_ & \all_features[2549] ;
  assign new_n16057_ = ~\all_features[2547]  & ~\all_features[2548]  & (~\all_features[2546]  | new_n16034_);
  assign new_n16058_ = new_n16031_ & new_n16045_;
  assign new_n16059_ = ~new_n16061_ & ~new_n16060_ & (~new_n15991_ | ~new_n15954_ | new_n15919_);
  assign new_n16060_ = new_n16024_ & (new_n16025_ ? ~new_n16026_ : ~new_n16028_);
  assign new_n16061_ = ~new_n15915_ & new_n15913_ & (new_n10099_ ? ~new_n8697_ : ~new_n15956_);
  assign new_n16062_ = new_n16107_ & (new_n16104_ ? (new_n16142_ ? ~new_n16148_ : new_n14654_) : new_n16063_);
  assign new_n16063_ = ~new_n16102_ & new_n16064_;
  assign new_n16064_ = new_n16065_ & new_n16097_;
  assign new_n16065_ = new_n16066_ & (new_n16080_ | (~new_n16083_ & (new_n16084_ | new_n16093_)));
  assign new_n16066_ = new_n16067_ & (\all_features[4363]  | \all_features[4364]  | \all_features[4365]  | \all_features[4366]  | \all_features[4367] );
  assign new_n16067_ = new_n16079_ & (~new_n16082_ | (new_n16085_ & (~new_n16089_ | new_n16068_)));
  assign new_n16068_ = new_n16069_ & (~new_n16073_ | (~new_n16078_ & \all_features[4365]  & \all_features[4366]  & \all_features[4367] ));
  assign new_n16069_ = \all_features[4367]  & (\all_features[4366]  | (~new_n16070_ & \all_features[4365] ));
  assign new_n16070_ = new_n16071_ & ~\all_features[4364]  & new_n16072_;
  assign new_n16071_ = ~\all_features[4360]  & ~\all_features[4361] ;
  assign new_n16072_ = ~\all_features[4362]  & ~\all_features[4363] ;
  assign new_n16073_ = \all_features[4367]  & \all_features[4366]  & ~new_n16076_ & new_n16074_;
  assign new_n16074_ = \all_features[4367]  & (\all_features[4366]  | (new_n16075_ & (\all_features[4362]  | \all_features[4363]  | \all_features[4361] )));
  assign new_n16075_ = \all_features[4364]  & \all_features[4365] ;
  assign new_n16076_ = new_n16072_ & ~\all_features[4365]  & ~new_n16077_ & ~\all_features[4364] ;
  assign new_n16077_ = \all_features[4360]  & \all_features[4361] ;
  assign new_n16078_ = ~\all_features[4363]  & ~\all_features[4364]  & (~\all_features[4362]  | new_n16071_);
  assign new_n16079_ = ~new_n16080_ & (\all_features[4363]  | \all_features[4364]  | \all_features[4365]  | \all_features[4366]  | \all_features[4367] );
  assign new_n16080_ = ~\all_features[4365]  & new_n16081_ & ((~\all_features[4362]  & new_n16071_) | ~\all_features[4364]  | ~\all_features[4363] );
  assign new_n16081_ = ~\all_features[4366]  & ~\all_features[4367] ;
  assign new_n16082_ = ~new_n16083_ & ~new_n16084_;
  assign new_n16083_ = new_n16081_ & (~\all_features[4365]  | (~\all_features[4364]  & (~\all_features[4363]  | (~\all_features[4362]  & ~\all_features[4361] ))));
  assign new_n16084_ = new_n16081_ & (~\all_features[4363]  | ~new_n16075_ | (~\all_features[4362]  & ~new_n16077_));
  assign new_n16085_ = ~new_n16086_ & ~new_n16088_;
  assign new_n16086_ = ~\all_features[4367]  & (~\all_features[4366]  | (~\all_features[4364]  & ~\all_features[4365]  & ~new_n16087_));
  assign new_n16087_ = \all_features[4362]  & \all_features[4363] ;
  assign new_n16088_ = ~\all_features[4367]  & (~\all_features[4366]  | (~\all_features[4365]  & (new_n16071_ | ~new_n16087_ | ~\all_features[4364] )));
  assign new_n16089_ = ~new_n16090_ & ~new_n16092_;
  assign new_n16090_ = ~new_n16091_ & ~\all_features[4367] ;
  assign new_n16091_ = \all_features[4365]  & \all_features[4366]  & (\all_features[4364]  | (\all_features[4362]  & \all_features[4363]  & \all_features[4361] ));
  assign new_n16092_ = ~\all_features[4367]  & (~\all_features[4366]  | ~new_n16077_ | ~new_n16075_ | ~new_n16087_);
  assign new_n16093_ = ~new_n16086_ & (new_n16088_ | (~new_n16090_ & (new_n16092_ | (~new_n16094_ & new_n16096_))));
  assign new_n16094_ = \all_features[4367]  & ((~new_n16095_ & ~\all_features[4365]  & \all_features[4366] ) | (~new_n16074_ & (\all_features[4366]  | (~new_n16070_ & \all_features[4365] ))));
  assign new_n16095_ = (\all_features[4364]  & ~new_n16072_) | (~new_n16077_ & ~\all_features[4364]  & new_n16072_);
  assign new_n16096_ = \all_features[4367]  & (\all_features[4365]  | \all_features[4366]  | \all_features[4364] );
  assign new_n16097_ = new_n16098_ & new_n16101_;
  assign new_n16098_ = new_n16099_ & (new_n16088_ | new_n16090_ | ~new_n16100_ | (new_n16073_ & new_n16069_));
  assign new_n16099_ = new_n16079_ & new_n16082_;
  assign new_n16100_ = ~new_n16086_ & ~new_n16092_;
  assign new_n16101_ = new_n16089_ & new_n16099_ & new_n16085_;
  assign new_n16102_ = new_n15408_ & new_n16103_;
  assign new_n16103_ = ~new_n15437_ & ~new_n15441_;
  assign new_n16104_ = ~new_n16105_ & new_n16106_;
  assign new_n16105_ = new_n15832_ & new_n15853_;
  assign new_n16106_ = ~new_n15860_ & ~new_n15862_;
  assign new_n16107_ = ~new_n16140_ & (~new_n16136_ | ~new_n16108_);
  assign new_n16108_ = new_n16109_ & new_n16133_;
  assign new_n16109_ = new_n16130_ & (~new_n16124_ | (~new_n16110_ & ~new_n16128_ & ~new_n16132_));
  assign new_n16110_ = ~new_n16119_ & ~new_n16120_ & (~new_n16123_ | ~new_n16122_ | new_n16111_);
  assign new_n16111_ = new_n16112_ & new_n16114_ & (new_n16117_ | ~\all_features[4453]  | ~\all_features[4454]  | ~\all_features[4455] );
  assign new_n16112_ = \all_features[4455]  & (\all_features[4454]  | (new_n16113_ & (\all_features[4450]  | \all_features[4451]  | \all_features[4449] )));
  assign new_n16113_ = \all_features[4452]  & \all_features[4453] ;
  assign new_n16114_ = \all_features[4454]  & \all_features[4455]  & (\all_features[4452]  | \all_features[4453]  | new_n16115_ | ~new_n16116_);
  assign new_n16115_ = \all_features[4448]  & \all_features[4449] ;
  assign new_n16116_ = ~\all_features[4450]  & ~\all_features[4451] ;
  assign new_n16117_ = ~\all_features[4451]  & ~\all_features[4452]  & (~\all_features[4450]  | new_n16118_);
  assign new_n16118_ = ~\all_features[4448]  & ~\all_features[4449] ;
  assign new_n16119_ = ~\all_features[4455]  & (~new_n16113_ | ~\all_features[4450]  | ~\all_features[4451]  | ~\all_features[4454]  | ~new_n16115_);
  assign new_n16120_ = ~new_n16121_ & ~\all_features[4455] ;
  assign new_n16121_ = \all_features[4453]  & \all_features[4454]  & (\all_features[4452]  | (\all_features[4450]  & \all_features[4451]  & \all_features[4449] ));
  assign new_n16122_ = \all_features[4455]  & (\all_features[4454]  | (\all_features[4453]  & (\all_features[4452]  | ~new_n16116_ | ~new_n16118_)));
  assign new_n16123_ = \all_features[4455]  & (\all_features[4453]  | \all_features[4454]  | \all_features[4452] );
  assign new_n16124_ = ~new_n16125_ & ~new_n16127_;
  assign new_n16125_ = new_n16126_ & (~\all_features[4451]  | ~new_n16113_ | (~\all_features[4450]  & ~new_n16115_));
  assign new_n16126_ = ~\all_features[4454]  & ~\all_features[4455] ;
  assign new_n16127_ = new_n16126_ & (~\all_features[4453]  | (~\all_features[4452]  & (~\all_features[4451]  | (~\all_features[4450]  & ~\all_features[4449] ))));
  assign new_n16128_ = ~\all_features[4455]  & (~\all_features[4454]  | new_n16129_);
  assign new_n16129_ = ~\all_features[4453]  & (new_n16118_ | ~\all_features[4451]  | ~\all_features[4452]  | ~\all_features[4450] );
  assign new_n16130_ = ~new_n16131_ & (\all_features[4451]  | \all_features[4452]  | \all_features[4453]  | \all_features[4454]  | \all_features[4455] );
  assign new_n16131_ = ~\all_features[4453]  & new_n16126_ & ((~\all_features[4450]  & new_n16118_) | ~\all_features[4452]  | ~\all_features[4451] );
  assign new_n16132_ = ~\all_features[4455]  & (~\all_features[4454]  | (~\all_features[4453]  & ~\all_features[4452]  & (~\all_features[4451]  | ~\all_features[4450] )));
  assign new_n16133_ = new_n16124_ & new_n16130_ & (new_n16128_ | new_n16135_ | new_n16119_ | ~new_n16134_);
  assign new_n16134_ = ~new_n16120_ & ~new_n16132_;
  assign new_n16135_ = new_n16123_ & new_n16114_ & new_n16122_ & new_n16112_;
  assign new_n16136_ = ~new_n16137_ & (\all_features[4451]  | \all_features[4452]  | \all_features[4453]  | \all_features[4454]  | \all_features[4455] );
  assign new_n16137_ = ~new_n16131_ & (new_n16127_ | (~new_n16125_ & (new_n16132_ | (~new_n16128_ & ~new_n16138_))));
  assign new_n16138_ = ~new_n16120_ & (new_n16119_ | (new_n16123_ & (~new_n16122_ | (~new_n16139_ & new_n16112_))));
  assign new_n16139_ = ~\all_features[4453]  & \all_features[4454]  & \all_features[4455]  & (\all_features[4452]  ? new_n16116_ : (new_n16115_ | ~new_n16116_));
  assign new_n16140_ = new_n16141_ & new_n16134_ & new_n16124_ & ~new_n16128_ & ~new_n16131_;
  assign new_n16141_ = ~new_n16119_ & (\all_features[4451]  | \all_features[4452]  | \all_features[4453]  | \all_features[4454]  | \all_features[4455] );
  assign new_n16142_ = new_n15628_ & (new_n15600_ | new_n16143_);
  assign new_n16143_ = new_n15623_ & new_n16144_;
  assign new_n16144_ = ~new_n16145_ & ~new_n15622_;
  assign new_n16145_ = ~new_n15621_ & (new_n15620_ | (~new_n15618_ & (new_n15608_ | (~new_n15602_ & ~new_n16146_))));
  assign new_n16146_ = ~new_n15606_ & (new_n15616_ | (new_n15615_ & (~new_n15617_ | (~new_n16147_ & new_n15610_))));
  assign new_n16147_ = ~\all_features[5069]  & \all_features[5070]  & \all_features[5071]  & (\all_features[5068]  ? new_n15614_ : (new_n15613_ | ~new_n15614_));
  assign new_n16148_ = new_n10677_ & (new_n10679_ | ~new_n10648_);
  assign new_n16149_ = new_n16320_ & (new_n16323_ | ~new_n16150_);
  assign new_n16150_ = new_n16151_ & ((new_n16281_ & new_n10489_) | ~new_n16319_ | new_n16280_);
  assign new_n16151_ = new_n16152_ & (~new_n16278_ | ~new_n16265_) & (~new_n16275_ | ~new_n16266_);
  assign new_n16152_ = (~new_n16153_ | new_n16264_) & (~new_n16229_ | (new_n16232_ ? ~new_n16233_ : ~new_n16230_));
  assign new_n16153_ = new_n16154_ & new_n16227_;
  assign new_n16154_ = ~new_n16155_ & ~new_n16192_;
  assign new_n16155_ = new_n16190_ & new_n16156_ & new_n16188_;
  assign new_n16156_ = new_n16157_ & (new_n16183_ | new_n16184_);
  assign new_n16157_ = new_n16158_ & (\all_features[4603]  | \all_features[4604]  | \all_features[4605]  | \all_features[4606]  | \all_features[4607] );
  assign new_n16158_ = new_n16182_ & (~new_n16170_ | (new_n16179_ & (~new_n16174_ | new_n16159_)));
  assign new_n16159_ = new_n16169_ & ~new_n16163_ & new_n16160_;
  assign new_n16160_ = \all_features[4607]  & (\all_features[4606]  | new_n16161_);
  assign new_n16161_ = \all_features[4605]  & (\all_features[4602]  | \all_features[4603]  | \all_features[4604]  | ~new_n16162_);
  assign new_n16162_ = ~\all_features[4600]  & ~\all_features[4601] ;
  assign new_n16163_ = ~new_n16166_ & new_n16164_ & \all_features[4606]  & \all_features[4607]  & (~\all_features[4605]  | new_n16168_);
  assign new_n16164_ = \all_features[4607]  & (\all_features[4606]  | (new_n16165_ & (\all_features[4602]  | \all_features[4603]  | \all_features[4601] )));
  assign new_n16165_ = \all_features[4604]  & \all_features[4605] ;
  assign new_n16166_ = ~\all_features[4605]  & ~\all_features[4604]  & ~\all_features[4603]  & ~new_n16167_ & ~\all_features[4602] ;
  assign new_n16167_ = \all_features[4600]  & \all_features[4601] ;
  assign new_n16168_ = ~\all_features[4603]  & ~\all_features[4604]  & (~\all_features[4602]  | new_n16162_);
  assign new_n16169_ = \all_features[4607]  & (\all_features[4605]  | \all_features[4606]  | \all_features[4604] );
  assign new_n16170_ = ~new_n16171_ & ~new_n16173_;
  assign new_n16171_ = new_n16172_ & (~\all_features[4605]  | (~\all_features[4604]  & (~\all_features[4603]  | (~\all_features[4602]  & ~\all_features[4601] ))));
  assign new_n16172_ = ~\all_features[4606]  & ~\all_features[4607] ;
  assign new_n16173_ = new_n16172_ & (~\all_features[4603]  | ~new_n16165_ | (~\all_features[4602]  & ~new_n16167_));
  assign new_n16174_ = ~new_n16175_ & ~new_n16177_;
  assign new_n16175_ = ~new_n16176_ & ~\all_features[4607] ;
  assign new_n16176_ = \all_features[4605]  & \all_features[4606]  & (\all_features[4604]  | (\all_features[4602]  & \all_features[4603]  & \all_features[4601] ));
  assign new_n16177_ = ~\all_features[4607]  & (~\all_features[4606]  | ~new_n16167_ | ~new_n16165_ | ~new_n16178_);
  assign new_n16178_ = \all_features[4602]  & \all_features[4603] ;
  assign new_n16179_ = ~new_n16180_ & ~new_n16181_;
  assign new_n16180_ = ~\all_features[4607]  & (~\all_features[4606]  | (~\all_features[4604]  & ~\all_features[4605]  & ~new_n16178_));
  assign new_n16181_ = ~\all_features[4607]  & (~\all_features[4606]  | (~\all_features[4605]  & (new_n16162_ | ~new_n16178_ | ~\all_features[4604] )));
  assign new_n16182_ = ~new_n16183_ & (\all_features[4603]  | \all_features[4604]  | \all_features[4605]  | \all_features[4606]  | \all_features[4607] );
  assign new_n16183_ = ~\all_features[4605]  & new_n16172_ & ((~\all_features[4602]  & new_n16162_) | ~\all_features[4604]  | ~\all_features[4603] );
  assign new_n16184_ = ~new_n16171_ & (new_n16173_ | (~new_n16180_ & (new_n16181_ | (~new_n16185_ & ~new_n16175_))));
  assign new_n16185_ = ~new_n16177_ & (~new_n16169_ | (new_n16160_ & (~new_n16164_ | (~new_n16187_ & new_n16186_))));
  assign new_n16186_ = \all_features[4607]  & ~new_n16166_ & \all_features[4606] ;
  assign new_n16187_ = \all_features[4606]  & \all_features[4607]  & (\all_features[4605]  | (\all_features[4604]  & (\all_features[4603]  | \all_features[4602] )));
  assign new_n16188_ = new_n16170_ & new_n16182_ & (~new_n16179_ | ~new_n16174_ | (new_n16189_ & new_n16160_));
  assign new_n16189_ = new_n16169_ & new_n16186_ & new_n16164_;
  assign new_n16190_ = new_n16191_ & new_n16170_ & ~new_n16175_ & ~new_n16181_ & ~new_n16183_ & ~new_n16180_;
  assign new_n16191_ = ~new_n16177_ & (\all_features[4603]  | \all_features[4604]  | \all_features[4605]  | \all_features[4606]  | \all_features[4607] );
  assign new_n16192_ = new_n16215_ & ~new_n16193_ & ~new_n16224_;
  assign new_n16193_ = ~new_n16194_ & (\all_features[3939]  | \all_features[3940]  | \all_features[3941]  | \all_features[3942]  | \all_features[3943] );
  assign new_n16194_ = ~new_n16209_ & (new_n16211_ | (~new_n16212_ & (new_n16213_ | (~new_n16195_ & ~new_n16214_))));
  assign new_n16195_ = ~new_n16205_ & (new_n16207_ | new_n16196_);
  assign new_n16196_ = \all_features[3943]  & ((new_n16197_ & (\all_features[3942]  | \all_features[3941] )) | (~\all_features[3942]  & (\all_features[3941]  ? new_n16203_ : \all_features[3940] )));
  assign new_n16197_ = new_n16198_ & (\all_features[3941]  | ~new_n16202_ | (~new_n16200_ & ~\all_features[3940]  & new_n16201_) | (\all_features[3940]  & ~new_n16201_));
  assign new_n16198_ = \all_features[3943]  & (\all_features[3942]  | (new_n16199_ & (\all_features[3938]  | \all_features[3939]  | \all_features[3937] )));
  assign new_n16199_ = \all_features[3940]  & \all_features[3941] ;
  assign new_n16200_ = \all_features[3936]  & \all_features[3937] ;
  assign new_n16201_ = ~\all_features[3938]  & ~\all_features[3939] ;
  assign new_n16202_ = \all_features[3942]  & \all_features[3943] ;
  assign new_n16203_ = new_n16204_ & ~\all_features[3940]  & new_n16201_;
  assign new_n16204_ = ~\all_features[3936]  & ~\all_features[3937] ;
  assign new_n16205_ = ~new_n16206_ & ~\all_features[3943] ;
  assign new_n16206_ = \all_features[3941]  & \all_features[3942]  & (\all_features[3940]  | (\all_features[3938]  & \all_features[3939]  & \all_features[3937] ));
  assign new_n16207_ = ~\all_features[3943]  & (~\all_features[3942]  | ~new_n16200_ | ~new_n16199_ | ~new_n16208_);
  assign new_n16208_ = \all_features[3938]  & \all_features[3939] ;
  assign new_n16209_ = ~\all_features[3941]  & new_n16210_ & ((~\all_features[3938]  & new_n16204_) | ~\all_features[3940]  | ~\all_features[3939] );
  assign new_n16210_ = ~\all_features[3942]  & ~\all_features[3943] ;
  assign new_n16211_ = new_n16210_ & (~\all_features[3941]  | (~\all_features[3940]  & (~\all_features[3939]  | (~\all_features[3938]  & ~\all_features[3937] ))));
  assign new_n16212_ = new_n16210_ & (~\all_features[3939]  | ~new_n16199_ | (~\all_features[3938]  & ~new_n16200_));
  assign new_n16213_ = ~\all_features[3943]  & (~\all_features[3942]  | (~\all_features[3940]  & ~\all_features[3941]  & ~new_n16208_));
  assign new_n16214_ = ~\all_features[3943]  & (~\all_features[3942]  | (~\all_features[3941]  & (new_n16204_ | ~new_n16208_ | ~\all_features[3940] )));
  assign new_n16215_ = ~new_n16216_ & ~new_n16222_;
  assign new_n16216_ = new_n16221_ & ~new_n16212_ & ~new_n16217_ & ~new_n16211_;
  assign new_n16217_ = new_n16219_ & (~new_n16218_ | ~new_n16198_ | ~new_n16220_);
  assign new_n16218_ = \all_features[3943]  & (\all_features[3942]  | (~new_n16203_ & \all_features[3941] ));
  assign new_n16219_ = ~new_n16207_ & ~new_n16205_ & ~new_n16213_ & ~new_n16214_;
  assign new_n16220_ = new_n16202_ & (new_n16200_ | \all_features[3940]  | \all_features[3941]  | ~new_n16201_);
  assign new_n16221_ = ~new_n16209_ & (\all_features[3939]  | \all_features[3940]  | \all_features[3941]  | \all_features[3942]  | \all_features[3943] );
  assign new_n16222_ = new_n16223_ & new_n16221_ & ~new_n16211_ & ~new_n16205_;
  assign new_n16223_ = ~new_n16207_ & ~new_n16214_ & ~new_n16212_ & ~new_n16213_;
  assign new_n16224_ = new_n16221_ & (new_n16212_ | new_n16211_ | (~new_n16225_ & ~new_n16213_ & ~new_n16214_));
  assign new_n16225_ = ~new_n16207_ & ~new_n16205_ & (~new_n16218_ | (~new_n16226_ & new_n16198_ & new_n16220_));
  assign new_n16226_ = new_n16202_ & \all_features[3941]  & ((~new_n16204_ & \all_features[3938] ) | \all_features[3940]  | \all_features[3939] );
  assign new_n16227_ = new_n16228_ & new_n8768_;
  assign new_n16228_ = new_n8743_ & new_n8765_;
  assign new_n16229_ = ~new_n16155_ & new_n16192_;
  assign new_n16230_ = new_n16231_ & new_n9018_;
  assign new_n16231_ = new_n9023_ & new_n8993_;
  assign new_n16232_ = ~new_n14834_ & new_n15589_;
  assign new_n16233_ = ~new_n16263_ & new_n16234_;
  assign new_n16234_ = ~new_n16235_ & ~new_n16261_;
  assign new_n16235_ = new_n16255_ & (~new_n16251_ | (new_n16247_ & (new_n16236_ | new_n16258_ | new_n16260_)));
  assign new_n16236_ = new_n16237_ & (~new_n16241_ | (~new_n16246_ & \all_features[2773]  & \all_features[2774]  & \all_features[2775] ));
  assign new_n16237_ = \all_features[2775]  & (\all_features[2774]  | (~new_n16238_ & \all_features[2773] ));
  assign new_n16238_ = new_n16239_ & ~\all_features[2772]  & new_n16240_;
  assign new_n16239_ = ~\all_features[2768]  & ~\all_features[2769] ;
  assign new_n16240_ = ~\all_features[2770]  & ~\all_features[2771] ;
  assign new_n16241_ = \all_features[2775]  & \all_features[2774]  & ~new_n16244_ & new_n16242_;
  assign new_n16242_ = \all_features[2775]  & (\all_features[2774]  | (new_n16243_ & (\all_features[2770]  | \all_features[2771]  | \all_features[2769] )));
  assign new_n16243_ = \all_features[2772]  & \all_features[2773] ;
  assign new_n16244_ = new_n16240_ & ~\all_features[2773]  & ~new_n16245_ & ~\all_features[2772] ;
  assign new_n16245_ = \all_features[2768]  & \all_features[2769] ;
  assign new_n16246_ = ~\all_features[2771]  & ~\all_features[2772]  & (~\all_features[2770]  | new_n16239_);
  assign new_n16247_ = ~new_n16248_ & ~new_n16250_;
  assign new_n16248_ = ~\all_features[2775]  & (~\all_features[2774]  | (~\all_features[2772]  & ~\all_features[2773]  & ~new_n16249_));
  assign new_n16249_ = \all_features[2770]  & \all_features[2771] ;
  assign new_n16250_ = ~\all_features[2775]  & (~\all_features[2774]  | (~\all_features[2773]  & (new_n16239_ | ~\all_features[2772]  | ~new_n16249_)));
  assign new_n16251_ = ~new_n16252_ & ~new_n16254_;
  assign new_n16252_ = new_n16253_ & (~\all_features[2771]  | ~new_n16243_ | (~\all_features[2770]  & ~new_n16245_));
  assign new_n16253_ = ~\all_features[2774]  & ~\all_features[2775] ;
  assign new_n16254_ = new_n16253_ & (~\all_features[2773]  | (~\all_features[2772]  & (~\all_features[2771]  | (~\all_features[2770]  & ~\all_features[2769] ))));
  assign new_n16255_ = ~new_n16256_ & ~new_n16257_;
  assign new_n16256_ = ~\all_features[2773]  & new_n16253_ & ((~\all_features[2770]  & new_n16239_) | ~\all_features[2772]  | ~\all_features[2771] );
  assign new_n16257_ = ~\all_features[2775]  & ~\all_features[2774]  & ~\all_features[2773]  & ~\all_features[2771]  & ~\all_features[2772] ;
  assign new_n16258_ = ~new_n16259_ & ~\all_features[2775] ;
  assign new_n16259_ = \all_features[2773]  & \all_features[2774]  & (\all_features[2772]  | (\all_features[2770]  & \all_features[2771]  & \all_features[2769] ));
  assign new_n16260_ = ~\all_features[2775]  & (~\all_features[2774]  | ~new_n16249_ | ~new_n16245_ | ~new_n16243_);
  assign new_n16261_ = new_n16255_ & ~new_n16262_ & new_n16251_;
  assign new_n16262_ = ~new_n16248_ & ~new_n16250_ & ~new_n16258_ & ~new_n16260_ & (~new_n16241_ | ~new_n16237_);
  assign new_n16263_ = new_n16251_ & new_n16247_ & new_n16255_ & ~new_n16258_ & ~new_n16260_;
  assign new_n16264_ = ~new_n15953_ & (~new_n15951_ | ~new_n15942_);
  assign new_n16265_ = ~new_n16227_ & new_n16154_;
  assign new_n16266_ = new_n16155_ & new_n16267_;
  assign new_n16267_ = new_n14626_ & new_n16268_;
  assign new_n16268_ = ~new_n16269_ & (new_n14650_ | (~new_n16272_ & ~new_n14648_));
  assign new_n16269_ = ~new_n14648_ & ~new_n14650_ & (~new_n14653_ | (~new_n16270_ & new_n14632_));
  assign new_n16270_ = new_n14636_ & ((~new_n16271_ & new_n14643_ & new_n14642_) | ~new_n14645_ | ~new_n14629_);
  assign new_n16271_ = new_n14644_ & \all_features[4845]  & ((~new_n14631_ & \all_features[4842] ) | \all_features[4844]  | \all_features[4843] );
  assign new_n16272_ = ~new_n14646_ & (new_n14649_ | (~new_n14633_ & (new_n14635_ | (~new_n14640_ & ~new_n16273_))));
  assign new_n16273_ = ~new_n14637_ & (~new_n14645_ | (new_n14629_ & (~new_n14642_ | (~new_n16274_ & new_n14643_))));
  assign new_n16274_ = new_n14644_ & (\all_features[4845]  | (\all_features[4844]  & (\all_features[4843]  | \all_features[4842] )));
  assign new_n16275_ = new_n16276_ & new_n16277_;
  assign new_n16276_ = new_n9653_ & new_n9686_;
  assign new_n16277_ = ~new_n9241_ & new_n9210_;
  assign new_n16278_ = new_n10644_ & new_n16279_;
  assign new_n16279_ = new_n6385_ & new_n6388_;
  assign new_n16280_ = new_n16316_ & new_n16304_ & ~new_n16281_ & new_n16283_;
  assign new_n16281_ = ~new_n12454_ & new_n16282_;
  assign new_n16282_ = ~new_n12487_ & ~new_n12490_;
  assign new_n16283_ = ~new_n16284_ & (\all_features[5275]  | \all_features[5276]  | \all_features[5277]  | \all_features[5278]  | \all_features[5279] );
  assign new_n16284_ = ~new_n16298_ & (new_n16300_ | (~new_n16301_ & (new_n16302_ | (~new_n16285_ & ~new_n16303_))));
  assign new_n16285_ = ~new_n16293_ & (new_n16295_ | (~new_n16286_ & new_n16297_));
  assign new_n16286_ = \all_features[5279]  & ((~new_n16291_ & ~\all_features[5277]  & \all_features[5278] ) | (~new_n16289_ & (\all_features[5278]  | (~new_n16287_ & \all_features[5277] ))));
  assign new_n16287_ = new_n16288_ & ~\all_features[5276]  & ~\all_features[5274]  & ~\all_features[5275] ;
  assign new_n16288_ = ~\all_features[5272]  & ~\all_features[5273] ;
  assign new_n16289_ = \all_features[5279]  & (\all_features[5278]  | (new_n16290_ & (\all_features[5274]  | \all_features[5275]  | \all_features[5273] )));
  assign new_n16290_ = \all_features[5276]  & \all_features[5277] ;
  assign new_n16291_ = (\all_features[5276]  & (\all_features[5274]  | \all_features[5275] )) | (~new_n16292_ & ~\all_features[5274]  & ~\all_features[5275]  & ~\all_features[5276] );
  assign new_n16292_ = \all_features[5272]  & \all_features[5273] ;
  assign new_n16293_ = ~new_n16294_ & ~\all_features[5279] ;
  assign new_n16294_ = \all_features[5277]  & \all_features[5278]  & (\all_features[5276]  | (\all_features[5274]  & \all_features[5275]  & \all_features[5273] ));
  assign new_n16295_ = ~\all_features[5279]  & (~\all_features[5278]  | ~new_n16292_ | ~new_n16290_ | ~new_n16296_);
  assign new_n16296_ = \all_features[5274]  & \all_features[5275] ;
  assign new_n16297_ = \all_features[5279]  & (\all_features[5277]  | \all_features[5278]  | \all_features[5276] );
  assign new_n16298_ = ~\all_features[5277]  & new_n16299_ & ((~\all_features[5274]  & new_n16288_) | ~\all_features[5276]  | ~\all_features[5275] );
  assign new_n16299_ = ~\all_features[5278]  & ~\all_features[5279] ;
  assign new_n16300_ = new_n16299_ & (~\all_features[5277]  | (~\all_features[5276]  & (~\all_features[5275]  | (~\all_features[5274]  & ~\all_features[5273] ))));
  assign new_n16301_ = new_n16299_ & (~\all_features[5275]  | ~new_n16290_ | (~\all_features[5274]  & ~new_n16292_));
  assign new_n16302_ = ~\all_features[5279]  & (~\all_features[5278]  | (~\all_features[5276]  & ~\all_features[5277]  & ~new_n16296_));
  assign new_n16303_ = ~\all_features[5279]  & (~\all_features[5278]  | (~\all_features[5277]  & (new_n16288_ | ~new_n16296_ | ~\all_features[5276] )));
  assign new_n16304_ = new_n16305_ & new_n16313_;
  assign new_n16305_ = new_n16306_ & (new_n16303_ | new_n16293_ | ~new_n16312_ | (new_n16310_ & new_n16309_));
  assign new_n16306_ = new_n16307_ & new_n16308_;
  assign new_n16307_ = ~new_n16298_ & (\all_features[5275]  | \all_features[5276]  | \all_features[5277]  | \all_features[5278]  | \all_features[5279] );
  assign new_n16308_ = ~new_n16300_ & ~new_n16301_;
  assign new_n16309_ = \all_features[5279]  & (\all_features[5278]  | (~new_n16287_ & \all_features[5277] ));
  assign new_n16310_ = \all_features[5279]  & \all_features[5278]  & ~new_n16311_ & new_n16289_;
  assign new_n16311_ = ~\all_features[5277]  & ~\all_features[5276]  & ~\all_features[5275]  & ~new_n16292_ & ~\all_features[5274] ;
  assign new_n16312_ = ~new_n16302_ & ~new_n16295_;
  assign new_n16313_ = new_n16315_ & new_n16306_ & new_n16314_;
  assign new_n16314_ = ~new_n16302_ & ~new_n16303_;
  assign new_n16315_ = ~new_n16293_ & ~new_n16295_;
  assign new_n16316_ = new_n16307_ & (~new_n16308_ | (new_n16314_ & (~new_n16315_ | new_n16317_)));
  assign new_n16317_ = new_n16309_ & (~new_n16310_ | (~new_n16318_ & \all_features[5277]  & \all_features[5278]  & \all_features[5279] ));
  assign new_n16318_ = ~\all_features[5275]  & ~\all_features[5276]  & (~\all_features[5274]  | new_n16288_);
  assign new_n16319_ = ~new_n16267_ & new_n16155_;
  assign new_n16320_ = new_n16321_ & (new_n16322_ | new_n16275_ | ~new_n16266_);
  assign new_n16321_ = (~new_n16229_ | (new_n16232_ ? new_n16233_ : new_n16230_)) & (~new_n16265_ | new_n16278_);
  assign new_n16322_ = ~new_n16276_ & ~new_n15598_;
  assign new_n16323_ = (~new_n16266_ | ~new_n16322_) & (~new_n16319_ | ~new_n16280_) & (~new_n16153_ | ~new_n16264_);
  assign new_n16324_ = new_n16325_ ? (~new_n16654_ ^ new_n16751_) : (new_n16654_ ^ new_n16751_);
  assign new_n16325_ = new_n16326_ ? (~new_n16520_ ^ new_n16644_) : (new_n16520_ ^ new_n16644_);
  assign new_n16326_ = new_n16327_ ? (new_n15907_ ^ new_n16451_) : (~new_n15907_ ^ new_n16451_);
  assign new_n16327_ = new_n16328_ ? (new_n16372_ ^ new_n16373_) : (~new_n16372_ ^ new_n16373_);
  assign new_n16328_ = ~new_n16329_ & new_n16368_;
  assign new_n16329_ = new_n16330_ & (~new_n16362_ | ~new_n16352_);
  assign new_n16330_ = ~new_n16346_ & ~new_n16331_ & (~new_n16342_ | (new_n16351_ & new_n13922_) | (new_n16349_ & ~new_n13922_));
  assign new_n16331_ = new_n16332_ & (new_n15671_ ? ~new_n7991_ : ~new_n16336_);
  assign new_n16332_ = ~new_n16335_ & new_n16333_;
  assign new_n16333_ = new_n9867_ & (new_n9864_ | ~new_n16334_);
  assign new_n16334_ = ~new_n9836_ & ~new_n9860_;
  assign new_n16335_ = ~new_n10596_ & new_n12152_;
  assign new_n16336_ = ~new_n16338_ & new_n16337_;
  assign new_n16337_ = ~new_n15797_ & ~new_n15819_;
  assign new_n16338_ = new_n15814_ & (new_n15818_ | new_n15817_ | (~new_n15800_ & ~new_n15805_ & ~new_n16339_));
  assign new_n16339_ = ~new_n15806_ & ~new_n15803_ & (~new_n15813_ | ~new_n15809_ | new_n16340_);
  assign new_n16340_ = new_n15811_ & new_n15812_ & (new_n16341_ | ~\all_features[989]  | ~\all_features[990]  | ~\all_features[991] );
  assign new_n16341_ = ~\all_features[987]  & ~\all_features[988]  & (~\all_features[986]  | new_n15801_);
  assign new_n16342_ = ~new_n16333_ & ~new_n16343_;
  assign new_n16343_ = new_n16344_ & new_n16345_;
  assign new_n16344_ = new_n10002_ & new_n10024_;
  assign new_n16345_ = new_n10028_ & new_n10032_;
  assign new_n16346_ = new_n16335_ & new_n16333_ & new_n16347_;
  assign new_n16347_ = new_n16348_ & new_n9640_;
  assign new_n16348_ = new_n9612_ & new_n9634_;
  assign new_n16349_ = new_n14235_ & (new_n14212_ | ~new_n16350_);
  assign new_n16350_ = ~new_n14620_ & ~new_n14237_;
  assign new_n16351_ = new_n9129_ & (new_n9131_ | ~new_n12448_);
  assign new_n16352_ = ~new_n16353_ & new_n16361_;
  assign new_n16353_ = new_n16354_ & new_n9995_;
  assign new_n16354_ = ~new_n16355_ & new_n9993_;
  assign new_n16355_ = ~new_n9968_ & ~new_n16356_;
  assign new_n16356_ = ~new_n9974_ & (new_n9970_ | (~new_n9989_ & (new_n9988_ | (~new_n9984_ & ~new_n16357_))));
  assign new_n16357_ = ~new_n9986_ & (new_n9990_ | (~new_n9992_ & (~new_n16360_ | new_n16358_)));
  assign new_n16358_ = \all_features[2991]  & ((~new_n16359_ & ~\all_features[2989]  & \all_features[2990] ) | (~new_n9979_ & (\all_features[2990]  | (~new_n9977_ & \all_features[2989] ))));
  assign new_n16359_ = (~\all_features[2986]  & ~\all_features[2987]  & ~\all_features[2988]  & (~\all_features[2985]  | ~\all_features[2984] )) | (\all_features[2988]  & (\all_features[2986]  | \all_features[2987] ));
  assign new_n16360_ = \all_features[2991]  & (\all_features[2989]  | \all_features[2990]  | \all_features[2988] );
  assign new_n16361_ = ~new_n16333_ & new_n16343_;
  assign new_n16362_ = ~new_n16363_ & new_n14038_;
  assign new_n16363_ = new_n14014_ & new_n16364_;
  assign new_n16364_ = ~new_n16365_ & (\all_features[2555]  | \all_features[2556]  | \all_features[2557]  | \all_features[2558]  | \all_features[2559] );
  assign new_n16365_ = ~new_n14036_ & (new_n14032_ | (~new_n14030_ & (new_n14037_ | (~new_n14033_ & ~new_n16366_))));
  assign new_n16366_ = ~new_n14026_ & (new_n14025_ | (new_n14028_ & (~new_n14024_ | (~new_n16367_ & new_n14017_))));
  assign new_n16367_ = ~\all_features[2557]  & \all_features[2558]  & \all_features[2559]  & (\all_features[2556]  ? new_n14021_ : (new_n14020_ | ~new_n14021_));
  assign new_n16368_ = new_n16371_ & new_n16369_ & new_n16370_;
  assign new_n16369_ = (~new_n16352_ | new_n16362_) & (~new_n16342_ | (new_n13922_ ? ~new_n16351_ : ~new_n16349_));
  assign new_n16370_ = (~new_n16332_ | ~new_n15671_ | ~new_n7991_) & (new_n12758_ | ~new_n16361_ | ~new_n16353_);
  assign new_n16371_ = ~new_n16333_ | ((new_n16347_ | ~new_n16335_) & (new_n15671_ | ~new_n16336_ | new_n16335_));
  assign new_n16372_ = ~new_n14614_ & new_n14865_;
  assign new_n16373_ = new_n16417_ & (new_n16374_ | new_n16446_ | ~new_n16450_);
  assign new_n16374_ = new_n16410_ ? new_n16375_ : (new_n15082_ | (new_n15049_ & new_n15079_));
  assign new_n16375_ = ~new_n16406_ & new_n16376_;
  assign new_n16376_ = ~new_n16402_ & new_n16377_;
  assign new_n16377_ = ~new_n16378_ & ~new_n16400_;
  assign new_n16378_ = new_n16395_ & ~new_n16399_ & ~new_n16379_ & ~new_n16398_;
  assign new_n16379_ = new_n16380_ & (~new_n16393_ | ~new_n16394_ | ~new_n16390_ | ~new_n16392_);
  assign new_n16380_ = ~new_n16387_ & ~new_n16385_ & ~new_n16381_ & ~new_n16383_;
  assign new_n16381_ = ~\all_features[2863]  & (~\all_features[2862]  | (~\all_features[2860]  & ~\all_features[2861]  & ~new_n16382_));
  assign new_n16382_ = \all_features[2858]  & \all_features[2859] ;
  assign new_n16383_ = ~\all_features[2863]  & (~\all_features[2862]  | (~\all_features[2861]  & (new_n16384_ | ~new_n16382_ | ~\all_features[2860] )));
  assign new_n16384_ = ~\all_features[2856]  & ~\all_features[2857] ;
  assign new_n16385_ = ~new_n16386_ & ~\all_features[2863] ;
  assign new_n16386_ = \all_features[2861]  & \all_features[2862]  & (\all_features[2860]  | (\all_features[2858]  & \all_features[2859]  & \all_features[2857] ));
  assign new_n16387_ = ~\all_features[2863]  & (~\all_features[2862]  | ~new_n16388_ | ~new_n16389_ | ~new_n16382_);
  assign new_n16388_ = \all_features[2856]  & \all_features[2857] ;
  assign new_n16389_ = \all_features[2860]  & \all_features[2861] ;
  assign new_n16390_ = \all_features[2863]  & (\all_features[2862]  | (\all_features[2861]  & (\all_features[2860]  | ~new_n16391_ | ~new_n16384_)));
  assign new_n16391_ = ~\all_features[2858]  & ~\all_features[2859] ;
  assign new_n16392_ = \all_features[2863]  & (\all_features[2862]  | (new_n16389_ & (\all_features[2858]  | \all_features[2859]  | \all_features[2857] )));
  assign new_n16393_ = \all_features[2862]  & \all_features[2863]  & (\all_features[2860]  | \all_features[2861]  | new_n16388_ | ~new_n16391_);
  assign new_n16394_ = \all_features[2863]  & (\all_features[2861]  | \all_features[2862]  | \all_features[2860] );
  assign new_n16395_ = ~new_n16396_ & (\all_features[2859]  | \all_features[2860]  | \all_features[2861]  | \all_features[2862]  | \all_features[2863] );
  assign new_n16396_ = ~\all_features[2861]  & new_n16397_ & ((~\all_features[2858]  & new_n16384_) | ~\all_features[2860]  | ~\all_features[2859] );
  assign new_n16397_ = ~\all_features[2862]  & ~\all_features[2863] ;
  assign new_n16398_ = new_n16397_ & (~\all_features[2861]  | (~\all_features[2860]  & (~\all_features[2859]  | (~\all_features[2858]  & ~\all_features[2857] ))));
  assign new_n16399_ = new_n16397_ & (~\all_features[2859]  | ~new_n16389_ | (~\all_features[2858]  & ~new_n16388_));
  assign new_n16400_ = new_n16401_ & new_n16395_ & ~new_n16398_ & ~new_n16385_;
  assign new_n16401_ = ~new_n16387_ & ~new_n16383_ & ~new_n16399_ & ~new_n16381_;
  assign new_n16402_ = new_n16395_ & (new_n16399_ | new_n16398_ | (~new_n16403_ & ~new_n16381_ & ~new_n16383_));
  assign new_n16403_ = ~new_n16385_ & ~new_n16387_ & (~new_n16394_ | ~new_n16390_ | new_n16404_);
  assign new_n16404_ = new_n16392_ & new_n16393_ & (new_n16405_ | ~\all_features[2861]  | ~\all_features[2862]  | ~\all_features[2863] );
  assign new_n16405_ = ~\all_features[2859]  & ~\all_features[2860]  & (~\all_features[2858]  | new_n16384_);
  assign new_n16406_ = ~new_n16407_ & (\all_features[2859]  | \all_features[2860]  | \all_features[2861]  | \all_features[2862]  | \all_features[2863] );
  assign new_n16407_ = ~new_n16396_ & (new_n16398_ | (~new_n16399_ & (new_n16381_ | (~new_n16408_ & ~new_n16383_))));
  assign new_n16408_ = ~new_n16385_ & (new_n16387_ | (new_n16394_ & (~new_n16390_ | (~new_n16409_ & new_n16392_))));
  assign new_n16409_ = ~\all_features[2861]  & \all_features[2862]  & \all_features[2863]  & (\all_features[2860]  ? new_n16391_ : (new_n16388_ | ~new_n16391_));
  assign new_n16410_ = ~new_n16411_ & new_n8268_;
  assign new_n16411_ = new_n16412_ & new_n8295_;
  assign new_n16412_ = (new_n16413_ | (new_n8279_ & (~\all_features[3203]  | ~\all_features[3204]  | (~\all_features[3202]  & new_n8278_)))) & (~new_n8279_ | \all_features[3203]  | \all_features[3204] );
  assign new_n16413_ = ~new_n8275_ & (new_n8272_ | (~new_n8286_ & (new_n8289_ | (~new_n16414_ & ~new_n8290_))));
  assign new_n16414_ = ~new_n8288_ & (~\all_features[3207]  | new_n16415_ | (~\all_features[3204]  & ~\all_features[3205]  & ~\all_features[3206] ));
  assign new_n16415_ = \all_features[3207]  & ((~new_n16416_ & ~\all_features[3205]  & \all_features[3206] ) | (~new_n8283_ & (\all_features[3206]  | (~new_n8281_ & \all_features[3205] ))));
  assign new_n16416_ = (\all_features[3204]  & (\all_features[3202]  | \all_features[3203] )) | (~new_n8273_ & ~\all_features[3202]  & ~\all_features[3203]  & ~\all_features[3204] );
  assign new_n16417_ = ~new_n16446_ & (~new_n16448_ | (~new_n16442_ & ~new_n16418_));
  assign new_n16418_ = new_n16434_ & (~new_n16437_ | (~new_n16419_ & ~new_n16440_ & ~new_n16441_));
  assign new_n16419_ = ~new_n16428_ & ~new_n16430_ & (~new_n16433_ | ~new_n16432_ | new_n16420_);
  assign new_n16420_ = new_n16421_ & new_n16423_ & (new_n16426_ | ~\all_features[5733]  | ~\all_features[5734]  | ~\all_features[5735] );
  assign new_n16421_ = \all_features[5735]  & (\all_features[5734]  | (new_n16422_ & (\all_features[5730]  | \all_features[5731]  | \all_features[5729] )));
  assign new_n16422_ = \all_features[5732]  & \all_features[5733] ;
  assign new_n16423_ = \all_features[5734]  & \all_features[5735]  & (\all_features[5732]  | \all_features[5733]  | new_n16424_ | ~new_n16425_);
  assign new_n16424_ = \all_features[5728]  & \all_features[5729] ;
  assign new_n16425_ = ~\all_features[5730]  & ~\all_features[5731] ;
  assign new_n16426_ = ~\all_features[5731]  & ~\all_features[5732]  & (~\all_features[5730]  | new_n16427_);
  assign new_n16427_ = ~\all_features[5728]  & ~\all_features[5729] ;
  assign new_n16428_ = ~new_n16429_ & ~\all_features[5735] ;
  assign new_n16429_ = \all_features[5733]  & \all_features[5734]  & (\all_features[5732]  | (\all_features[5730]  & \all_features[5731]  & \all_features[5729] ));
  assign new_n16430_ = ~\all_features[5735]  & (~\all_features[5734]  | ~new_n16431_ | ~new_n16424_ | ~new_n16422_);
  assign new_n16431_ = \all_features[5730]  & \all_features[5731] ;
  assign new_n16432_ = \all_features[5735]  & (\all_features[5734]  | (\all_features[5733]  & (\all_features[5732]  | ~new_n16425_ | ~new_n16427_)));
  assign new_n16433_ = \all_features[5735]  & (\all_features[5733]  | \all_features[5734]  | \all_features[5732] );
  assign new_n16434_ = ~new_n16435_ & (\all_features[5731]  | \all_features[5732]  | \all_features[5733]  | \all_features[5734]  | \all_features[5735] );
  assign new_n16435_ = ~\all_features[5733]  & new_n16436_ & ((~\all_features[5730]  & new_n16427_) | ~\all_features[5732]  | ~\all_features[5731] );
  assign new_n16436_ = ~\all_features[5734]  & ~\all_features[5735] ;
  assign new_n16437_ = ~new_n16438_ & ~new_n16439_;
  assign new_n16438_ = new_n16436_ & (~\all_features[5733]  | (~\all_features[5732]  & (~\all_features[5731]  | (~\all_features[5730]  & ~\all_features[5729] ))));
  assign new_n16439_ = new_n16436_ & (~\all_features[5731]  | ~new_n16422_ | (~\all_features[5730]  & ~new_n16424_));
  assign new_n16440_ = ~\all_features[5735]  & (~\all_features[5734]  | (~\all_features[5733]  & (new_n16427_ | ~new_n16431_ | ~\all_features[5732] )));
  assign new_n16441_ = ~\all_features[5735]  & (~\all_features[5734]  | (~\all_features[5732]  & ~\all_features[5733]  & ~new_n16431_));
  assign new_n16442_ = ~new_n16443_ & (\all_features[5731]  | \all_features[5732]  | \all_features[5733]  | \all_features[5734]  | \all_features[5735] );
  assign new_n16443_ = ~new_n16435_ & (new_n16438_ | (~new_n16439_ & (new_n16441_ | (~new_n16440_ & ~new_n16444_))));
  assign new_n16444_ = ~new_n16428_ & (new_n16430_ | (new_n16433_ & (~new_n16432_ | (~new_n16445_ & new_n16421_))));
  assign new_n16445_ = ~\all_features[5733]  & \all_features[5734]  & \all_features[5735]  & (\all_features[5732]  ? new_n16425_ : (new_n16424_ | ~new_n16425_));
  assign new_n16446_ = new_n16447_ & new_n16434_ & ~new_n16439_ & ~new_n16440_ & ~new_n16428_ & ~new_n16438_;
  assign new_n16447_ = ~new_n16430_ & ~new_n16441_;
  assign new_n16448_ = new_n16434_ & new_n16437_ & (new_n16449_ | new_n16428_ | new_n16440_ | ~new_n16447_);
  assign new_n16449_ = new_n16433_ & new_n16423_ & new_n16432_ & new_n16421_;
  assign new_n16450_ = ~new_n16418_ & ~new_n16448_;
  assign new_n16451_ = (~new_n12825_ | ~new_n12834_) & ((~new_n16519_ & ~new_n8164_ & new_n16485_) | (~new_n16452_ & ~new_n16485_));
  assign new_n16452_ = (new_n16453_ & new_n13328_) | (new_n16455_ & new_n16482_ & ~new_n13328_);
  assign new_n16453_ = ~new_n6461_ & new_n16454_;
  assign new_n16454_ = ~new_n6491_ & ~new_n6495_;
  assign new_n16455_ = new_n16456_ & new_n16479_;
  assign new_n16456_ = new_n16457_ & (new_n16476_ | new_n16477_ | ~new_n16472_ | (new_n16469_ & new_n16467_));
  assign new_n16457_ = new_n16458_ & new_n16464_;
  assign new_n16458_ = ~new_n16459_ & ~new_n16462_;
  assign new_n16459_ = ~\all_features[1462]  & ~\all_features[1463]  & (~\all_features[1459]  | ~new_n16461_ | (~\all_features[1458]  & ~new_n16460_));
  assign new_n16460_ = \all_features[1456]  & \all_features[1457] ;
  assign new_n16461_ = \all_features[1460]  & \all_features[1461] ;
  assign new_n16462_ = ~\all_features[1463]  & ~new_n16463_ & ~\all_features[1462] ;
  assign new_n16463_ = \all_features[1461]  & (\all_features[1460]  | (\all_features[1459]  & (\all_features[1458]  | \all_features[1457] )));
  assign new_n16464_ = ~new_n16466_ | (\all_features[1459]  & \all_features[1460]  & (\all_features[1458]  | ~new_n16465_));
  assign new_n16465_ = ~\all_features[1456]  & ~\all_features[1457] ;
  assign new_n16466_ = ~\all_features[1463]  & ~\all_features[1461]  & ~\all_features[1462] ;
  assign new_n16467_ = \all_features[1463]  & (\all_features[1462]  | (~new_n16468_ & \all_features[1461] ));
  assign new_n16468_ = new_n16465_ & ~\all_features[1460]  & ~\all_features[1458]  & ~\all_features[1459] ;
  assign new_n16469_ = \all_features[1463]  & \all_features[1462]  & ~new_n16471_ & new_n16470_;
  assign new_n16470_ = \all_features[1463]  & (\all_features[1462]  | (new_n16461_ & (\all_features[1458]  | \all_features[1459]  | \all_features[1457] )));
  assign new_n16471_ = ~\all_features[1461]  & ~\all_features[1460]  & ~\all_features[1459]  & ~new_n16460_ & ~\all_features[1458] ;
  assign new_n16472_ = ~new_n16473_ & ~new_n16475_;
  assign new_n16473_ = ~\all_features[1463]  & (~\all_features[1462]  | (~\all_features[1460]  & ~\all_features[1461]  & ~new_n16474_));
  assign new_n16474_ = \all_features[1458]  & \all_features[1459] ;
  assign new_n16475_ = ~\all_features[1463]  & (~\all_features[1462]  | ~new_n16460_ | ~new_n16461_ | ~new_n16474_);
  assign new_n16476_ = ~\all_features[1463]  & (~\all_features[1462]  | (~\all_features[1461]  & (new_n16465_ | ~new_n16474_ | ~\all_features[1460] )));
  assign new_n16477_ = ~new_n16478_ & ~\all_features[1463] ;
  assign new_n16478_ = \all_features[1461]  & \all_features[1462]  & (\all_features[1460]  | (\all_features[1458]  & \all_features[1459]  & \all_features[1457] ));
  assign new_n16479_ = new_n16481_ & new_n16457_ & new_n16480_;
  assign new_n16480_ = ~new_n16473_ & ~new_n16476_;
  assign new_n16481_ = ~new_n16475_ & ~new_n16477_;
  assign new_n16482_ = new_n16464_ & (~new_n16458_ | (new_n16480_ & (~new_n16481_ | new_n16483_)));
  assign new_n16483_ = new_n16467_ & (~new_n16469_ | (~new_n16484_ & \all_features[1461]  & \all_features[1462]  & \all_features[1463] ));
  assign new_n16484_ = ~\all_features[1459]  & ~\all_features[1460]  & (~\all_features[1458]  | new_n16465_);
  assign new_n16485_ = new_n16486_ & ~new_n16515_ & ~new_n16518_;
  assign new_n16486_ = ~new_n16487_ & ~new_n16508_;
  assign new_n16487_ = ~new_n16488_ & (\all_features[4083]  | \all_features[4084]  | \all_features[4085]  | \all_features[4086]  | \all_features[4087] );
  assign new_n16488_ = ~new_n16502_ & (new_n16504_ | (~new_n16505_ & (new_n16506_ | (~new_n16489_ & ~new_n16507_))));
  assign new_n16489_ = ~new_n16490_ & (new_n16492_ | (new_n16501_ & (~new_n16496_ | (~new_n16500_ & new_n16499_))));
  assign new_n16490_ = ~new_n16491_ & ~\all_features[4087] ;
  assign new_n16491_ = \all_features[4085]  & \all_features[4086]  & (\all_features[4084]  | (\all_features[4082]  & \all_features[4083]  & \all_features[4081] ));
  assign new_n16492_ = ~\all_features[4087]  & (~\all_features[4086]  | ~new_n16493_ | ~new_n16494_ | ~new_n16495_);
  assign new_n16493_ = \all_features[4080]  & \all_features[4081] ;
  assign new_n16494_ = \all_features[4084]  & \all_features[4085] ;
  assign new_n16495_ = \all_features[4082]  & \all_features[4083] ;
  assign new_n16496_ = \all_features[4087]  & (\all_features[4086]  | (\all_features[4085]  & (\all_features[4084]  | ~new_n16498_ | ~new_n16497_)));
  assign new_n16497_ = ~\all_features[4080]  & ~\all_features[4081] ;
  assign new_n16498_ = ~\all_features[4082]  & ~\all_features[4083] ;
  assign new_n16499_ = \all_features[4087]  & (\all_features[4086]  | (new_n16494_ & (\all_features[4082]  | \all_features[4083]  | \all_features[4081] )));
  assign new_n16500_ = ~\all_features[4085]  & \all_features[4086]  & \all_features[4087]  & (\all_features[4084]  ? new_n16498_ : (new_n16493_ | ~new_n16498_));
  assign new_n16501_ = \all_features[4087]  & (\all_features[4085]  | \all_features[4086]  | \all_features[4084] );
  assign new_n16502_ = ~\all_features[4085]  & new_n16503_ & ((~\all_features[4082]  & new_n16497_) | ~\all_features[4084]  | ~\all_features[4083] );
  assign new_n16503_ = ~\all_features[4086]  & ~\all_features[4087] ;
  assign new_n16504_ = new_n16503_ & (~\all_features[4085]  | (~\all_features[4084]  & (~\all_features[4083]  | (~\all_features[4082]  & ~\all_features[4081] ))));
  assign new_n16505_ = new_n16503_ & (~\all_features[4083]  | ~new_n16494_ | (~\all_features[4082]  & ~new_n16493_));
  assign new_n16506_ = ~\all_features[4087]  & (~\all_features[4086]  | (~\all_features[4084]  & ~\all_features[4085]  & ~new_n16495_));
  assign new_n16507_ = ~\all_features[4087]  & (~\all_features[4086]  | (~\all_features[4085]  & (new_n16497_ | ~new_n16495_ | ~\all_features[4084] )));
  assign new_n16508_ = new_n16514_ & (~new_n16513_ | (~new_n16509_ & ~new_n16506_ & ~new_n16507_));
  assign new_n16509_ = ~new_n16490_ & ~new_n16492_ & (~new_n16501_ | ~new_n16496_ | new_n16510_);
  assign new_n16510_ = new_n16499_ & new_n16511_ & (new_n16512_ | ~\all_features[4085]  | ~\all_features[4086]  | ~\all_features[4087] );
  assign new_n16511_ = \all_features[4086]  & \all_features[4087]  & (\all_features[4084]  | \all_features[4085]  | new_n16493_ | ~new_n16498_);
  assign new_n16512_ = ~\all_features[4083]  & ~\all_features[4084]  & (~\all_features[4082]  | new_n16497_);
  assign new_n16513_ = ~new_n16504_ & ~new_n16505_;
  assign new_n16514_ = ~new_n16502_ & (\all_features[4083]  | \all_features[4084]  | \all_features[4085]  | \all_features[4086]  | \all_features[4087] );
  assign new_n16515_ = new_n16513_ & new_n16514_ & (new_n16516_ | new_n16507_ | new_n16492_ | ~new_n16517_);
  assign new_n16516_ = new_n16501_ & new_n16511_ & new_n16496_ & new_n16499_;
  assign new_n16517_ = ~new_n16506_ & ~new_n16490_;
  assign new_n16518_ = new_n16514_ & new_n16513_ & new_n16517_ & ~new_n16507_ & ~new_n16492_;
  assign new_n16519_ = ~new_n11823_ & new_n11793_;
  assign new_n16520_ = new_n16572_ & (~new_n16521_ | ((~new_n16609_ | ~new_n16574_) & (~new_n16568_ | ~new_n16610_)));
  assign new_n16521_ = ~new_n16563_ & new_n16522_ & (~new_n16569_ | ~new_n16568_);
  assign new_n16522_ = (~new_n16523_ | new_n13349_ | ~new_n16524_) & (new_n16527_ | ~new_n16525_ | ~new_n13405_ | new_n16524_);
  assign new_n16523_ = ~new_n15713_ & new_n9058_;
  assign new_n16524_ = new_n9690_ & new_n12906_;
  assign new_n16525_ = new_n16526_ & new_n10729_;
  assign new_n16526_ = new_n10703_ & new_n10726_;
  assign new_n16527_ = ~new_n16528_ & new_n16558_;
  assign new_n16528_ = new_n16529_ & new_n16550_;
  assign new_n16529_ = ~new_n16530_ & (\all_features[3235]  | \all_features[3236]  | \all_features[3237]  | \all_features[3238]  | \all_features[3239] );
  assign new_n16530_ = ~new_n16544_ & (new_n16549_ | (~new_n16546_ & (new_n16547_ | (~new_n16548_ & ~new_n16531_))));
  assign new_n16531_ = ~new_n16532_ & (new_n16541_ | (new_n16543_ & (~new_n16534_ | (~new_n16539_ & new_n16537_))));
  assign new_n16532_ = ~new_n16533_ & ~\all_features[3239] ;
  assign new_n16533_ = \all_features[3237]  & \all_features[3238]  & (\all_features[3236]  | (\all_features[3234]  & \all_features[3235]  & \all_features[3233] ));
  assign new_n16534_ = \all_features[3239]  & (\all_features[3238]  | (\all_features[3237]  & (\all_features[3236]  | ~new_n16536_ | ~new_n16535_)));
  assign new_n16535_ = ~\all_features[3232]  & ~\all_features[3233] ;
  assign new_n16536_ = ~\all_features[3234]  & ~\all_features[3235] ;
  assign new_n16537_ = \all_features[3239]  & (\all_features[3238]  | (new_n16538_ & (\all_features[3234]  | \all_features[3235]  | \all_features[3233] )));
  assign new_n16538_ = \all_features[3236]  & \all_features[3237] ;
  assign new_n16539_ = ~\all_features[3237]  & \all_features[3238]  & \all_features[3239]  & (\all_features[3236]  ? new_n16536_ : (new_n16540_ | ~new_n16536_));
  assign new_n16540_ = \all_features[3232]  & \all_features[3233] ;
  assign new_n16541_ = ~\all_features[3239]  & (~\all_features[3238]  | ~new_n16540_ | ~new_n16538_ | ~new_n16542_);
  assign new_n16542_ = \all_features[3234]  & \all_features[3235] ;
  assign new_n16543_ = \all_features[3239]  & (\all_features[3237]  | \all_features[3238]  | \all_features[3236] );
  assign new_n16544_ = ~\all_features[3237]  & new_n16545_ & ((~\all_features[3234]  & new_n16535_) | ~\all_features[3236]  | ~\all_features[3235] );
  assign new_n16545_ = ~\all_features[3238]  & ~\all_features[3239] ;
  assign new_n16546_ = new_n16545_ & (~\all_features[3235]  | ~new_n16538_ | (~\all_features[3234]  & ~new_n16540_));
  assign new_n16547_ = ~\all_features[3239]  & (~\all_features[3238]  | (~\all_features[3236]  & ~\all_features[3237]  & ~new_n16542_));
  assign new_n16548_ = ~\all_features[3239]  & (~\all_features[3238]  | (~\all_features[3237]  & (new_n16535_ | ~new_n16542_ | ~\all_features[3236] )));
  assign new_n16549_ = new_n16545_ & (~\all_features[3237]  | (~\all_features[3236]  & (~\all_features[3235]  | (~\all_features[3234]  & ~\all_features[3233] ))));
  assign new_n16550_ = new_n16556_ & (~new_n16557_ | (~new_n16551_ & ~new_n16547_ & ~new_n16548_));
  assign new_n16551_ = new_n16554_ & ((~new_n16552_ & new_n16537_ & new_n16555_) | ~new_n16543_ | ~new_n16534_);
  assign new_n16552_ = \all_features[3239]  & \all_features[3238]  & ~new_n16553_ & \all_features[3237] ;
  assign new_n16553_ = ~\all_features[3235]  & ~\all_features[3236]  & (~\all_features[3234]  | new_n16535_);
  assign new_n16554_ = ~new_n16532_ & ~new_n16541_;
  assign new_n16555_ = \all_features[3238]  & \all_features[3239]  & (\all_features[3236]  | \all_features[3237]  | new_n16540_ | ~new_n16536_);
  assign new_n16556_ = ~new_n16544_ & (\all_features[3235]  | \all_features[3236]  | \all_features[3237]  | \all_features[3238]  | \all_features[3239] );
  assign new_n16557_ = ~new_n16546_ & ~new_n16549_;
  assign new_n16558_ = ~new_n16559_ & ~new_n16562_;
  assign new_n16559_ = new_n16557_ & ~new_n16560_ & new_n16556_;
  assign new_n16560_ = new_n16561_ & (~new_n16555_ | ~new_n16543_ | ~new_n16534_ | ~new_n16537_);
  assign new_n16561_ = ~new_n16541_ & ~new_n16532_ & ~new_n16547_ & ~new_n16548_;
  assign new_n16562_ = new_n16554_ & new_n16556_ & ~new_n16549_ & ~new_n16548_ & ~new_n16546_ & ~new_n16547_;
  assign new_n16563_ = ~new_n16524_ & (new_n16527_ ? ~new_n16564_ : ~new_n16525_);
  assign new_n16564_ = (new_n16565_ & new_n16567_) | (~new_n16268_ & new_n14627_ & new_n14651_ & ~new_n16567_);
  assign new_n16565_ = new_n12187_ & (new_n12185_ | ~new_n16566_);
  assign new_n16566_ = ~new_n12155_ & ~new_n12175_;
  assign new_n16567_ = ~new_n13971_ & ~new_n13975_;
  assign new_n16568_ = new_n16524_ & new_n13349_;
  assign new_n16569_ = ~new_n7445_ & new_n16570_;
  assign new_n16570_ = ~new_n13921_ & new_n16571_;
  assign new_n16571_ = ~new_n13909_ & ~new_n13918_;
  assign new_n16572_ = new_n16573_ & (new_n16569_ | new_n16610_ | ~new_n16568_);
  assign new_n16573_ = new_n16608_ & (new_n16574_ | new_n16523_ | ~new_n16609_);
  assign new_n16574_ = new_n15713_ & (~new_n16607_ | ~new_n16603_ | (~new_n16596_ & ~new_n16575_));
  assign new_n16575_ = ~new_n16576_ & (\all_features[4611]  | \all_features[4612]  | \all_features[4613]  | \all_features[4614]  | \all_features[4615] );
  assign new_n16576_ = ~new_n16590_ & (new_n16592_ | (~new_n16593_ & (new_n16594_ | (~new_n16577_ & ~new_n16595_))));
  assign new_n16577_ = ~new_n16578_ & (new_n16580_ | (new_n16589_ & (~new_n16584_ | (~new_n16588_ & new_n16587_))));
  assign new_n16578_ = ~new_n16579_ & ~\all_features[4615] ;
  assign new_n16579_ = \all_features[4613]  & \all_features[4614]  & (\all_features[4612]  | (\all_features[4610]  & \all_features[4611]  & \all_features[4609] ));
  assign new_n16580_ = ~\all_features[4615]  & (~\all_features[4614]  | ~new_n16581_ | ~new_n16582_ | ~new_n16583_);
  assign new_n16581_ = \all_features[4608]  & \all_features[4609] ;
  assign new_n16582_ = \all_features[4612]  & \all_features[4613] ;
  assign new_n16583_ = \all_features[4610]  & \all_features[4611] ;
  assign new_n16584_ = \all_features[4615]  & (\all_features[4614]  | (\all_features[4613]  & (\all_features[4612]  | ~new_n16586_ | ~new_n16585_)));
  assign new_n16585_ = ~\all_features[4608]  & ~\all_features[4609] ;
  assign new_n16586_ = ~\all_features[4610]  & ~\all_features[4611] ;
  assign new_n16587_ = \all_features[4615]  & (\all_features[4614]  | (new_n16582_ & (\all_features[4610]  | \all_features[4611]  | \all_features[4609] )));
  assign new_n16588_ = ~\all_features[4613]  & \all_features[4614]  & \all_features[4615]  & (\all_features[4612]  ? new_n16586_ : (new_n16581_ | ~new_n16586_));
  assign new_n16589_ = \all_features[4615]  & (\all_features[4613]  | \all_features[4614]  | \all_features[4612] );
  assign new_n16590_ = ~\all_features[4613]  & new_n16591_ & ((~\all_features[4610]  & new_n16585_) | ~\all_features[4612]  | ~\all_features[4611] );
  assign new_n16591_ = ~\all_features[4614]  & ~\all_features[4615] ;
  assign new_n16592_ = new_n16591_ & (~\all_features[4613]  | (~\all_features[4612]  & (~\all_features[4611]  | (~\all_features[4610]  & ~\all_features[4609] ))));
  assign new_n16593_ = new_n16591_ & (~\all_features[4611]  | ~new_n16582_ | (~\all_features[4610]  & ~new_n16581_));
  assign new_n16594_ = ~\all_features[4615]  & (~\all_features[4614]  | (~\all_features[4612]  & ~\all_features[4613]  & ~new_n16583_));
  assign new_n16595_ = ~\all_features[4615]  & (~\all_features[4614]  | (~\all_features[4613]  & (new_n16585_ | ~new_n16583_ | ~\all_features[4612] )));
  assign new_n16596_ = new_n16601_ & (~new_n16602_ | (~new_n16597_ & ~new_n16594_ & ~new_n16595_));
  assign new_n16597_ = ~new_n16578_ & ~new_n16580_ & (~new_n16589_ | ~new_n16584_ | new_n16598_);
  assign new_n16598_ = new_n16587_ & new_n16599_ & (new_n16600_ | ~\all_features[4613]  | ~\all_features[4614]  | ~\all_features[4615] );
  assign new_n16599_ = \all_features[4614]  & \all_features[4615]  & (\all_features[4612]  | \all_features[4613]  | new_n16581_ | ~new_n16586_);
  assign new_n16600_ = ~\all_features[4611]  & ~\all_features[4612]  & (~\all_features[4610]  | new_n16585_);
  assign new_n16601_ = ~new_n16590_ & (\all_features[4611]  | \all_features[4612]  | \all_features[4613]  | \all_features[4614]  | \all_features[4615] );
  assign new_n16602_ = ~new_n16592_ & ~new_n16593_;
  assign new_n16603_ = new_n16606_ & ~new_n16592_ & ~new_n16604_ & ~new_n16590_;
  assign new_n16604_ = new_n16605_ & ~new_n16595_ & (~new_n16599_ | ~new_n16589_ | ~new_n16584_ | ~new_n16587_);
  assign new_n16605_ = ~new_n16580_ & ~new_n16594_ & ~new_n16578_;
  assign new_n16606_ = ~new_n16593_ & (\all_features[4611]  | \all_features[4612]  | \all_features[4613]  | \all_features[4614]  | \all_features[4615] );
  assign new_n16607_ = new_n16601_ & new_n16605_ & ~new_n16595_ & new_n16602_;
  assign new_n16608_ = new_n16524_ | ((~new_n16565_ | ~new_n16567_ | ~new_n16527_) & (new_n13405_ | ~new_n16525_ | new_n16527_));
  assign new_n16609_ = ~new_n13349_ & new_n16524_;
  assign new_n16610_ = new_n7445_ & new_n16611_;
  assign new_n16611_ = ~new_n16640_ & new_n16612_;
  assign new_n16612_ = ~new_n16613_ & ~new_n16639_;
  assign new_n16613_ = new_n16626_ & (~new_n16614_ | (new_n16637_ & new_n16638_ & new_n16634_ & new_n16635_));
  assign new_n16614_ = new_n16615_ & new_n16622_;
  assign new_n16615_ = ~new_n16616_ & ~new_n16618_;
  assign new_n16616_ = ~new_n16617_ & ~\all_features[4431] ;
  assign new_n16617_ = \all_features[4429]  & \all_features[4430]  & (\all_features[4428]  | (\all_features[4426]  & \all_features[4427]  & \all_features[4425] ));
  assign new_n16618_ = ~\all_features[4431]  & (~\all_features[4430]  | ~new_n16619_ | ~new_n16620_ | ~new_n16621_);
  assign new_n16619_ = \all_features[4428]  & \all_features[4429] ;
  assign new_n16620_ = \all_features[4424]  & \all_features[4425] ;
  assign new_n16621_ = \all_features[4426]  & \all_features[4427] ;
  assign new_n16622_ = ~new_n16623_ & ~new_n16624_;
  assign new_n16623_ = ~\all_features[4431]  & (~\all_features[4430]  | (~\all_features[4428]  & ~\all_features[4429]  & ~new_n16621_));
  assign new_n16624_ = ~\all_features[4431]  & (~\all_features[4430]  | (~\all_features[4429]  & (new_n16625_ | ~new_n16621_ | ~\all_features[4428] )));
  assign new_n16625_ = ~\all_features[4424]  & ~\all_features[4425] ;
  assign new_n16626_ = new_n16627_ & new_n16631_;
  assign new_n16627_ = ~new_n16628_ & ~new_n16630_;
  assign new_n16628_ = new_n16629_ & (~\all_features[4429]  | (~\all_features[4428]  & (~\all_features[4427]  | (~\all_features[4426]  & ~\all_features[4425] ))));
  assign new_n16629_ = ~\all_features[4430]  & ~\all_features[4431] ;
  assign new_n16630_ = new_n16629_ & (~\all_features[4427]  | ~new_n16619_ | (~\all_features[4426]  & ~new_n16620_));
  assign new_n16631_ = ~new_n16632_ & ~new_n16633_;
  assign new_n16632_ = ~\all_features[4429]  & new_n16629_ & ((~\all_features[4426]  & new_n16625_) | ~\all_features[4428]  | ~\all_features[4427] );
  assign new_n16633_ = ~\all_features[4431]  & ~\all_features[4430]  & ~\all_features[4429]  & ~\all_features[4427]  & ~\all_features[4428] ;
  assign new_n16634_ = \all_features[4431]  & (\all_features[4430]  | (new_n16619_ & (\all_features[4426]  | \all_features[4427]  | \all_features[4425] )));
  assign new_n16635_ = \all_features[4430]  & \all_features[4431]  & (\all_features[4428]  | \all_features[4429]  | new_n16620_ | ~new_n16636_);
  assign new_n16636_ = ~\all_features[4426]  & ~\all_features[4427] ;
  assign new_n16637_ = \all_features[4431]  & (\all_features[4430]  | (\all_features[4429]  & (\all_features[4428]  | ~new_n16636_ | ~new_n16625_)));
  assign new_n16638_ = \all_features[4431]  & (\all_features[4429]  | \all_features[4430]  | \all_features[4428] );
  assign new_n16639_ = new_n16614_ & new_n16626_;
  assign new_n16640_ = new_n16631_ & (~new_n16627_ | (~new_n16641_ & new_n16622_));
  assign new_n16641_ = new_n16615_ & ((~new_n16642_ & new_n16635_ & new_n16634_) | ~new_n16638_ | ~new_n16637_);
  assign new_n16642_ = \all_features[4431]  & \all_features[4430]  & ~new_n16643_ & \all_features[4429] ;
  assign new_n16643_ = ~\all_features[4427]  & ~\all_features[4428]  & (~\all_features[4426]  | new_n16625_);
  assign new_n16644_ = new_n15365_ & (new_n16649_ | new_n16645_);
  assign new_n16645_ = ~new_n8630_ & ((~new_n12448_ & new_n16648_) ? (~new_n10027_ & new_n16344_) : new_n16646_);
  assign new_n16646_ = ~new_n8482_ & new_n16647_;
  assign new_n16647_ = ~new_n7899_ & ~new_n7902_;
  assign new_n16648_ = new_n9129_ & new_n9131_;
  assign new_n16649_ = new_n8630_ & ((new_n16650_ & new_n16651_) | (~new_n12006_ & ~new_n16651_ & (~new_n16653_ | new_n16652_)));
  assign new_n16650_ = new_n8739_ & (new_n8736_ | new_n8704_);
  assign new_n16651_ = new_n6801_ & ~new_n6770_ & new_n6799_;
  assign new_n16652_ = ~new_n12031_ & ~new_n12035_;
  assign new_n16653_ = ~new_n12007_ & new_n12029_;
  assign new_n16654_ = ~new_n16655_ & new_n16747_;
  assign new_n16655_ = new_n16656_ & new_n16678_ & (~new_n10737_ | ~new_n16746_);
  assign new_n16656_ = (~new_n16104_ | (new_n13807_ ? ~new_n15752_ : ~new_n10701_)) & (~new_n16657_ | new_n16677_ | new_n16104_);
  assign new_n16657_ = new_n16658_ & (new_n11504_ | (~new_n16674_ & ~new_n11512_));
  assign new_n16658_ = ~new_n16670_ & new_n16659_;
  assign new_n16659_ = ~new_n16660_ & ~new_n11498_;
  assign new_n16660_ = new_n16669_ & ~new_n16661_ & new_n11505_;
  assign new_n16661_ = new_n16666_ & (~new_n16667_ | ~new_n16668_ | ~new_n16664_ | ~new_n16662_);
  assign new_n16662_ = \all_features[799]  & (\all_features[798]  | new_n16663_);
  assign new_n16663_ = \all_features[797]  & (\all_features[794]  | \all_features[795]  | \all_features[796]  | ~new_n11513_);
  assign new_n16664_ = \all_features[799]  & ~new_n16665_ & \all_features[798] ;
  assign new_n16665_ = ~\all_features[797]  & ~\all_features[796]  & ~\all_features[795]  & ~new_n11501_ & ~\all_features[794] ;
  assign new_n16666_ = ~new_n11514_ & ~new_n11511_ & ~new_n11509_ & ~new_n11500_;
  assign new_n16667_ = \all_features[799]  & (\all_features[798]  | (new_n11502_ & (\all_features[794]  | \all_features[795]  | \all_features[793] )));
  assign new_n16668_ = \all_features[799]  & (\all_features[797]  | \all_features[798]  | \all_features[796] );
  assign new_n16669_ = ~new_n11512_ & ~new_n11504_;
  assign new_n16670_ = new_n16669_ & (~new_n11505_ | (~new_n16671_ & ~new_n11511_ & ~new_n11514_));
  assign new_n16671_ = ~new_n11500_ & ~new_n11509_ & (~new_n16668_ | new_n16672_ | ~new_n16662_);
  assign new_n16672_ = ~new_n16665_ & new_n16667_ & \all_features[798]  & \all_features[799]  & (~\all_features[797]  | new_n16673_);
  assign new_n16673_ = ~\all_features[795]  & ~\all_features[796]  & (~\all_features[794]  | new_n11513_);
  assign new_n16674_ = ~new_n11508_ & (new_n11506_ | (~new_n11511_ & (new_n11514_ | (~new_n16675_ & ~new_n11509_))));
  assign new_n16675_ = ~new_n11500_ & (~new_n16668_ | (new_n16662_ & (~new_n16667_ | (~new_n16676_ & new_n16664_))));
  assign new_n16676_ = \all_features[798]  & \all_features[799]  & (\all_features[797]  | (\all_features[796]  & (\all_features[795]  | \all_features[794] )));
  assign new_n16677_ = ~new_n15017_ & new_n14989_;
  assign new_n16678_ = new_n16104_ | ((new_n16711_ | ~new_n8165_ | new_n16657_) & (new_n16679_ | ~new_n16677_ | ~new_n16657_));
  assign new_n16679_ = ~new_n16707_ & (~new_n16709_ | ~new_n16680_);
  assign new_n16680_ = new_n16701_ & (new_n16706_ | new_n16681_);
  assign new_n16681_ = ~new_n16697_ & ~new_n16695_ & ~new_n16700_ & (new_n16699_ | (new_n16693_ & new_n16682_));
  assign new_n16682_ = new_n16683_ & (~new_n16688_ | (~new_n16692_ & \all_features[5205]  & \all_features[5206]  & \all_features[5207] ));
  assign new_n16683_ = \all_features[5207]  & (\all_features[5206]  | (~new_n16687_ & new_n16684_));
  assign new_n16684_ = \all_features[5205]  & (\all_features[5204]  | ~new_n16686_ | ~new_n16685_);
  assign new_n16685_ = ~\all_features[5200]  & ~\all_features[5201] ;
  assign new_n16686_ = ~\all_features[5202]  & ~\all_features[5203] ;
  assign new_n16687_ = ~\all_features[5204]  & ~\all_features[5205] ;
  assign new_n16688_ = new_n16689_ & \all_features[5206]  & \all_features[5207]  & (~new_n16686_ | ~new_n16687_ | new_n16691_);
  assign new_n16689_ = \all_features[5207]  & (\all_features[5206]  | (new_n16690_ & (\all_features[5202]  | \all_features[5203]  | \all_features[5201] )));
  assign new_n16690_ = \all_features[5204]  & \all_features[5205] ;
  assign new_n16691_ = \all_features[5200]  & \all_features[5201] ;
  assign new_n16692_ = ~\all_features[5203]  & ~\all_features[5204]  & (~\all_features[5202]  | new_n16685_);
  assign new_n16693_ = \all_features[5207]  & ((~new_n16694_ & \all_features[5206]  & new_n16689_) | (~new_n16687_ & ((~new_n16694_ & new_n16689_) | (~new_n16684_ & ~\all_features[5206] ))));
  assign new_n16694_ = ~\all_features[5205]  & \all_features[5206]  & \all_features[5207]  & (\all_features[5204]  ? new_n16686_ : (new_n16691_ | ~new_n16686_));
  assign new_n16695_ = ~new_n16696_ & ~\all_features[5207] ;
  assign new_n16696_ = \all_features[5205]  & \all_features[5206]  & (\all_features[5204]  | (\all_features[5202]  & \all_features[5203]  & \all_features[5201] ));
  assign new_n16697_ = ~\all_features[5207]  & (~\all_features[5206]  | (~\all_features[5205]  & (new_n16685_ | ~new_n16698_ | ~\all_features[5204] )));
  assign new_n16698_ = \all_features[5202]  & \all_features[5203] ;
  assign new_n16699_ = ~\all_features[5207]  & (~\all_features[5206]  | ~new_n16698_ | ~new_n16691_ | ~new_n16690_);
  assign new_n16700_ = ~\all_features[5207]  & (~\all_features[5206]  | (~new_n16698_ & new_n16687_));
  assign new_n16701_ = ~new_n16704_ & new_n16702_;
  assign new_n16702_ = \all_features[5205]  | \all_features[5206]  | \all_features[5207]  | (\all_features[5204]  & \all_features[5203]  & ~new_n16703_);
  assign new_n16703_ = ~\all_features[5202]  & new_n16685_;
  assign new_n16704_ = ~\all_features[5207]  & ~new_n16705_ & ~\all_features[5206] ;
  assign new_n16705_ = \all_features[5205]  & (\all_features[5204]  | (\all_features[5203]  & (\all_features[5202]  | \all_features[5201] )));
  assign new_n16706_ = ~\all_features[5206]  & ~\all_features[5207]  & (~\all_features[5203]  | ~new_n16690_ | (~\all_features[5202]  & ~new_n16691_));
  assign new_n16707_ = new_n16701_ & new_n16708_ & ~new_n16706_ & ~new_n16695_ & ~new_n16697_;
  assign new_n16708_ = ~new_n16699_ & ~new_n16700_;
  assign new_n16709_ = new_n16702_ & ~new_n16706_ & ~new_n16710_ & ~new_n16704_;
  assign new_n16710_ = ~new_n16695_ & ~new_n16697_ & new_n16708_ & (~new_n16688_ | ~new_n16683_);
  assign new_n16711_ = new_n16744_ & (new_n16712_ | (new_n16735_ & new_n16740_));
  assign new_n16712_ = ~new_n16734_ & ~new_n16733_ & ~new_n16732_ & ~new_n16713_ & ~new_n16730_;
  assign new_n16713_ = new_n16714_ & new_n16719_ & (~new_n16728_ | ~new_n16729_ | ~new_n16725_ | ~new_n16727_);
  assign new_n16714_ = ~new_n16715_ & ~new_n16717_;
  assign new_n16715_ = ~\all_features[2311]  & (~\all_features[2310]  | (~\all_features[2308]  & ~\all_features[2309]  & ~new_n16716_));
  assign new_n16716_ = \all_features[2306]  & \all_features[2307] ;
  assign new_n16717_ = ~\all_features[2311]  & (~\all_features[2310]  | (~\all_features[2309]  & (new_n16718_ | ~\all_features[2308]  | ~new_n16716_)));
  assign new_n16718_ = ~\all_features[2304]  & ~\all_features[2305] ;
  assign new_n16719_ = ~new_n16720_ & ~new_n16722_;
  assign new_n16720_ = ~new_n16721_ & ~\all_features[2311] ;
  assign new_n16721_ = \all_features[2309]  & \all_features[2310]  & (\all_features[2308]  | (\all_features[2306]  & \all_features[2307]  & \all_features[2305] ));
  assign new_n16722_ = ~\all_features[2311]  & (~\all_features[2310]  | ~new_n16723_ | ~new_n16716_ | ~new_n16724_);
  assign new_n16723_ = \all_features[2304]  & \all_features[2305] ;
  assign new_n16724_ = \all_features[2308]  & \all_features[2309] ;
  assign new_n16725_ = \all_features[2311]  & (\all_features[2310]  | (\all_features[2309]  & (\all_features[2308]  | ~new_n16726_ | ~new_n16718_)));
  assign new_n16726_ = ~\all_features[2306]  & ~\all_features[2307] ;
  assign new_n16727_ = \all_features[2311]  & (\all_features[2310]  | (new_n16724_ & (\all_features[2306]  | \all_features[2307]  | \all_features[2305] )));
  assign new_n16728_ = \all_features[2310]  & \all_features[2311]  & (\all_features[2308]  | \all_features[2309]  | new_n16723_ | ~new_n16726_);
  assign new_n16729_ = \all_features[2311]  & (\all_features[2309]  | \all_features[2310]  | \all_features[2308] );
  assign new_n16730_ = ~\all_features[2309]  & new_n16731_ & ((~\all_features[2306]  & new_n16718_) | ~\all_features[2308]  | ~\all_features[2307] );
  assign new_n16731_ = ~\all_features[2310]  & ~\all_features[2311] ;
  assign new_n16732_ = new_n16731_ & (~\all_features[2309]  | (~\all_features[2308]  & (~\all_features[2307]  | (~\all_features[2306]  & ~\all_features[2305] ))));
  assign new_n16733_ = new_n16731_ & (~\all_features[2307]  | ~new_n16724_ | (~\all_features[2306]  & ~new_n16723_));
  assign new_n16734_ = ~\all_features[2311]  & ~\all_features[2310]  & ~\all_features[2309]  & ~\all_features[2307]  & ~\all_features[2308] ;
  assign new_n16735_ = ~new_n16730_ & ~new_n16734_ & (~new_n16739_ | (~new_n16736_ & new_n16714_));
  assign new_n16736_ = new_n16719_ & ((~new_n16737_ & new_n16727_ & new_n16728_) | ~new_n16729_ | ~new_n16725_);
  assign new_n16737_ = \all_features[2311]  & \all_features[2310]  & ~new_n16738_ & \all_features[2309] ;
  assign new_n16738_ = ~\all_features[2307]  & ~\all_features[2308]  & (~\all_features[2306]  | new_n16718_);
  assign new_n16739_ = ~new_n16732_ & ~new_n16733_;
  assign new_n16740_ = ~new_n16741_ & ~new_n16734_;
  assign new_n16741_ = ~new_n16730_ & (new_n16732_ | (~new_n16733_ & (new_n16715_ | (~new_n16717_ & ~new_n16742_))));
  assign new_n16742_ = ~new_n16720_ & (new_n16722_ | (new_n16729_ & (~new_n16725_ | (~new_n16743_ & new_n16727_))));
  assign new_n16743_ = ~\all_features[2309]  & \all_features[2310]  & \all_features[2311]  & (\all_features[2308]  ? new_n16726_ : (new_n16723_ | ~new_n16726_));
  assign new_n16744_ = new_n16739_ & new_n16745_ & ~new_n16717_ & ~new_n16730_ & ~new_n16720_ & ~new_n16715_;
  assign new_n16745_ = ~new_n16722_ & ~new_n16734_;
  assign new_n16746_ = new_n16104_ & ~new_n10701_ & ~new_n13807_;
  assign new_n16747_ = new_n16748_ & new_n16750_;
  assign new_n16748_ = (new_n16749_ | new_n15752_ | ~new_n13807_ | ~new_n16104_) & (new_n8165_ | new_n16657_ | new_n16104_);
  assign new_n16749_ = new_n13269_ & (new_n13245_ | ~new_n13270_);
  assign new_n16750_ = (new_n16104_ | ~new_n16657_ | ~new_n16677_ | ~new_n16679_) & (new_n10737_ | ~new_n16746_);
  assign new_n16751_ = ~new_n16752_ & new_n16768_;
  assign new_n16752_ = (~new_n16760_ & ~new_n16767_ & ~new_n16765_) | (new_n16765_ & (new_n16762_ ? new_n16753_ : ~new_n16756_));
  assign new_n16753_ = new_n14336_ ? new_n9547_ : new_n16754_;
  assign new_n16754_ = new_n16755_ & (~new_n14600_ | ~new_n14579_);
  assign new_n16755_ = ~new_n14607_ & ~new_n14609_;
  assign new_n16756_ = ~new_n16757_ & new_n16758_;
  assign new_n16757_ = ~new_n15530_ & (~new_n15528_ | new_n15497_);
  assign new_n16758_ = ~new_n10833_ & new_n16759_;
  assign new_n16759_ = ~new_n10805_ & ~new_n10830_;
  assign new_n16760_ = new_n11051_ & new_n11027_ & new_n11859_ & new_n16761_;
  assign new_n16761_ = new_n11055_ & new_n11059_;
  assign new_n16762_ = new_n16763_ & new_n16764_;
  assign new_n16763_ = ~new_n15216_ & ~new_n15237_;
  assign new_n16764_ = ~new_n15264_ & ~new_n15244_;
  assign new_n16765_ = new_n12900_ & new_n16766_;
  assign new_n16766_ = ~new_n12872_ & ~new_n12896_;
  assign new_n16767_ = new_n16140_ & (new_n16109_ | new_n16136_ | new_n16133_);
  assign new_n16768_ = ~new_n16770_ & (new_n16765_ ? new_n16769_ : (new_n16767_ | new_n16760_));
  assign new_n16769_ = (new_n14336_ | ~new_n16754_ | ~new_n16762_) & (~new_n16757_ | ~new_n16758_ | new_n16762_);
  assign new_n16770_ = new_n9279_ & new_n16765_ & ~new_n16762_ & ~new_n16758_;
  assign new_n16771_ = ~new_n16892_ & (~new_n16772_ | (new_n16893_ & new_n16894_));
  assign new_n16772_ = new_n16773_ & (~new_n16853_ | (new_n16856_ & new_n16854_) | (~new_n16857_ & ~new_n16854_));
  assign new_n16773_ = ~new_n16774_ & (new_n16849_ | ~new_n16485_ | ~new_n16775_) & (new_n16851_ | ~new_n16848_);
  assign new_n16774_ = ~new_n16775_ & (new_n16812_ ? new_n16814_ : (~new_n16810_ | ~new_n16276_));
  assign new_n16775_ = ~new_n16806_ & new_n16776_;
  assign new_n16776_ = ~new_n16802_ & new_n16777_;
  assign new_n16777_ = ~new_n16778_ & ~new_n16800_;
  assign new_n16778_ = new_n16795_ & ~new_n16799_ & ~new_n16779_ & ~new_n16798_;
  assign new_n16779_ = new_n16780_ & (~new_n16793_ | ~new_n16794_ | ~new_n16790_ | ~new_n16792_);
  assign new_n16780_ = ~new_n16787_ & ~new_n16785_ & ~new_n16781_ & ~new_n16783_;
  assign new_n16781_ = ~\all_features[2543]  & (~\all_features[2542]  | (~\all_features[2540]  & ~\all_features[2541]  & ~new_n16782_));
  assign new_n16782_ = \all_features[2538]  & \all_features[2539] ;
  assign new_n16783_ = ~\all_features[2543]  & (~\all_features[2542]  | (~\all_features[2541]  & (new_n16784_ | ~new_n16782_ | ~\all_features[2540] )));
  assign new_n16784_ = ~\all_features[2536]  & ~\all_features[2537] ;
  assign new_n16785_ = ~new_n16786_ & ~\all_features[2543] ;
  assign new_n16786_ = \all_features[2541]  & \all_features[2542]  & (\all_features[2540]  | (\all_features[2538]  & \all_features[2539]  & \all_features[2537] ));
  assign new_n16787_ = ~\all_features[2543]  & (~\all_features[2542]  | ~new_n16788_ | ~new_n16789_ | ~new_n16782_);
  assign new_n16788_ = \all_features[2536]  & \all_features[2537] ;
  assign new_n16789_ = \all_features[2540]  & \all_features[2541] ;
  assign new_n16790_ = \all_features[2543]  & (\all_features[2542]  | (\all_features[2541]  & (\all_features[2540]  | ~new_n16791_ | ~new_n16784_)));
  assign new_n16791_ = ~\all_features[2538]  & ~\all_features[2539] ;
  assign new_n16792_ = \all_features[2543]  & (\all_features[2542]  | (new_n16789_ & (\all_features[2538]  | \all_features[2539]  | \all_features[2537] )));
  assign new_n16793_ = \all_features[2542]  & \all_features[2543]  & (\all_features[2540]  | \all_features[2541]  | new_n16788_ | ~new_n16791_);
  assign new_n16794_ = \all_features[2543]  & (\all_features[2541]  | \all_features[2542]  | \all_features[2540] );
  assign new_n16795_ = ~new_n16796_ & (\all_features[2539]  | \all_features[2540]  | \all_features[2541]  | \all_features[2542]  | \all_features[2543] );
  assign new_n16796_ = ~\all_features[2541]  & new_n16797_ & ((~\all_features[2538]  & new_n16784_) | ~\all_features[2540]  | ~\all_features[2539] );
  assign new_n16797_ = ~\all_features[2542]  & ~\all_features[2543] ;
  assign new_n16798_ = new_n16797_ & (~\all_features[2541]  | (~\all_features[2540]  & (~\all_features[2539]  | (~\all_features[2538]  & ~\all_features[2537] ))));
  assign new_n16799_ = new_n16797_ & (~\all_features[2539]  | ~new_n16789_ | (~\all_features[2538]  & ~new_n16788_));
  assign new_n16800_ = new_n16801_ & new_n16795_ & ~new_n16798_ & ~new_n16785_;
  assign new_n16801_ = ~new_n16787_ & ~new_n16783_ & ~new_n16799_ & ~new_n16781_;
  assign new_n16802_ = new_n16795_ & (new_n16799_ | new_n16798_ | (~new_n16803_ & ~new_n16781_ & ~new_n16783_));
  assign new_n16803_ = ~new_n16785_ & ~new_n16787_ & (~new_n16794_ | ~new_n16790_ | new_n16804_);
  assign new_n16804_ = new_n16792_ & new_n16793_ & (new_n16805_ | ~\all_features[2541]  | ~\all_features[2542]  | ~\all_features[2543] );
  assign new_n16805_ = ~\all_features[2539]  & ~\all_features[2540]  & (~\all_features[2538]  | new_n16784_);
  assign new_n16806_ = ~new_n16807_ & (\all_features[2539]  | \all_features[2540]  | \all_features[2541]  | \all_features[2542]  | \all_features[2543] );
  assign new_n16807_ = ~new_n16796_ & (new_n16798_ | (~new_n16799_ & (new_n16781_ | (~new_n16808_ & ~new_n16783_))));
  assign new_n16808_ = ~new_n16785_ & (new_n16787_ | (new_n16794_ & (~new_n16790_ | (~new_n16809_ & new_n16792_))));
  assign new_n16809_ = ~\all_features[2541]  & \all_features[2542]  & \all_features[2543]  & (\all_features[2540]  ? new_n16791_ : (new_n16788_ | ~new_n16791_));
  assign new_n16810_ = ~new_n16811_ & new_n8856_;
  assign new_n16811_ = new_n8881_ & new_n8885_;
  assign new_n16812_ = new_n16813_ & ~new_n15823_ & ~new_n15013_;
  assign new_n16813_ = ~new_n14990_ & ~new_n15017_;
  assign new_n16814_ = new_n16815_ & (~new_n16844_ | ~new_n16840_);
  assign new_n16815_ = ~new_n16816_ & ~new_n16838_;
  assign new_n16816_ = new_n16833_ & ~new_n16837_ & ~new_n16817_ & ~new_n16836_;
  assign new_n16817_ = new_n16818_ & (~new_n16831_ | ~new_n16832_ | ~new_n16828_ | ~new_n16830_);
  assign new_n16818_ = ~new_n16827_ & ~new_n16824_ & ~new_n16819_ & ~new_n16822_;
  assign new_n16819_ = ~\all_features[807]  & (~\all_features[806]  | (~\all_features[805]  & (new_n16820_ | ~new_n16821_ | ~\all_features[804] )));
  assign new_n16820_ = ~\all_features[800]  & ~\all_features[801] ;
  assign new_n16821_ = \all_features[802]  & \all_features[803] ;
  assign new_n16822_ = ~new_n16823_ & ~\all_features[807] ;
  assign new_n16823_ = \all_features[805]  & \all_features[806]  & (\all_features[804]  | (\all_features[802]  & \all_features[803]  & \all_features[801] ));
  assign new_n16824_ = ~\all_features[807]  & (~\all_features[806]  | ~new_n16825_ | ~new_n16826_ | ~new_n16821_);
  assign new_n16825_ = \all_features[804]  & \all_features[805] ;
  assign new_n16826_ = \all_features[800]  & \all_features[801] ;
  assign new_n16827_ = ~\all_features[807]  & (~\all_features[806]  | (~\all_features[804]  & ~\all_features[805]  & ~new_n16821_));
  assign new_n16828_ = \all_features[807]  & (\all_features[806]  | (\all_features[805]  & (\all_features[804]  | ~new_n16820_ | ~new_n16829_)));
  assign new_n16829_ = ~\all_features[802]  & ~\all_features[803] ;
  assign new_n16830_ = \all_features[807]  & (\all_features[806]  | (new_n16825_ & (\all_features[802]  | \all_features[803]  | \all_features[801] )));
  assign new_n16831_ = \all_features[806]  & \all_features[807]  & (\all_features[804]  | \all_features[805]  | new_n16826_ | ~new_n16829_);
  assign new_n16832_ = \all_features[807]  & (\all_features[805]  | \all_features[806]  | \all_features[804] );
  assign new_n16833_ = ~new_n16834_ & (\all_features[803]  | \all_features[804]  | \all_features[805]  | \all_features[806]  | \all_features[807] );
  assign new_n16834_ = ~\all_features[805]  & new_n16835_ & ((~\all_features[802]  & new_n16820_) | ~\all_features[804]  | ~\all_features[803] );
  assign new_n16835_ = ~\all_features[806]  & ~\all_features[807] ;
  assign new_n16836_ = new_n16835_ & (~\all_features[805]  | (~\all_features[804]  & (~\all_features[803]  | (~\all_features[802]  & ~\all_features[801] ))));
  assign new_n16837_ = new_n16835_ & (~\all_features[803]  | ~new_n16825_ | (~\all_features[802]  & ~new_n16826_));
  assign new_n16838_ = new_n16839_ & new_n16833_ & ~new_n16822_ & ~new_n16836_;
  assign new_n16839_ = ~new_n16837_ & ~new_n16827_ & ~new_n16819_ & ~new_n16824_;
  assign new_n16840_ = new_n16833_ & (new_n16837_ | new_n16836_ | (~new_n16819_ & ~new_n16827_ & ~new_n16841_));
  assign new_n16841_ = ~new_n16824_ & ~new_n16822_ & (~new_n16832_ | ~new_n16828_ | new_n16842_);
  assign new_n16842_ = new_n16830_ & new_n16831_ & (new_n16843_ | ~\all_features[805]  | ~\all_features[806]  | ~\all_features[807] );
  assign new_n16843_ = ~\all_features[803]  & ~\all_features[804]  & (~\all_features[802]  | new_n16820_);
  assign new_n16844_ = ~new_n16845_ & (\all_features[803]  | \all_features[804]  | \all_features[805]  | \all_features[806]  | \all_features[807] );
  assign new_n16845_ = ~new_n16834_ & (new_n16836_ | (~new_n16837_ & (new_n16827_ | (~new_n16819_ & ~new_n16846_))));
  assign new_n16846_ = ~new_n16822_ & (new_n16824_ | (new_n16832_ & (~new_n16828_ | (~new_n16847_ & new_n16830_))));
  assign new_n16847_ = ~\all_features[805]  & \all_features[806]  & \all_features[807]  & (\all_features[804]  ? new_n16829_ : (new_n16826_ | ~new_n16829_));
  assign new_n16848_ = new_n16812_ & ~new_n16775_ & ~new_n16814_;
  assign new_n16849_ = new_n15152_ & new_n16850_;
  assign new_n16850_ = ~new_n11598_ & new_n11904_;
  assign new_n16851_ = ~new_n16852_ & new_n6495_;
  assign new_n16852_ = ~new_n6491_ & ~new_n6484_;
  assign new_n16853_ = ~new_n16485_ & new_n16775_;
  assign new_n16854_ = ~new_n9579_ & new_n16855_;
  assign new_n16855_ = ~new_n9572_ & ~new_n9581_;
  assign new_n16856_ = ~new_n9836_ & new_n10637_;
  assign new_n16857_ = ~new_n16890_ & ~new_n16879_ & ~new_n16887_ & (new_n16885_ | (~new_n16884_ & ~new_n16858_));
  assign new_n16858_ = ~new_n16872_ & (new_n16874_ | (~new_n16875_ & (new_n16876_ | (~new_n16859_ & ~new_n16877_))));
  assign new_n16859_ = ~new_n16866_ & (~new_n16870_ | (new_n16860_ & (~new_n16869_ | (~new_n16871_ & new_n16863_))));
  assign new_n16860_ = \all_features[5423]  & (\all_features[5422]  | new_n16861_);
  assign new_n16861_ = \all_features[5421]  & (\all_features[5418]  | \all_features[5419]  | \all_features[5420]  | ~new_n16862_);
  assign new_n16862_ = ~\all_features[5416]  & ~\all_features[5417] ;
  assign new_n16863_ = \all_features[5423]  & ~new_n16864_ & \all_features[5422] ;
  assign new_n16864_ = ~\all_features[5421]  & ~\all_features[5420]  & ~\all_features[5419]  & ~new_n16865_ & ~\all_features[5418] ;
  assign new_n16865_ = \all_features[5416]  & \all_features[5417] ;
  assign new_n16866_ = ~\all_features[5423]  & (~\all_features[5422]  | ~new_n16865_ | ~new_n16867_ | ~new_n16868_);
  assign new_n16867_ = \all_features[5420]  & \all_features[5421] ;
  assign new_n16868_ = \all_features[5418]  & \all_features[5419] ;
  assign new_n16869_ = \all_features[5423]  & (\all_features[5422]  | (new_n16867_ & (\all_features[5418]  | \all_features[5419]  | \all_features[5417] )));
  assign new_n16870_ = \all_features[5423]  & (\all_features[5421]  | \all_features[5422]  | \all_features[5420] );
  assign new_n16871_ = \all_features[5422]  & \all_features[5423]  & (\all_features[5421]  | (\all_features[5420]  & (\all_features[5419]  | \all_features[5418] )));
  assign new_n16872_ = new_n16873_ & (~\all_features[5421]  | (~\all_features[5420]  & (~\all_features[5419]  | (~\all_features[5418]  & ~\all_features[5417] ))));
  assign new_n16873_ = ~\all_features[5422]  & ~\all_features[5423] ;
  assign new_n16874_ = new_n16873_ & (~\all_features[5419]  | ~new_n16867_ | (~\all_features[5418]  & ~new_n16865_));
  assign new_n16875_ = ~\all_features[5423]  & (~\all_features[5422]  | (~\all_features[5420]  & ~\all_features[5421]  & ~new_n16868_));
  assign new_n16876_ = ~\all_features[5423]  & (~\all_features[5422]  | (~\all_features[5421]  & (new_n16862_ | ~new_n16868_ | ~\all_features[5420] )));
  assign new_n16877_ = ~new_n16878_ & ~\all_features[5423] ;
  assign new_n16878_ = \all_features[5421]  & \all_features[5422]  & (\all_features[5420]  | (\all_features[5418]  & \all_features[5419]  & \all_features[5417] ));
  assign new_n16879_ = new_n16883_ & (~new_n16886_ | (~new_n16880_ & ~new_n16875_ & ~new_n16876_));
  assign new_n16880_ = ~new_n16866_ & ~new_n16877_ & (~new_n16870_ | new_n16881_ | ~new_n16860_);
  assign new_n16881_ = ~new_n16864_ & new_n16869_ & \all_features[5422]  & \all_features[5423]  & (~\all_features[5421]  | new_n16882_);
  assign new_n16882_ = ~\all_features[5419]  & ~\all_features[5420]  & (~\all_features[5418]  | new_n16862_);
  assign new_n16883_ = ~new_n16884_ & ~new_n16885_;
  assign new_n16884_ = ~\all_features[5421]  & new_n16873_ & ((~\all_features[5418]  & new_n16862_) | ~\all_features[5420]  | ~\all_features[5419] );
  assign new_n16885_ = ~\all_features[5423]  & ~\all_features[5422]  & ~\all_features[5421]  & ~\all_features[5419]  & ~\all_features[5420] ;
  assign new_n16886_ = ~new_n16872_ & ~new_n16874_;
  assign new_n16887_ = new_n16886_ & ~new_n16888_ & new_n16883_;
  assign new_n16888_ = new_n16889_ & (~new_n16869_ | ~new_n16870_ | ~new_n16863_ | ~new_n16860_);
  assign new_n16889_ = ~new_n16866_ & ~new_n16877_ & ~new_n16875_ & ~new_n16876_;
  assign new_n16890_ = new_n16891_ & new_n16883_ & ~new_n16872_ & ~new_n16877_;
  assign new_n16891_ = ~new_n16866_ & ~new_n16876_ & ~new_n16874_ & ~new_n16875_;
  assign new_n16892_ = new_n16856_ & new_n16853_ & new_n16854_;
  assign new_n16893_ = new_n16848_ & new_n16851_;
  assign new_n16894_ = ~new_n16775_ | ((~new_n16849_ | ~new_n16485_) & (new_n16854_ | new_n16857_ | new_n16485_));
  assign new_n16895_ = ~new_n16896_ & new_n16950_;
  assign new_n16896_ = ~new_n16941_ & ~new_n16947_ & new_n16897_ & (~new_n16944_ | (~new_n16945_ & ~new_n16949_));
  assign new_n16897_ = ~new_n16898_ & (new_n11095_ | ~new_n16907_ | ~new_n16910_);
  assign new_n16898_ = new_n12117_ & new_n14469_ & ~new_n16899_ & new_n15671_;
  assign new_n16899_ = new_n16900_ & new_n16906_;
  assign new_n16900_ = ~new_n7805_ & ~new_n16901_;
  assign new_n16901_ = ~new_n7811_ & (new_n7807_ | (~new_n7826_ & (new_n7825_ | (~new_n7821_ & ~new_n16902_))));
  assign new_n16902_ = ~new_n7823_ & (new_n7827_ | (~new_n7829_ & (~new_n16905_ | new_n16903_)));
  assign new_n16903_ = \all_features[3447]  & ((~new_n16904_ & ~\all_features[3445]  & \all_features[3446] ) | (~new_n7816_ & (\all_features[3446]  | (~new_n7814_ & \all_features[3445] ))));
  assign new_n16904_ = (~\all_features[3442]  & ~\all_features[3443]  & ~\all_features[3444]  & (~\all_features[3441]  | ~\all_features[3440] )) | (\all_features[3444]  & (\all_features[3442]  | \all_features[3443] ));
  assign new_n16905_ = \all_features[3447]  & (\all_features[3445]  | \all_features[3446]  | \all_features[3444] );
  assign new_n16906_ = ~new_n7830_ & ~new_n7832_;
  assign new_n16907_ = ~new_n12117_ & ~new_n16908_;
  assign new_n16908_ = ~new_n13209_ & new_n16909_;
  assign new_n16909_ = new_n13238_ & new_n13242_;
  assign new_n16910_ = ~new_n16911_ & new_n16933_ & (new_n16940_ | new_n16916_ | new_n16918_ | ~new_n16938_);
  assign new_n16911_ = ~new_n16926_ & (new_n16928_ | (~new_n16930_ & (new_n16931_ | (~new_n16912_ & ~new_n16932_))));
  assign new_n16912_ = ~new_n16916_ & (new_n16918_ | (new_n16925_ & (~new_n16913_ | (~new_n16922_ & new_n16924_))));
  assign new_n16913_ = \all_features[1167]  & (\all_features[1166]  | new_n16914_);
  assign new_n16914_ = \all_features[1165]  & (\all_features[1162]  | \all_features[1163]  | \all_features[1164]  | ~new_n16915_);
  assign new_n16915_ = ~\all_features[1160]  & ~\all_features[1161] ;
  assign new_n16916_ = ~new_n16917_ & ~\all_features[1167] ;
  assign new_n16917_ = \all_features[1165]  & \all_features[1166]  & (\all_features[1164]  | (\all_features[1162]  & \all_features[1163]  & \all_features[1161] ));
  assign new_n16918_ = ~\all_features[1167]  & (~\all_features[1166]  | ~new_n16919_ | ~new_n16920_ | ~new_n16921_);
  assign new_n16919_ = \all_features[1160]  & \all_features[1161] ;
  assign new_n16920_ = \all_features[1164]  & \all_features[1165] ;
  assign new_n16921_ = \all_features[1162]  & \all_features[1163] ;
  assign new_n16922_ = ~\all_features[1165]  & new_n16923_ & ((~\all_features[1164]  & (new_n16919_ | \all_features[1162]  | \all_features[1163] )) | (~\all_features[1162]  & ~\all_features[1163]  & \all_features[1164] ));
  assign new_n16923_ = \all_features[1166]  & \all_features[1167] ;
  assign new_n16924_ = \all_features[1167]  & (\all_features[1166]  | (new_n16920_ & (\all_features[1162]  | \all_features[1163]  | \all_features[1161] )));
  assign new_n16925_ = \all_features[1167]  & (\all_features[1165]  | \all_features[1166]  | \all_features[1164] );
  assign new_n16926_ = new_n16927_ & ((~\all_features[1162]  & new_n16915_) | ~\all_features[1164]  | ~\all_features[1163] );
  assign new_n16927_ = ~\all_features[1167]  & ~\all_features[1165]  & ~\all_features[1166] ;
  assign new_n16928_ = ~\all_features[1167]  & ~new_n16929_ & ~\all_features[1166] ;
  assign new_n16929_ = \all_features[1165]  & (\all_features[1164]  | (\all_features[1163]  & (\all_features[1162]  | \all_features[1161] )));
  assign new_n16930_ = ~\all_features[1166]  & ~\all_features[1167]  & (~\all_features[1163]  | ~new_n16920_ | (~\all_features[1162]  & ~new_n16919_));
  assign new_n16931_ = ~\all_features[1167]  & (~\all_features[1166]  | (~\all_features[1164]  & ~\all_features[1165]  & ~new_n16921_));
  assign new_n16932_ = ~\all_features[1167]  & (~\all_features[1166]  | (~\all_features[1165]  & (new_n16915_ | ~new_n16921_ | ~\all_features[1164] )));
  assign new_n16933_ = ~new_n16928_ & ~new_n16916_ & new_n16939_ & new_n16938_ & (new_n16918_ | new_n16934_);
  assign new_n16934_ = new_n16925_ & ~new_n16935_ & new_n16913_;
  assign new_n16935_ = new_n16924_ & new_n16936_ & (~\all_features[1165]  | ~new_n16923_ | new_n16937_);
  assign new_n16936_ = new_n16923_ & (new_n16919_ | \all_features[1162]  | \all_features[1163]  | \all_features[1164]  | \all_features[1165] );
  assign new_n16937_ = ~\all_features[1163]  & ~\all_features[1164]  & (~\all_features[1162]  | new_n16915_);
  assign new_n16938_ = ~new_n16931_ & ~new_n16932_;
  assign new_n16939_ = ~new_n16926_ & ~new_n16930_ & ~new_n16918_ & (\all_features[1164]  | \all_features[1163]  | ~new_n16927_);
  assign new_n16940_ = new_n16925_ & new_n16924_ & new_n16913_ & new_n16936_;
  assign new_n16941_ = new_n16942_ & new_n15039_;
  assign new_n16942_ = new_n12117_ & ~new_n14469_ & ~new_n16943_;
  assign new_n16943_ = new_n16660_ & new_n11498_;
  assign new_n16944_ = ~new_n12117_ & new_n16908_;
  assign new_n16945_ = new_n14293_ & new_n16946_;
  assign new_n16946_ = new_n14545_ & new_n6674_ & new_n14541_;
  assign new_n16947_ = new_n16948_ & new_n16943_ & new_n12117_ & ~new_n14469_ & ~new_n14277_;
  assign new_n16948_ = ~new_n12718_ & ~new_n12721_;
  assign new_n16949_ = ~new_n16946_ & new_n13800_;
  assign new_n16950_ = new_n16951_ & (~new_n16907_ | (~new_n11095_ & new_n16910_));
  assign new_n16951_ = ~new_n16952_ & (new_n15039_ | ~new_n16942_) & (new_n16949_ | new_n16945_ | ~new_n16944_);
  assign new_n16952_ = new_n14469_ & new_n12117_ & (new_n16899_ ? ~new_n15595_ : ~new_n15671_);
  assign new_n16953_ = ~new_n16954_ & new_n17008_;
  assign new_n16954_ = ~new_n16994_ & (new_n16955_ | new_n16997_) & (new_n16956_ | new_n16765_ | ~new_n17000_ | ~new_n16997_);
  assign new_n16955_ = (new_n16957_ | ~new_n13807_ | ~new_n16956_) & (new_n14290_ | ~new_n16963_ | new_n16956_);
  assign new_n16956_ = ~new_n13707_ & ~new_n13676_ & ~new_n13703_;
  assign new_n16957_ = new_n16958_ & ~new_n16054_ & ~new_n16959_;
  assign new_n16958_ = ~new_n16030_ & ~new_n16058_;
  assign new_n16959_ = ~new_n16036_ & (new_n16033_ | (~new_n16037_ & ~new_n16960_));
  assign new_n16960_ = ~new_n16038_ & (new_n16051_ | (~new_n16046_ & (new_n16048_ | (~new_n16050_ & ~new_n16961_))));
  assign new_n16961_ = new_n16044_ & (~new_n16042_ | (new_n16053_ & (new_n16962_ | ~new_n16052_)));
  assign new_n16962_ = \all_features[2550]  & \all_features[2551]  & (\all_features[2549]  | (~new_n16043_ & \all_features[2548] ));
  assign new_n16963_ = ~new_n16964_ & new_n16986_ & (new_n16993_ | new_n16969_ | new_n16971_ | ~new_n16991_);
  assign new_n16964_ = ~new_n16979_ & (new_n16981_ | (~new_n16983_ & (new_n16984_ | (~new_n16965_ & ~new_n16985_))));
  assign new_n16965_ = ~new_n16969_ & (new_n16971_ | (new_n16978_ & (~new_n16966_ | (~new_n16975_ & new_n16977_))));
  assign new_n16966_ = \all_features[4967]  & (\all_features[4966]  | new_n16967_);
  assign new_n16967_ = \all_features[4965]  & (\all_features[4962]  | \all_features[4963]  | \all_features[4964]  | ~new_n16968_);
  assign new_n16968_ = ~\all_features[4960]  & ~\all_features[4961] ;
  assign new_n16969_ = ~new_n16970_ & ~\all_features[4967] ;
  assign new_n16970_ = \all_features[4965]  & \all_features[4966]  & (\all_features[4964]  | (\all_features[4962]  & \all_features[4963]  & \all_features[4961] ));
  assign new_n16971_ = ~\all_features[4967]  & (~\all_features[4966]  | ~new_n16972_ | ~new_n16973_ | ~new_n16974_);
  assign new_n16972_ = \all_features[4960]  & \all_features[4961] ;
  assign new_n16973_ = \all_features[4964]  & \all_features[4965] ;
  assign new_n16974_ = \all_features[4962]  & \all_features[4963] ;
  assign new_n16975_ = ~\all_features[4965]  & new_n16976_ & ((~\all_features[4964]  & (new_n16972_ | \all_features[4962]  | \all_features[4963] )) | (~\all_features[4962]  & ~\all_features[4963]  & \all_features[4964] ));
  assign new_n16976_ = \all_features[4966]  & \all_features[4967] ;
  assign new_n16977_ = \all_features[4967]  & (\all_features[4966]  | (new_n16973_ & (\all_features[4962]  | \all_features[4963]  | \all_features[4961] )));
  assign new_n16978_ = \all_features[4967]  & (\all_features[4965]  | \all_features[4966]  | \all_features[4964] );
  assign new_n16979_ = new_n16980_ & ((~\all_features[4962]  & new_n16968_) | ~\all_features[4964]  | ~\all_features[4963] );
  assign new_n16980_ = ~\all_features[4967]  & ~\all_features[4965]  & ~\all_features[4966] ;
  assign new_n16981_ = ~\all_features[4967]  & ~new_n16982_ & ~\all_features[4966] ;
  assign new_n16982_ = \all_features[4965]  & (\all_features[4964]  | (\all_features[4963]  & (\all_features[4962]  | \all_features[4961] )));
  assign new_n16983_ = ~\all_features[4966]  & ~\all_features[4967]  & (~\all_features[4963]  | ~new_n16973_ | (~\all_features[4962]  & ~new_n16972_));
  assign new_n16984_ = ~\all_features[4967]  & (~\all_features[4966]  | (~\all_features[4964]  & ~\all_features[4965]  & ~new_n16974_));
  assign new_n16985_ = ~\all_features[4967]  & (~\all_features[4966]  | (~\all_features[4965]  & (new_n16968_ | ~new_n16974_ | ~\all_features[4964] )));
  assign new_n16986_ = ~new_n16981_ & ~new_n16969_ & new_n16992_ & new_n16991_ & (new_n16971_ | new_n16987_);
  assign new_n16987_ = new_n16978_ & ~new_n16988_ & new_n16966_;
  assign new_n16988_ = new_n16977_ & new_n16989_ & (~\all_features[4965]  | ~new_n16976_ | new_n16990_);
  assign new_n16989_ = new_n16976_ & (new_n16972_ | \all_features[4962]  | \all_features[4963]  | \all_features[4964]  | \all_features[4965] );
  assign new_n16990_ = ~\all_features[4963]  & ~\all_features[4964]  & (~\all_features[4962]  | new_n16968_);
  assign new_n16991_ = ~new_n16984_ & ~new_n16985_;
  assign new_n16992_ = ~new_n16979_ & ~new_n16983_ & ~new_n16971_ & (\all_features[4964]  | \all_features[4963]  | ~new_n16980_);
  assign new_n16993_ = new_n16978_ & new_n16977_ & new_n16966_ & new_n16989_;
  assign new_n16994_ = new_n16956_ & new_n16957_ & (new_n16996_ | new_n16995_);
  assign new_n16995_ = new_n14211_ & new_n16350_;
  assign new_n16996_ = ~new_n7375_ & new_n7591_;
  assign new_n16997_ = new_n16998_ & new_n16999_;
  assign new_n16998_ = new_n6640_ & new_n6662_;
  assign new_n16999_ = new_n6666_ & new_n6670_;
  assign new_n17000_ = new_n13708_ & new_n17001_;
  assign new_n17001_ = ~new_n13732_ & (~new_n17007_ | (~new_n13726_ & (new_n13721_ | new_n17005_ | ~new_n17002_)));
  assign new_n17002_ = ~new_n13723_ & ~new_n13725_ & (~new_n13716_ | (~new_n17003_ & new_n13710_));
  assign new_n17003_ = \all_features[4671]  & \all_features[4670]  & ~new_n17004_ & \all_features[4669] ;
  assign new_n17004_ = ~\all_features[4667]  & ~\all_features[4668]  & (~\all_features[4666]  | new_n13718_);
  assign new_n17005_ = ~new_n13723_ & (new_n13725_ | (new_n13719_ & (~new_n13717_ | (~new_n17006_ & new_n13714_))));
  assign new_n17006_ = ~\all_features[4669]  & \all_features[4670]  & \all_features[4671]  & (\all_features[4668]  ? new_n13712_ : (new_n13713_ | ~new_n13712_));
  assign new_n17007_ = ~new_n13731_ & ~new_n13728_ & ~new_n13730_;
  assign new_n17008_ = new_n17009_ & (new_n17011_ | new_n16956_) & (new_n16957_ | new_n17012_ | ~new_n16997_ | ~new_n16956_);
  assign new_n17009_ = new_n16956_ ? new_n17010_ : ((new_n16064_ | ~new_n16765_ | ~new_n16997_) & (~new_n14290_ | new_n16997_));
  assign new_n17010_ = (new_n13807_ | new_n16997_ | new_n16957_) & (new_n16995_ | new_n16996_ | ~new_n16957_);
  assign new_n17011_ = (new_n14290_ | new_n16963_ | new_n16997_) & (new_n16765_ | new_n17000_ | ~new_n16997_);
  assign new_n17012_ = new_n17013_ & new_n11901_;
  assign new_n17013_ = new_n6535_ & new_n6556_;
  assign \o[8]  = ~new_n17015_ ^ new_n17016_;
  assign new_n17015_ = (new_n16895_ & new_n16953_) | (~new_n13664_ & (new_n16895_ | new_n16953_));
  assign new_n17016_ = new_n17017_ ? (~new_n17018_ ^ new_n17070_) : (new_n17018_ ^ new_n17070_);
  assign new_n17017_ = (~new_n16324_ & new_n16771_) | (~new_n13665_ & (~new_n16324_ | new_n16771_));
  assign new_n17018_ = new_n17019_ ? (new_n17020_ ^ new_n17057_) : (~new_n17020_ ^ new_n17057_);
  assign new_n17019_ = (~new_n15400_ & new_n16149_) | (~new_n13666_ & (~new_n15400_ | new_n16149_));
  assign new_n17020_ = new_n17021_ ? (new_n17034_ ^ new_n17035_) : (~new_n17034_ ^ new_n17035_);
  assign new_n17021_ = new_n17022_ ? (~new_n17032_ ^ new_n17033_) : (new_n17032_ ^ new_n17033_);
  assign new_n17022_ = new_n17023_ ? (new_n17027_ ^ new_n17028_) : (~new_n17027_ ^ new_n17028_);
  assign new_n17023_ = new_n17024_ ? (new_n17025_ ^ new_n17026_) : (~new_n17025_ ^ new_n17026_);
  assign new_n17024_ = new_n16150_ & new_n16320_;
  assign new_n17025_ = new_n16521_ & new_n16572_;
  assign new_n17026_ = new_n15150_ & new_n15209_;
  assign new_n17027_ = (new_n15544_ & new_n15666_) | (new_n15403_ & (new_n15544_ | new_n15666_));
  assign new_n17028_ = new_n17029_ ? (~new_n17030_ ^ new_n16107_) : (new_n17030_ ^ new_n16107_);
  assign new_n17029_ = new_n15909_ & new_n16059_;
  assign new_n17030_ = new_n15026_ & new_n15111_;
  assign new_n17032_ = (~new_n15708_ & new_n15907_) | (~new_n15402_ & (~new_n15708_ | new_n15907_));
  assign new_n17033_ = (new_n14613_ & new_n15211_) | (~new_n14870_ & (new_n14613_ | new_n15211_));
  assign new_n17034_ = (~new_n14869_ & ~new_n15350_) | (~new_n13667_ & (~new_n14869_ | ~new_n15350_));
  assign new_n17035_ = new_n17036_ ? (new_n17043_ ^ new_n17044_) : (~new_n17043_ ^ new_n17044_);
  assign new_n17036_ = new_n17037_ ? (~new_n17038_ ^ new_n17039_) : (new_n17038_ ^ new_n17039_);
  assign new_n17037_ = (new_n13884_ & new_n14081_) | (new_n13669_ & (new_n13884_ | new_n14081_));
  assign new_n17038_ = (new_n15025_ & new_n15149_) | (new_n14871_ & (new_n15025_ | new_n15149_));
  assign new_n17039_ = new_n17040_ ? (new_n17041_ ^ new_n17042_) : (~new_n17041_ ^ new_n17042_);
  assign new_n17040_ = new_n14872_ & new_n15019_;
  assign new_n17041_ = new_n16655_ & new_n16747_;
  assign new_n17042_ = new_n16752_ & new_n16768_;
  assign new_n17043_ = (~new_n14284_ & new_n14613_) | (~new_n13668_ & (~new_n14284_ | new_n14613_));
  assign new_n17044_ = new_n17045_ ? (~new_n17051_ ^ new_n17052_) : (new_n17051_ ^ new_n17052_);
  assign new_n17045_ = new_n17046_ ? (new_n17047_ ^ new_n17050_) : (~new_n17047_ ^ new_n17050_);
  assign new_n17046_ = new_n13670_ & new_n13847_;
  assign new_n17047_ = ~new_n17049_ & new_n17048_;
  assign new_n17048_ = ~new_n16892_ & new_n16772_;
  assign new_n17049_ = ~new_n16893_ & new_n16894_;
  assign new_n17050_ = new_n16954_ & new_n17008_;
  assign new_n17051_ = ~new_n14285_ & ~new_n14432_;
  assign new_n17052_ = new_n17053_ ? (new_n17054_ ^ new_n17055_) : (~new_n17054_ ^ new_n17055_);
  assign new_n17053_ = new_n14286_ & new_n14430_ & (new_n14429_ | ~new_n14428_ | ~new_n14427_);
  assign new_n17054_ = new_n14433_ & new_n14611_;
  assign new_n17055_ = new_n17056_ & new_n16896_ & new_n16950_;
  assign new_n17056_ = new_n15595_ & new_n16899_ & new_n12117_ & new_n14469_;
  assign new_n17057_ = new_n17058_ ? (~new_n17059_ ^ new_n17060_) : (new_n17059_ ^ new_n17060_);
  assign new_n17058_ = (new_n15908_ & new_n16062_) | (~new_n15401_ & (new_n15908_ | new_n16062_));
  assign new_n17059_ = (new_n16520_ & new_n16644_) | (~new_n16326_ & (new_n16520_ | new_n16644_));
  assign new_n17060_ = new_n17061_ ? (~new_n17062_ ^ new_n17069_) : (new_n17062_ ^ new_n17069_);
  assign new_n17061_ = (~new_n16451_ & new_n15907_) | (~new_n16327_ & (~new_n16451_ | new_n15907_));
  assign new_n17062_ = new_n17063_ ? (~new_n17064_ ^ new_n17068_) : (new_n17064_ ^ new_n17068_);
  assign new_n17063_ = (new_n16372_ & new_n16373_) | (new_n16328_ & (new_n16372_ | new_n16373_));
  assign new_n17064_ = new_n17065_ ? (new_n17066_ ^ new_n17067_) : (~new_n17066_ ^ new_n17067_);
  assign new_n17065_ = new_n16329_ & new_n16368_;
  assign new_n17066_ = new_n15545_ & new_n15629_;
  assign new_n17067_ = new_n15710_ & new_n15758_;
  assign new_n17068_ = (new_n15759_ & new_n15865_) | (new_n15709_ & (new_n15759_ | new_n15865_));
  assign new_n17069_ = new_n15212_ & new_n15349_;
  assign new_n17070_ = (new_n16654_ & new_n16751_) | (~new_n16325_ & (new_n16654_ | new_n16751_));
  assign \o[9]  = ~new_n17072_ ^ new_n17073_;
  assign new_n17072_ = ~new_n17016_ & new_n17015_;
  assign new_n17073_ = new_n17074_ ^ new_n17075_;
  assign new_n17074_ = (~new_n17018_ & new_n17070_) | (new_n17017_ & (~new_n17018_ | new_n17070_));
  assign new_n17075_ = new_n17076_ ? (~new_n17077_ ^ new_n17104_) : (new_n17077_ ^ new_n17104_);
  assign new_n17076_ = (~new_n17020_ & ~new_n17057_) | (new_n17019_ & (~new_n17020_ | ~new_n17057_));
  assign new_n17077_ = new_n17078_ ? (new_n17086_ ^ new_n17087_) : (~new_n17086_ ^ new_n17087_);
  assign new_n17078_ = new_n17079_ ? (~new_n17080_ ^ new_n17081_) : (new_n17080_ ^ new_n17081_);
  assign new_n17079_ = (new_n17032_ & new_n17033_) | (~new_n17022_ & (new_n17032_ | new_n17033_));
  assign new_n17080_ = (~new_n17062_ & new_n17069_) | (new_n17061_ & (~new_n17062_ | new_n17069_));
  assign new_n17081_ = ~new_n17082_ ^ new_n17083_;
  assign new_n17082_ = (~new_n17064_ & new_n17068_) | (new_n17063_ & (~new_n17064_ | new_n17068_));
  assign new_n17083_ = new_n17084_ ^ new_n17085_;
  assign new_n17084_ = (new_n17066_ & new_n17067_) | (new_n17065_ & (new_n17066_ | new_n17067_));
  assign new_n17085_ = (~new_n16107_ & new_n17030_) | (new_n17029_ & (~new_n16107_ | new_n17030_));
  assign new_n17086_ = (~new_n17035_ & new_n17034_) | (~new_n17021_ & (~new_n17035_ | new_n17034_));
  assign new_n17087_ = new_n17088_ ? (new_n17092_ ^ new_n17093_) : (~new_n17092_ ^ new_n17093_);
  assign new_n17088_ = new_n17089_ ? (new_n17090_ ^ new_n17091_) : (~new_n17090_ ^ new_n17091_);
  assign new_n17089_ = (~new_n17028_ & new_n17027_) | (~new_n17023_ & (~new_n17028_ | new_n17027_));
  assign new_n17090_ = (~new_n17039_ & new_n17038_) | (new_n17037_ & (~new_n17039_ | new_n17038_));
  assign new_n17091_ = (new_n17025_ & new_n17026_) | (new_n17024_ & (new_n17025_ | new_n17026_));
  assign new_n17092_ = (~new_n17044_ & new_n17043_) | (~new_n17036_ & (~new_n17044_ | new_n17043_));
  assign new_n17093_ = new_n17094_ ? (new_n17097_ ^ new_n17098_) : (~new_n17097_ ^ new_n17098_);
  assign new_n17094_ = ~new_n17095_ ^ new_n17096_;
  assign new_n17095_ = (new_n17047_ & new_n17050_) | (new_n17046_ & (new_n17047_ | new_n17050_));
  assign new_n17096_ = (new_n17041_ & new_n17042_) | (new_n17040_ & (new_n17041_ | new_n17042_));
  assign new_n17097_ = (~new_n17051_ & ~new_n17052_) | (~new_n17045_ & (~new_n17051_ | ~new_n17052_));
  assign new_n17098_ = new_n17099_ ^ new_n17100_;
  assign new_n17099_ = (new_n17054_ & new_n17055_) | (new_n17053_ & (new_n17054_ | new_n17055_));
  assign new_n17100_ = new_n17101_ ? (new_n17102_ ^ new_n17103_) : (~new_n17102_ ^ new_n17103_);
  assign new_n17101_ = new_n17048_ & new_n17049_;
  assign new_n17102_ = new_n14430_ & new_n14286_ & ~new_n14429_ & new_n14427_;
  assign new_n17103_ = new_n16896_ & ~new_n17056_ & new_n16950_;
  assign new_n17104_ = (~new_n17060_ & new_n17059_) | (new_n17058_ & (~new_n17060_ | new_n17059_));
  assign \o[10]  = ((new_n17106_ | new_n17107_) & (new_n17108_ ^ new_n17109_)) | (~new_n17106_ & ~new_n17107_ & (~new_n17108_ ^ new_n17109_));
  assign new_n17106_ = ~new_n17073_ & new_n17072_;
  assign new_n17107_ = ~new_n17075_ & new_n17074_;
  assign new_n17108_ = (~new_n17077_ & new_n17104_) | (new_n17076_ & (~new_n17077_ | new_n17104_));
  assign new_n17109_ = new_n17110_ ? (~new_n17111_ ^ new_n17123_) : (new_n17111_ ^ new_n17123_);
  assign new_n17110_ = (~new_n17087_ & new_n17086_) | (~new_n17078_ & (~new_n17087_ | new_n17086_));
  assign new_n17111_ = new_n17112_ ? (new_n17116_ ^ new_n17117_) : (~new_n17116_ ^ new_n17117_);
  assign new_n17112_ = new_n17113_ ? (new_n17114_ ^ new_n17115_) : (~new_n17114_ ^ new_n17115_);
  assign new_n17113_ = (new_n17090_ & new_n17091_) | (new_n17089_ & (new_n17090_ | new_n17091_));
  assign new_n17114_ = new_n17082_ & new_n17083_;
  assign new_n17115_ = new_n17084_ & new_n17085_;
  assign new_n17116_ = (~new_n17093_ & new_n17092_) | (~new_n17088_ & (~new_n17093_ | new_n17092_));
  assign new_n17117_ = new_n17118_ ? (~new_n17119_ ^ new_n17120_) : (new_n17119_ ^ new_n17120_);
  assign new_n17118_ = (~new_n17098_ & new_n17097_) | (~new_n17094_ & (~new_n17098_ | new_n17097_));
  assign new_n17119_ = new_n17095_ & new_n17096_;
  assign new_n17120_ = ~new_n17121_ ^ new_n17122_;
  assign new_n17121_ = ~new_n17100_ & new_n17099_;
  assign new_n17122_ = (new_n17102_ & new_n17103_) | (new_n17101_ & (new_n17102_ | new_n17103_));
  assign new_n17123_ = (~new_n17081_ & new_n17080_) | (new_n17079_ & (~new_n17081_ | new_n17080_));
  assign \o[11]  = ~new_n17125_ ^ new_n17126_;
  assign new_n17125_ = (new_n17108_ | (~new_n17109_ & (new_n17107_ | new_n17106_))) & (new_n17107_ | new_n17106_ | ~new_n17109_);
  assign new_n17126_ = new_n17127_ ^ new_n17128_;
  assign new_n17127_ = (~new_n17111_ & new_n17123_) | (new_n17110_ & (~new_n17111_ | new_n17123_));
  assign new_n17128_ = new_n17129_ ? (~new_n17130_ ^ new_n17133_) : (new_n17130_ ^ new_n17133_);
  assign new_n17129_ = (~new_n17117_ & new_n17116_) | (~new_n17112_ & (~new_n17117_ | new_n17116_));
  assign new_n17130_ = ~new_n17131_ ^ new_n17132_;
  assign new_n17131_ = (~new_n17120_ & new_n17119_) | (new_n17118_ & (~new_n17120_ | new_n17119_));
  assign new_n17132_ = new_n17121_ & new_n17122_;
  assign new_n17133_ = (new_n17114_ & new_n17115_) | (new_n17113_ & (new_n17114_ | new_n17115_));
  assign \o[12]  = ((new_n17135_ | new_n17136_) & (~new_n17137_ ^ new_n17138_)) | (~new_n17135_ & ~new_n17136_ & (new_n17137_ ^ new_n17138_));
  assign new_n17135_ = ~new_n17126_ & new_n17125_;
  assign new_n17136_ = ~new_n17128_ & new_n17127_;
  assign new_n17137_ = (~new_n17130_ & new_n17133_) | (new_n17129_ & (~new_n17130_ | new_n17133_));
  assign new_n17138_ = new_n17131_ & new_n17132_;
  assign \o[13]  = (new_n17138_ | new_n17135_ | new_n17136_) & (new_n17137_ | (new_n17138_ & (new_n17135_ | new_n17136_)));
  assign \o[14]  = new_n17141_ ? (new_n19816_ ^ new_n19879_) : (~new_n19816_ ^ new_n19879_);
  assign new_n17141_ = new_n17142_ ? (new_n19031_ ^ new_n19730_) : (~new_n19031_ ^ new_n19730_);
  assign new_n17142_ = new_n17143_ ? (new_n18112_ ^ new_n18957_) : (~new_n18112_ ^ new_n18957_);
  assign new_n17143_ = new_n17144_ ? (~new_n18009_ ^ new_n18106_) : (new_n18009_ ^ new_n18106_);
  assign new_n17144_ = new_n17145_ ? (new_n17671_ ^ new_n17809_) : (~new_n17671_ ^ new_n17809_);
  assign new_n17145_ = new_n17146_ ? (new_n17290_ ^ new_n17451_) : (~new_n17290_ ^ new_n17451_);
  assign new_n17146_ = ~new_n17147_ & new_n17286_;
  assign new_n17147_ = new_n17148_ & (~new_n17259_ | (~new_n17260_ & ~new_n17261_));
  assign new_n17148_ = new_n17149_ & (~new_n17257_ | (~new_n17258_ & new_n14384_) | (new_n17255_ & ~new_n14384_));
  assign new_n17149_ = (~new_n17249_ | new_n17150_) & (~new_n17213_ | (new_n9634_ ? ~new_n17248_ : new_n17250_));
  assign new_n17150_ = (~new_n17151_ & ~new_n17152_) | (~new_n17186_ & new_n17206_ & new_n17210_ & new_n17212_ & new_n17152_);
  assign new_n17151_ = new_n10368_ & new_n8093_;
  assign new_n17152_ = new_n17153_ & new_n17177_;
  assign new_n17153_ = ~new_n17154_ & ~new_n17176_;
  assign new_n17154_ = new_n17155_ & (~new_n17164_ | (new_n17174_ & new_n17175_ & new_n17171_ & new_n17173_));
  assign new_n17155_ = new_n17156_ & ~new_n17160_ & ~new_n17161_;
  assign new_n17156_ = ~new_n17157_ & (\all_features[4763]  | \all_features[4764]  | \all_features[4765]  | \all_features[4766]  | \all_features[4767] );
  assign new_n17157_ = ~\all_features[4765]  & new_n17159_ & ((~\all_features[4762]  & new_n17158_) | ~\all_features[4764]  | ~\all_features[4763] );
  assign new_n17158_ = ~\all_features[4760]  & ~\all_features[4761] ;
  assign new_n17159_ = ~\all_features[4766]  & ~\all_features[4767] ;
  assign new_n17160_ = new_n17159_ & (~\all_features[4765]  | (~\all_features[4764]  & (~\all_features[4763]  | (~\all_features[4762]  & ~\all_features[4761] ))));
  assign new_n17161_ = new_n17159_ & (~\all_features[4763]  | ~new_n17162_ | (~\all_features[4762]  & ~new_n17163_));
  assign new_n17162_ = \all_features[4764]  & \all_features[4765] ;
  assign new_n17163_ = \all_features[4760]  & \all_features[4761] ;
  assign new_n17164_ = ~new_n17170_ & ~new_n17169_ & ~new_n17165_ & ~new_n17167_;
  assign new_n17165_ = ~\all_features[4767]  & (~\all_features[4766]  | (~\all_features[4765]  & (new_n17158_ | ~new_n17166_ | ~\all_features[4764] )));
  assign new_n17166_ = \all_features[4762]  & \all_features[4763] ;
  assign new_n17167_ = ~new_n17168_ & ~\all_features[4767] ;
  assign new_n17168_ = \all_features[4765]  & \all_features[4766]  & (\all_features[4764]  | (\all_features[4762]  & \all_features[4763]  & \all_features[4761] ));
  assign new_n17169_ = ~\all_features[4767]  & (~\all_features[4766]  | ~new_n17162_ | ~new_n17163_ | ~new_n17166_);
  assign new_n17170_ = ~\all_features[4767]  & (~\all_features[4766]  | (~\all_features[4764]  & ~\all_features[4765]  & ~new_n17166_));
  assign new_n17171_ = \all_features[4767]  & (\all_features[4766]  | (\all_features[4765]  & (\all_features[4764]  | ~new_n17158_ | ~new_n17172_)));
  assign new_n17172_ = ~\all_features[4762]  & ~\all_features[4763] ;
  assign new_n17173_ = \all_features[4767]  & (\all_features[4766]  | (new_n17162_ & (\all_features[4762]  | \all_features[4763]  | \all_features[4761] )));
  assign new_n17174_ = \all_features[4766]  & \all_features[4767]  & (\all_features[4764]  | \all_features[4765]  | new_n17163_ | ~new_n17172_);
  assign new_n17175_ = \all_features[4767]  & (\all_features[4765]  | \all_features[4766]  | \all_features[4764] );
  assign new_n17176_ = new_n17155_ & new_n17164_;
  assign new_n17177_ = ~new_n17178_ & ~new_n17182_;
  assign new_n17178_ = new_n17156_ & (new_n17161_ | new_n17160_ | (~new_n17165_ & ~new_n17170_ & ~new_n17179_));
  assign new_n17179_ = ~new_n17169_ & ~new_n17167_ & (~new_n17175_ | ~new_n17171_ | new_n17180_);
  assign new_n17180_ = new_n17173_ & new_n17174_ & (new_n17181_ | ~\all_features[4765]  | ~\all_features[4766]  | ~\all_features[4767] );
  assign new_n17181_ = ~\all_features[4763]  & ~\all_features[4764]  & (~\all_features[4762]  | new_n17158_);
  assign new_n17182_ = ~new_n17183_ & (\all_features[4763]  | \all_features[4764]  | \all_features[4765]  | \all_features[4766]  | \all_features[4767] );
  assign new_n17183_ = ~new_n17157_ & (new_n17160_ | (~new_n17161_ & (new_n17170_ | (~new_n17165_ & ~new_n17184_))));
  assign new_n17184_ = ~new_n17167_ & (new_n17169_ | (new_n17175_ & (~new_n17171_ | (~new_n17185_ & new_n17173_))));
  assign new_n17185_ = ~\all_features[4765]  & \all_features[4766]  & \all_features[4767]  & (\all_features[4764]  ? new_n17172_ : (new_n17163_ | ~new_n17172_));
  assign new_n17186_ = new_n17187_ & (new_n17205_ | new_n17204_ | (~new_n17200_ & ~new_n17202_ & ~new_n17193_));
  assign new_n17187_ = ~new_n17188_ & ~new_n17192_;
  assign new_n17188_ = new_n17189_ & (~\all_features[3843]  | ~new_n17191_ | (~\all_features[3842]  & ~new_n17190_));
  assign new_n17189_ = ~\all_features[3846]  & ~\all_features[3847] ;
  assign new_n17190_ = \all_features[3840]  & \all_features[3841] ;
  assign new_n17191_ = \all_features[3844]  & \all_features[3845] ;
  assign new_n17192_ = new_n17189_ & (~\all_features[3845]  | (~\all_features[3844]  & (~\all_features[3843]  | (~\all_features[3842]  & ~\all_features[3841] ))));
  assign new_n17193_ = \all_features[3847]  & (new_n17197_ | ~new_n17195_ | ~new_n17194_) & (new_n17199_ | \all_features[3846] );
  assign new_n17194_ = \all_features[3847]  & (\all_features[3846]  | (new_n17191_ & (\all_features[3842]  | \all_features[3843]  | \all_features[3841] )));
  assign new_n17195_ = new_n17196_ & (new_n17190_ | \all_features[3842]  | \all_features[3843]  | \all_features[3844]  | \all_features[3845] );
  assign new_n17196_ = \all_features[3846]  & \all_features[3847] ;
  assign new_n17197_ = new_n17196_ & \all_features[3845]  & ((~new_n17198_ & \all_features[3842] ) | \all_features[3844]  | \all_features[3843] );
  assign new_n17198_ = ~\all_features[3840]  & ~\all_features[3841] ;
  assign new_n17199_ = \all_features[3845]  & (\all_features[3842]  | \all_features[3843]  | \all_features[3844]  | ~new_n17198_);
  assign new_n17200_ = ~\all_features[3847]  & (~\all_features[3846]  | ~new_n17190_ | ~new_n17191_ | ~new_n17201_);
  assign new_n17201_ = \all_features[3842]  & \all_features[3843] ;
  assign new_n17202_ = ~new_n17203_ & ~\all_features[3847] ;
  assign new_n17203_ = \all_features[3845]  & \all_features[3846]  & (\all_features[3844]  | (\all_features[3842]  & \all_features[3843]  & \all_features[3841] ));
  assign new_n17204_ = ~\all_features[3847]  & (~\all_features[3846]  | (~\all_features[3844]  & ~\all_features[3845]  & ~new_n17201_));
  assign new_n17205_ = ~\all_features[3847]  & (~\all_features[3846]  | (~\all_features[3845]  & (new_n17198_ | ~new_n17201_ | ~\all_features[3844] )));
  assign new_n17206_ = new_n17208_ & ~new_n17209_ & ~new_n17207_ & ~new_n17192_;
  assign new_n17207_ = ~new_n17200_ & ~new_n17202_ & ~new_n17204_ & ~new_n17205_ & (~new_n17195_ | ~new_n17194_);
  assign new_n17208_ = ~new_n17188_ & (\all_features[3843]  | \all_features[3844]  | \all_features[3845]  | \all_features[3846]  | \all_features[3847] );
  assign new_n17209_ = ~\all_features[3845]  & new_n17189_ & ((~\all_features[3842]  & new_n17198_) | ~\all_features[3844]  | ~\all_features[3843] );
  assign new_n17210_ = new_n17211_ & new_n17187_ & ~new_n17209_ & ~new_n17205_ & ~new_n17202_ & ~new_n17204_;
  assign new_n17211_ = ~new_n17200_ & (\all_features[3843]  | \all_features[3844]  | \all_features[3845]  | \all_features[3846]  | \all_features[3847] );
  assign new_n17212_ = ~new_n17209_ & (\all_features[3843]  | \all_features[3844]  | \all_features[3845]  | \all_features[3846]  | \all_features[3847] );
  assign new_n17213_ = ~new_n17214_ & ~new_n17217_;
  assign new_n17214_ = new_n17215_ & new_n17216_;
  assign new_n17215_ = new_n15986_ & new_n15990_;
  assign new_n17216_ = new_n15958_ & new_n15982_;
  assign new_n17217_ = ~new_n17247_ & (~new_n17244_ | ~new_n17218_);
  assign new_n17218_ = new_n17230_ & (~new_n17233_ | (new_n17236_ & (~new_n17240_ | new_n17219_)));
  assign new_n17219_ = new_n17220_ & (~new_n17225_ | (~new_n17229_ & \all_features[2317]  & \all_features[2318]  & \all_features[2319] ));
  assign new_n17220_ = \all_features[2319]  & (\all_features[2318]  | (~new_n17224_ & new_n17221_));
  assign new_n17221_ = \all_features[2317]  & (\all_features[2316]  | ~new_n17223_ | ~new_n17222_);
  assign new_n17222_ = ~\all_features[2312]  & ~\all_features[2313] ;
  assign new_n17223_ = ~\all_features[2314]  & ~\all_features[2315] ;
  assign new_n17224_ = ~\all_features[2316]  & ~\all_features[2317] ;
  assign new_n17225_ = new_n17226_ & \all_features[2318]  & \all_features[2319]  & (~new_n17223_ | ~new_n17224_ | new_n17228_);
  assign new_n17226_ = \all_features[2319]  & (\all_features[2318]  | (new_n17227_ & (\all_features[2314]  | \all_features[2315]  | \all_features[2313] )));
  assign new_n17227_ = \all_features[2316]  & \all_features[2317] ;
  assign new_n17228_ = \all_features[2312]  & \all_features[2313] ;
  assign new_n17229_ = ~\all_features[2315]  & ~\all_features[2316]  & (~\all_features[2314]  | new_n17222_);
  assign new_n17230_ = ~new_n17231_ & (\all_features[2315]  | \all_features[2316]  | \all_features[2317]  | \all_features[2318]  | \all_features[2319] );
  assign new_n17231_ = ~\all_features[2317]  & new_n17232_ & ((~\all_features[2314]  & new_n17222_) | ~\all_features[2316]  | ~\all_features[2315] );
  assign new_n17232_ = ~\all_features[2318]  & ~\all_features[2319] ;
  assign new_n17233_ = ~new_n17234_ & ~new_n17235_;
  assign new_n17234_ = new_n17232_ & (~\all_features[2315]  | ~new_n17227_ | (~\all_features[2314]  & ~new_n17228_));
  assign new_n17235_ = new_n17232_ & (~\all_features[2317]  | (~\all_features[2316]  & (~\all_features[2315]  | (~\all_features[2314]  & ~\all_features[2313] ))));
  assign new_n17236_ = ~new_n17237_ & ~new_n17239_;
  assign new_n17237_ = ~\all_features[2319]  & (~\all_features[2318]  | (~new_n17238_ & new_n17224_));
  assign new_n17238_ = \all_features[2314]  & \all_features[2315] ;
  assign new_n17239_ = ~\all_features[2319]  & (~\all_features[2318]  | (~\all_features[2317]  & (new_n17222_ | ~new_n17238_ | ~\all_features[2316] )));
  assign new_n17240_ = ~new_n17241_ & ~new_n17242_;
  assign new_n17241_ = ~\all_features[2319]  & (~\all_features[2318]  | ~new_n17228_ | ~new_n17227_ | ~new_n17238_);
  assign new_n17242_ = ~new_n17243_ & ~\all_features[2319] ;
  assign new_n17243_ = \all_features[2317]  & \all_features[2318]  & (\all_features[2316]  | (\all_features[2314]  & \all_features[2315]  & \all_features[2313] ));
  assign new_n17244_ = new_n17245_ & (new_n17239_ | new_n17242_ | ~new_n17246_ | (new_n17225_ & new_n17220_));
  assign new_n17245_ = new_n17230_ & new_n17233_;
  assign new_n17246_ = ~new_n17237_ & ~new_n17241_;
  assign new_n17247_ = new_n17240_ & new_n17245_ & new_n17236_;
  assign new_n17248_ = new_n10936_ & ~new_n10938_ & new_n10912_;
  assign new_n17249_ = new_n14923_ & new_n17217_;
  assign new_n17250_ = ~new_n12680_ & ~new_n12656_ & ~new_n17251_;
  assign new_n17251_ = new_n12674_ & (~new_n12681_ | (~new_n17252_ & ~new_n12670_ & ~new_n12672_));
  assign new_n17252_ = ~new_n12673_ & ~new_n12668_ & (~new_n12666_ | new_n17253_ | ~new_n12658_);
  assign new_n17253_ = ~new_n12665_ & new_n12662_ & \all_features[3782]  & \all_features[3783]  & (~\all_features[3781]  | new_n17254_);
  assign new_n17254_ = ~\all_features[3779]  & ~\all_features[3780]  & (~\all_features[3778]  | new_n12660_);
  assign new_n17255_ = ~new_n12834_ & (~new_n12825_ | ~new_n17256_);
  assign new_n17256_ = new_n12803_ & new_n12829_;
  assign new_n17257_ = ~new_n14923_ & new_n17217_;
  assign new_n17258_ = ~new_n11940_ & ~new_n11935_ & ~new_n11908_ & ~new_n11931_;
  assign new_n17259_ = ~new_n17217_ & new_n17214_;
  assign new_n17260_ = ~new_n12404_ & new_n12375_;
  assign new_n17261_ = new_n17262_ & new_n17284_;
  assign new_n17262_ = new_n17278_ & ~new_n17283_ & ~new_n17263_ & ~new_n17282_;
  assign new_n17263_ = ~new_n17272_ & ~new_n17274_ & ~new_n17276_ & ~new_n17277_ & (~new_n17267_ | ~new_n17264_);
  assign new_n17264_ = \all_features[3767]  & (\all_features[3766]  | (~new_n17265_ & \all_features[3765] ));
  assign new_n17265_ = new_n17266_ & ~\all_features[3764]  & ~\all_features[3762]  & ~\all_features[3763] ;
  assign new_n17266_ = ~\all_features[3760]  & ~\all_features[3761] ;
  assign new_n17267_ = \all_features[3767]  & \all_features[3766]  & ~new_n17270_ & new_n17268_;
  assign new_n17268_ = \all_features[3767]  & (\all_features[3766]  | (new_n17269_ & (\all_features[3762]  | \all_features[3763]  | \all_features[3761] )));
  assign new_n17269_ = \all_features[3764]  & \all_features[3765] ;
  assign new_n17270_ = ~\all_features[3765]  & ~\all_features[3764]  & ~\all_features[3763]  & ~new_n17271_ & ~\all_features[3762] ;
  assign new_n17271_ = \all_features[3760]  & \all_features[3761] ;
  assign new_n17272_ = ~\all_features[3767]  & (~\all_features[3766]  | (~\all_features[3765]  & (new_n17266_ | ~new_n17273_ | ~\all_features[3764] )));
  assign new_n17273_ = \all_features[3762]  & \all_features[3763] ;
  assign new_n17274_ = ~new_n17275_ & ~\all_features[3767] ;
  assign new_n17275_ = \all_features[3765]  & \all_features[3766]  & (\all_features[3764]  | (\all_features[3762]  & \all_features[3763]  & \all_features[3761] ));
  assign new_n17276_ = ~\all_features[3767]  & (~\all_features[3766]  | ~new_n17269_ | ~new_n17271_ | ~new_n17273_);
  assign new_n17277_ = ~\all_features[3767]  & (~\all_features[3766]  | (~\all_features[3764]  & ~\all_features[3765]  & ~new_n17273_));
  assign new_n17278_ = ~new_n17279_ & ~new_n17281_;
  assign new_n17279_ = ~\all_features[3765]  & new_n17280_ & ((~\all_features[3762]  & new_n17266_) | ~\all_features[3764]  | ~\all_features[3763] );
  assign new_n17280_ = ~\all_features[3766]  & ~\all_features[3767] ;
  assign new_n17281_ = ~\all_features[3767]  & ~\all_features[3766]  & ~\all_features[3765]  & ~\all_features[3763]  & ~\all_features[3764] ;
  assign new_n17282_ = new_n17280_ & (~\all_features[3765]  | (~\all_features[3764]  & (~\all_features[3763]  | (~\all_features[3762]  & ~\all_features[3761] ))));
  assign new_n17283_ = new_n17280_ & (~\all_features[3763]  | ~new_n17269_ | (~\all_features[3762]  & ~new_n17271_));
  assign new_n17284_ = new_n17285_ & new_n17278_ & ~new_n17274_ & ~new_n17282_;
  assign new_n17285_ = ~new_n17283_ & ~new_n17277_ & ~new_n17272_ & ~new_n17276_;
  assign new_n17286_ = ~new_n17289_ & new_n17287_ & (new_n17261_ | new_n17260_ | ~new_n17259_);
  assign new_n17287_ = ~new_n17288_ & (~new_n17213_ | (new_n17248_ & new_n9634_) | (~new_n17250_ & ~new_n9634_));
  assign new_n17288_ = new_n17249_ & ~new_n17151_ & ~new_n17152_;
  assign new_n17289_ = new_n17257_ & (new_n14384_ ? ~new_n17258_ : new_n17255_);
  assign new_n17290_ = new_n17324_ & (new_n17391_ | ((new_n17415_ | ~new_n14918_ | ~new_n14084_) & (new_n17291_ | new_n14084_)));
  assign new_n17291_ = (~new_n17320_ & (~new_n17322_ | (~new_n17292_ & ~new_n17313_))) ? new_n12562_ : new_n13674_;
  assign new_n17292_ = ~new_n17293_ & (\all_features[5283]  | \all_features[5284]  | \all_features[5285]  | \all_features[5286]  | \all_features[5287] );
  assign new_n17293_ = ~new_n17309_ & (new_n17307_ | (~new_n17311_ & (new_n17312_ | (~new_n17310_ & ~new_n17294_))));
  assign new_n17294_ = ~new_n17295_ & (new_n17297_ | (new_n17306_ & (~new_n17301_ | (~new_n17305_ & new_n17304_))));
  assign new_n17295_ = ~new_n17296_ & ~\all_features[5287] ;
  assign new_n17296_ = \all_features[5285]  & \all_features[5286]  & (\all_features[5284]  | (\all_features[5282]  & \all_features[5283]  & \all_features[5281] ));
  assign new_n17297_ = ~\all_features[5287]  & (~\all_features[5286]  | ~new_n17298_ | ~new_n17299_ | ~new_n17300_);
  assign new_n17298_ = \all_features[5282]  & \all_features[5283] ;
  assign new_n17299_ = \all_features[5280]  & \all_features[5281] ;
  assign new_n17300_ = \all_features[5284]  & \all_features[5285] ;
  assign new_n17301_ = \all_features[5287]  & (\all_features[5286]  | (\all_features[5285]  & (\all_features[5284]  | ~new_n17303_ | ~new_n17302_)));
  assign new_n17302_ = ~\all_features[5280]  & ~\all_features[5281] ;
  assign new_n17303_ = ~\all_features[5282]  & ~\all_features[5283] ;
  assign new_n17304_ = \all_features[5287]  & (\all_features[5286]  | (new_n17300_ & (\all_features[5282]  | \all_features[5283]  | \all_features[5281] )));
  assign new_n17305_ = ~\all_features[5285]  & \all_features[5286]  & \all_features[5287]  & (\all_features[5284]  ? new_n17303_ : (new_n17299_ | ~new_n17303_));
  assign new_n17306_ = \all_features[5287]  & (\all_features[5285]  | \all_features[5286]  | \all_features[5284] );
  assign new_n17307_ = new_n17308_ & (~\all_features[5285]  | (~\all_features[5284]  & (~\all_features[5283]  | (~\all_features[5282]  & ~\all_features[5281] ))));
  assign new_n17308_ = ~\all_features[5286]  & ~\all_features[5287] ;
  assign new_n17309_ = ~\all_features[5285]  & new_n17308_ & ((~\all_features[5282]  & new_n17302_) | ~\all_features[5284]  | ~\all_features[5283] );
  assign new_n17310_ = ~\all_features[5287]  & (~\all_features[5286]  | (~\all_features[5285]  & (new_n17302_ | ~new_n17298_ | ~\all_features[5284] )));
  assign new_n17311_ = new_n17308_ & (~\all_features[5283]  | ~new_n17300_ | (~\all_features[5282]  & ~new_n17299_));
  assign new_n17312_ = ~\all_features[5287]  & (~\all_features[5286]  | (~\all_features[5284]  & ~\all_features[5285]  & ~new_n17298_));
  assign new_n17313_ = new_n17318_ & (~new_n17319_ | (~new_n17314_ & ~new_n17310_ & ~new_n17312_));
  assign new_n17314_ = ~new_n17295_ & ~new_n17297_ & (~new_n17306_ | ~new_n17301_ | new_n17315_);
  assign new_n17315_ = new_n17304_ & new_n17316_ & (new_n17317_ | ~\all_features[5285]  | ~\all_features[5286]  | ~\all_features[5287] );
  assign new_n17316_ = \all_features[5286]  & \all_features[5287]  & (\all_features[5284]  | \all_features[5285]  | new_n17299_ | ~new_n17303_);
  assign new_n17317_ = ~\all_features[5283]  & ~\all_features[5284]  & (~\all_features[5282]  | new_n17302_);
  assign new_n17318_ = ~new_n17309_ & (\all_features[5283]  | \all_features[5284]  | \all_features[5285]  | \all_features[5286]  | \all_features[5287] );
  assign new_n17319_ = ~new_n17307_ & ~new_n17311_;
  assign new_n17320_ = new_n17321_ & new_n17318_ & ~new_n17311_ & ~new_n17310_ & ~new_n17295_ & ~new_n17307_;
  assign new_n17321_ = ~new_n17297_ & ~new_n17312_;
  assign new_n17322_ = new_n17318_ & new_n17319_ & (new_n17323_ | new_n17295_ | new_n17310_ | ~new_n17321_);
  assign new_n17323_ = new_n17306_ & new_n17316_ & new_n17301_ & new_n17304_;
  assign new_n17324_ = ~new_n17390_ & (~new_n17391_ | (new_n17325_ & ~new_n17448_) | (~new_n17449_ & ~new_n17358_ & new_n17448_));
  assign new_n17325_ = new_n17329_ ? new_n17328_ : new_n17326_;
  assign new_n17326_ = new_n11120_ & new_n17327_ & new_n11097_;
  assign new_n17327_ = new_n15486_ & new_n11123_;
  assign new_n17328_ = ~new_n6833_ & new_n9869_;
  assign new_n17329_ = new_n17357_ & (new_n17353_ | new_n17330_);
  assign new_n17330_ = new_n17350_ & ~new_n17331_ & new_n17345_;
  assign new_n17331_ = ~new_n17339_ & ~new_n17341_ & ~new_n17342_ & ~new_n17344_ & (~new_n17335_ | ~new_n17332_);
  assign new_n17332_ = \all_features[5047]  & (\all_features[5046]  | (~new_n17333_ & \all_features[5045] ));
  assign new_n17333_ = new_n17334_ & ~\all_features[5044]  & ~\all_features[5042]  & ~\all_features[5043] ;
  assign new_n17334_ = ~\all_features[5040]  & ~\all_features[5041] ;
  assign new_n17335_ = \all_features[5047]  & \all_features[5046]  & ~new_n17338_ & new_n17336_;
  assign new_n17336_ = \all_features[5047]  & (\all_features[5046]  | (new_n17337_ & (\all_features[5042]  | \all_features[5043]  | \all_features[5041] )));
  assign new_n17337_ = \all_features[5044]  & \all_features[5045] ;
  assign new_n17338_ = ~\all_features[5042]  & ~\all_features[5043]  & ~\all_features[5044]  & ~\all_features[5045]  & (~\all_features[5041]  | ~\all_features[5040] );
  assign new_n17339_ = ~\all_features[5047]  & (~\all_features[5046]  | (~\all_features[5044]  & ~\all_features[5045]  & ~new_n17340_));
  assign new_n17340_ = \all_features[5042]  & \all_features[5043] ;
  assign new_n17341_ = ~\all_features[5047]  & (~\all_features[5046]  | (~\all_features[5045]  & (new_n17334_ | ~\all_features[5044]  | ~new_n17340_)));
  assign new_n17342_ = ~new_n17343_ & ~\all_features[5047] ;
  assign new_n17343_ = \all_features[5045]  & \all_features[5046]  & (\all_features[5044]  | (\all_features[5042]  & \all_features[5043]  & \all_features[5041] ));
  assign new_n17344_ = ~\all_features[5047]  & (~new_n17337_ | ~\all_features[5040]  | ~\all_features[5041]  | ~\all_features[5046]  | ~new_n17340_);
  assign new_n17345_ = ~new_n17346_ & ~new_n17349_;
  assign new_n17346_ = new_n17347_ & ((~\all_features[5042]  & new_n17334_) | ~\all_features[5044]  | ~\all_features[5043] );
  assign new_n17347_ = ~\all_features[5045]  & new_n17348_;
  assign new_n17348_ = ~\all_features[5046]  & ~\all_features[5047] ;
  assign new_n17349_ = new_n17347_ & ~\all_features[5043]  & ~\all_features[5044] ;
  assign new_n17350_ = ~new_n17351_ & ~new_n17352_;
  assign new_n17351_ = new_n17348_ & (~new_n17337_ | ~\all_features[5043]  | (~\all_features[5042]  & (~\all_features[5040]  | ~\all_features[5041] )));
  assign new_n17352_ = new_n17348_ & (~\all_features[5045]  | (~\all_features[5044]  & (~\all_features[5043]  | (~\all_features[5042]  & ~\all_features[5041] ))));
  assign new_n17353_ = new_n17345_ & (~new_n17350_ | (new_n17356_ & (new_n17354_ | new_n17342_ | new_n17344_)));
  assign new_n17354_ = new_n17332_ & (~new_n17335_ | (~new_n17355_ & \all_features[5045]  & \all_features[5046]  & \all_features[5047] ));
  assign new_n17355_ = ~\all_features[5043]  & ~\all_features[5044]  & (~\all_features[5042]  | new_n17334_);
  assign new_n17356_ = ~new_n17339_ & ~new_n17341_;
  assign new_n17357_ = new_n17350_ & new_n17356_ & ~new_n17344_ & ~new_n17342_ & ~new_n17346_ & ~new_n17349_;
  assign new_n17358_ = ~new_n15167_ & new_n17359_;
  assign new_n17359_ = ~new_n17388_ & ~new_n17382_ & (~new_n17385_ | new_n17360_);
  assign new_n17360_ = new_n17374_ & (new_n17381_ | new_n17372_ | (~new_n17378_ & ~new_n17380_ & ~new_n17361_));
  assign new_n17361_ = new_n17370_ & new_n17371_ & (~new_n17367_ | ~new_n17365_ | new_n17362_);
  assign new_n17362_ = \all_features[3863]  & \all_features[3862]  & ~new_n17363_ & \all_features[3861] ;
  assign new_n17363_ = ~\all_features[3859]  & ~\all_features[3860]  & (~\all_features[3858]  | new_n17364_);
  assign new_n17364_ = ~\all_features[3856]  & ~\all_features[3857] ;
  assign new_n17365_ = \all_features[3863]  & (\all_features[3862]  | (new_n17366_ & (\all_features[3858]  | \all_features[3859]  | \all_features[3857] )));
  assign new_n17366_ = \all_features[3860]  & \all_features[3861] ;
  assign new_n17367_ = \all_features[3862]  & \all_features[3863]  & (\all_features[3860]  | \all_features[3861]  | new_n17369_ | ~new_n17368_);
  assign new_n17368_ = ~\all_features[3858]  & ~\all_features[3859] ;
  assign new_n17369_ = \all_features[3856]  & \all_features[3857] ;
  assign new_n17370_ = \all_features[3863]  & (\all_features[3862]  | (\all_features[3861]  & (\all_features[3860]  | ~new_n17368_ | ~new_n17364_)));
  assign new_n17371_ = \all_features[3863]  & (\all_features[3861]  | \all_features[3862]  | \all_features[3860] );
  assign new_n17372_ = ~\all_features[3863]  & (~\all_features[3862]  | new_n17373_);
  assign new_n17373_ = ~\all_features[3861]  & (new_n17364_ | ~\all_features[3859]  | ~\all_features[3860]  | ~\all_features[3858] );
  assign new_n17374_ = ~new_n17375_ & ~new_n17377_;
  assign new_n17375_ = new_n17376_ & (~\all_features[3861]  | (~\all_features[3860]  & (~\all_features[3859]  | (~\all_features[3858]  & ~\all_features[3857] ))));
  assign new_n17376_ = ~\all_features[3862]  & ~\all_features[3863] ;
  assign new_n17377_ = new_n17376_ & (~\all_features[3859]  | ~new_n17366_ | (~new_n17369_ & ~\all_features[3858] ));
  assign new_n17378_ = ~new_n17379_ & ~\all_features[3863] ;
  assign new_n17379_ = \all_features[3861]  & \all_features[3862]  & (\all_features[3860]  | (\all_features[3858]  & \all_features[3859]  & \all_features[3857] ));
  assign new_n17380_ = ~\all_features[3863]  & (~new_n17369_ | ~\all_features[3858]  | ~\all_features[3859]  | ~\all_features[3862]  | ~new_n17366_);
  assign new_n17381_ = ~\all_features[3863]  & (~\all_features[3862]  | (~\all_features[3861]  & ~\all_features[3860]  & (~\all_features[3859]  | ~\all_features[3858] )));
  assign new_n17382_ = new_n17374_ & ~new_n17383_ & new_n17385_;
  assign new_n17383_ = ~new_n17381_ & ~new_n17380_ & ~new_n17378_ & ~new_n17372_ & ~new_n17384_;
  assign new_n17384_ = new_n17371_ & new_n17370_ & new_n17365_ & new_n17367_;
  assign new_n17385_ = ~new_n17386_ & ~new_n17387_;
  assign new_n17386_ = ~\all_features[3861]  & new_n17376_ & ((~\all_features[3858]  & new_n17364_) | ~\all_features[3860]  | ~\all_features[3859] );
  assign new_n17387_ = ~\all_features[3863]  & ~\all_features[3862]  & ~\all_features[3861]  & ~\all_features[3859]  & ~\all_features[3860] ;
  assign new_n17388_ = new_n17385_ & new_n17389_ & ~new_n17378_ & ~new_n17375_;
  assign new_n17389_ = ~new_n17381_ & ~new_n17377_ & ~new_n17372_ & ~new_n17380_;
  assign new_n17390_ = new_n17415_ & new_n14084_ & ~new_n7097_ & ~new_n17391_;
  assign new_n17391_ = ~new_n17392_ & ~new_n17414_;
  assign new_n17392_ = new_n17393_ & (~new_n17407_ | (new_n17402_ & new_n17404_));
  assign new_n17393_ = new_n17394_ & ~new_n17399_ & ~new_n17400_;
  assign new_n17394_ = ~new_n17395_ & ~new_n17398_;
  assign new_n17395_ = ~\all_features[3885]  & new_n17397_ & ((~\all_features[3882]  & new_n17396_) | ~\all_features[3884]  | ~\all_features[3883] );
  assign new_n17396_ = ~\all_features[3880]  & ~\all_features[3881] ;
  assign new_n17397_ = ~\all_features[3886]  & ~\all_features[3887] ;
  assign new_n17398_ = ~\all_features[3887]  & ~\all_features[3886]  & ~\all_features[3885]  & ~\all_features[3883]  & ~\all_features[3884] ;
  assign new_n17399_ = new_n17397_ & (~\all_features[3885]  | (~\all_features[3884]  & (~\all_features[3883]  | (~\all_features[3882]  & ~\all_features[3881] ))));
  assign new_n17400_ = new_n17397_ & (~new_n17401_ | ~\all_features[3883]  | (~\all_features[3882]  & (~\all_features[3880]  | ~\all_features[3881] )));
  assign new_n17401_ = \all_features[3884]  & \all_features[3885] ;
  assign new_n17402_ = \all_features[3887]  & (\all_features[3886]  | (~new_n17403_ & \all_features[3885] ));
  assign new_n17403_ = new_n17396_ & ~\all_features[3884]  & ~\all_features[3882]  & ~\all_features[3883] ;
  assign new_n17404_ = \all_features[3887]  & \all_features[3886]  & ~new_n17406_ & new_n17405_;
  assign new_n17405_ = \all_features[3887]  & (\all_features[3886]  | (new_n17401_ & (\all_features[3882]  | \all_features[3883]  | \all_features[3881] )));
  assign new_n17406_ = ~\all_features[3882]  & ~\all_features[3883]  & ~\all_features[3884]  & ~\all_features[3885]  & (~\all_features[3881]  | ~\all_features[3880] );
  assign new_n17407_ = ~new_n17413_ & ~new_n17412_ & ~new_n17408_ & ~new_n17410_;
  assign new_n17408_ = ~\all_features[3887]  & (~\all_features[3886]  | (~\all_features[3885]  & (new_n17396_ | ~new_n17409_ | ~\all_features[3884] )));
  assign new_n17409_ = \all_features[3882]  & \all_features[3883] ;
  assign new_n17410_ = ~new_n17411_ & ~\all_features[3887] ;
  assign new_n17411_ = \all_features[3885]  & \all_features[3886]  & (\all_features[3884]  | (\all_features[3882]  & \all_features[3883]  & \all_features[3881] ));
  assign new_n17412_ = ~\all_features[3887]  & (~\all_features[3886]  | (~\all_features[3884]  & ~\all_features[3885]  & ~new_n17409_));
  assign new_n17413_ = ~\all_features[3887]  & (~new_n17409_ | ~\all_features[3880]  | ~\all_features[3881]  | ~\all_features[3886]  | ~new_n17401_);
  assign new_n17414_ = new_n17393_ & new_n17407_;
  assign new_n17415_ = ~new_n17446_ & ~new_n17444_ & ~new_n17416_ & ~new_n17437_;
  assign new_n17416_ = ~new_n17417_ & (\all_features[4411]  | \all_features[4412]  | \all_features[4413]  | \all_features[4414]  | \all_features[4415] );
  assign new_n17417_ = ~new_n17431_ & (new_n17433_ | (~new_n17434_ & (new_n17435_ | (~new_n17418_ & ~new_n17436_))));
  assign new_n17418_ = ~new_n17419_ & (new_n17421_ | (new_n17430_ & (~new_n17425_ | (~new_n17429_ & new_n17428_))));
  assign new_n17419_ = ~new_n17420_ & ~\all_features[4415] ;
  assign new_n17420_ = \all_features[4413]  & \all_features[4414]  & (\all_features[4412]  | (\all_features[4410]  & \all_features[4411]  & \all_features[4409] ));
  assign new_n17421_ = ~\all_features[4415]  & (~\all_features[4414]  | ~new_n17422_ | ~new_n17423_ | ~new_n17424_);
  assign new_n17422_ = \all_features[4408]  & \all_features[4409] ;
  assign new_n17423_ = \all_features[4412]  & \all_features[4413] ;
  assign new_n17424_ = \all_features[4410]  & \all_features[4411] ;
  assign new_n17425_ = \all_features[4415]  & (\all_features[4414]  | (\all_features[4413]  & (\all_features[4412]  | ~new_n17427_ | ~new_n17426_)));
  assign new_n17426_ = ~\all_features[4408]  & ~\all_features[4409] ;
  assign new_n17427_ = ~\all_features[4410]  & ~\all_features[4411] ;
  assign new_n17428_ = \all_features[4415]  & (\all_features[4414]  | (new_n17423_ & (\all_features[4410]  | \all_features[4411]  | \all_features[4409] )));
  assign new_n17429_ = ~\all_features[4413]  & \all_features[4414]  & \all_features[4415]  & (\all_features[4412]  ? new_n17427_ : (new_n17422_ | ~new_n17427_));
  assign new_n17430_ = \all_features[4415]  & (\all_features[4413]  | \all_features[4414]  | \all_features[4412] );
  assign new_n17431_ = ~\all_features[4413]  & new_n17432_ & ((~\all_features[4410]  & new_n17426_) | ~\all_features[4412]  | ~\all_features[4411] );
  assign new_n17432_ = ~\all_features[4414]  & ~\all_features[4415] ;
  assign new_n17433_ = new_n17432_ & (~\all_features[4413]  | (~\all_features[4412]  & (~\all_features[4411]  | (~\all_features[4410]  & ~\all_features[4409] ))));
  assign new_n17434_ = new_n17432_ & (~\all_features[4411]  | ~new_n17423_ | (~\all_features[4410]  & ~new_n17422_));
  assign new_n17435_ = ~\all_features[4415]  & (~\all_features[4414]  | (~\all_features[4412]  & ~\all_features[4413]  & ~new_n17424_));
  assign new_n17436_ = ~\all_features[4415]  & (~\all_features[4414]  | (~\all_features[4413]  & (new_n17426_ | ~new_n17424_ | ~\all_features[4412] )));
  assign new_n17437_ = new_n17442_ & (~new_n17443_ | (~new_n17438_ & ~new_n17435_ & ~new_n17436_));
  assign new_n17438_ = ~new_n17419_ & ~new_n17421_ & (~new_n17430_ | ~new_n17425_ | new_n17439_);
  assign new_n17439_ = new_n17428_ & new_n17440_ & (new_n17441_ | ~\all_features[4413]  | ~\all_features[4414]  | ~\all_features[4415] );
  assign new_n17440_ = \all_features[4414]  & \all_features[4415]  & (\all_features[4412]  | \all_features[4413]  | new_n17422_ | ~new_n17427_);
  assign new_n17441_ = ~\all_features[4411]  & ~\all_features[4412]  & (~\all_features[4410]  | new_n17426_);
  assign new_n17442_ = ~new_n17431_ & (\all_features[4411]  | \all_features[4412]  | \all_features[4413]  | \all_features[4414]  | \all_features[4415] );
  assign new_n17443_ = ~new_n17433_ & ~new_n17434_;
  assign new_n17444_ = new_n17445_ & new_n17442_ & ~new_n17419_ & ~new_n17436_ & ~new_n17433_ & ~new_n17434_;
  assign new_n17445_ = ~new_n17435_ & ~new_n17421_;
  assign new_n17446_ = new_n17442_ & new_n17443_ & (new_n17447_ | new_n17436_ | new_n17419_ | ~new_n17445_);
  assign new_n17447_ = new_n17430_ & new_n17440_ & new_n17425_ & new_n17428_;
  assign new_n17448_ = new_n12001_ & ~new_n14085_ & new_n11978_;
  assign new_n17449_ = ~new_n9649_ & ~new_n17359_ & (~new_n9650_ | new_n17450_);
  assign new_n17450_ = ~new_n8031_ & ~new_n9645_;
  assign new_n17451_ = ~new_n17452_ & new_n17632_;
  assign new_n17452_ = new_n17453_ & (new_n17454_ | (~new_n17587_ & ~new_n17630_) | (~new_n17623_ & new_n17630_));
  assign new_n17453_ = ~new_n17454_ | ((new_n16611_ | ~new_n17489_ | ~new_n17471_) & (new_n17471_ | (~new_n17554_ & ~new_n17520_)));
  assign new_n17454_ = new_n17455_ & (new_n8333_ | (~new_n17468_ & ~new_n8341_));
  assign new_n17455_ = ~new_n8327_ & ((~new_n17456_ & new_n8334_ & new_n17465_) | new_n8333_ | new_n8341_);
  assign new_n17456_ = ~new_n8340_ & ~new_n8343_ & (new_n8329_ | new_n8338_ | new_n17457_);
  assign new_n17457_ = new_n17464_ & ~new_n17460_ & new_n17458_;
  assign new_n17458_ = \all_features[3335]  & (\all_features[3334]  | new_n17459_);
  assign new_n17459_ = \all_features[3333]  & (\all_features[3330]  | \all_features[3331]  | \all_features[3332]  | ~new_n8342_);
  assign new_n17460_ = ~new_n17462_ & new_n17461_ & \all_features[3334]  & \all_features[3335]  & (~\all_features[3333]  | new_n17463_);
  assign new_n17461_ = \all_features[3335]  & (\all_features[3334]  | (new_n8331_ & (\all_features[3330]  | \all_features[3331]  | \all_features[3329] )));
  assign new_n17462_ = ~\all_features[3333]  & ~\all_features[3332]  & ~\all_features[3331]  & ~new_n8330_ & ~\all_features[3330] ;
  assign new_n17463_ = ~\all_features[3331]  & ~\all_features[3332]  & (~\all_features[3330]  | new_n8342_);
  assign new_n17464_ = \all_features[3335]  & (\all_features[3333]  | \all_features[3334]  | \all_features[3332] );
  assign new_n17465_ = new_n17467_ & (~new_n17461_ | ~new_n17464_ | ~new_n17466_ | ~new_n17458_);
  assign new_n17466_ = \all_features[3335]  & ~new_n17462_ & \all_features[3334] ;
  assign new_n17467_ = ~new_n8343_ & ~new_n8340_ & ~new_n8338_ & ~new_n8329_;
  assign new_n17468_ = ~new_n8337_ & (new_n8335_ | (~new_n8340_ & (new_n8343_ | (~new_n17469_ & ~new_n8338_))));
  assign new_n17469_ = ~new_n8329_ & (~new_n17464_ | (new_n17458_ & (~new_n17461_ | (~new_n17470_ & new_n17466_))));
  assign new_n17470_ = \all_features[3334]  & \all_features[3335]  & (\all_features[3333]  | (\all_features[3332]  & (\all_features[3331]  | \all_features[3330] )));
  assign new_n17471_ = new_n17480_ & ~new_n17472_ & ~new_n17485_;
  assign new_n17472_ = ~new_n17473_ & (\all_features[4859]  | \all_features[4860]  | \all_features[4861]  | \all_features[4862]  | \all_features[4863] );
  assign new_n17473_ = ~new_n14851_ & (new_n14862_ | (~new_n14864_ & (new_n14859_ | (~new_n14863_ & ~new_n17474_))));
  assign new_n17474_ = ~new_n14860_ & (new_n14855_ | (new_n17479_ & (~new_n17475_ | (~new_n17478_ & new_n17477_))));
  assign new_n17475_ = \all_features[4863]  & (\all_features[4862]  | (\all_features[4861]  & (\all_features[4860]  | ~new_n17476_ | ~new_n14853_)));
  assign new_n17476_ = ~\all_features[4858]  & ~\all_features[4859] ;
  assign new_n17477_ = \all_features[4863]  & (\all_features[4862]  | (new_n14858_ & (\all_features[4858]  | \all_features[4859]  | \all_features[4857] )));
  assign new_n17478_ = ~\all_features[4861]  & \all_features[4862]  & \all_features[4863]  & (\all_features[4860]  ? new_n17476_ : (new_n14857_ | ~new_n17476_));
  assign new_n17479_ = \all_features[4863]  & (\all_features[4861]  | \all_features[4862]  | \all_features[4860] );
  assign new_n17480_ = ~new_n14849_ & (new_n17481_ | ~new_n14850_ | ~new_n17484_);
  assign new_n17481_ = ~new_n14860_ & ~new_n14863_ & new_n14854_ & (~new_n17475_ | ~new_n17482_);
  assign new_n17482_ = new_n17479_ & new_n17477_ & new_n17483_;
  assign new_n17483_ = \all_features[4862]  & \all_features[4863]  & (\all_features[4860]  | \all_features[4861]  | new_n14857_ | ~new_n17476_);
  assign new_n17484_ = ~new_n14862_ & ~new_n14864_;
  assign new_n17485_ = new_n14850_ & (~new_n17484_ | (~new_n17486_ & ~new_n14863_ & ~new_n14859_));
  assign new_n17486_ = ~new_n14860_ & ~new_n14855_ & (~new_n17479_ | ~new_n17475_ | new_n17487_);
  assign new_n17487_ = new_n17477_ & new_n17483_ & (new_n17488_ | ~\all_features[4861]  | ~\all_features[4862]  | ~\all_features[4863] );
  assign new_n17488_ = ~\all_features[4859]  & ~\all_features[4860]  & (~\all_features[4858]  | new_n14853_);
  assign new_n17489_ = ~new_n17518_ & (new_n17519_ | new_n17490_);
  assign new_n17490_ = new_n17509_ & (new_n17514_ | (~new_n17515_ & new_n17491_ & (new_n17501_ | new_n17507_)));
  assign new_n17491_ = ~new_n17501_ & ~new_n17503_ & (~new_n17506_ | ~new_n17505_ | new_n17492_);
  assign new_n17492_ = new_n17493_ & ~new_n17499_ & new_n17495_;
  assign new_n17493_ = \all_features[5535]  & (\all_features[5534]  | (new_n17494_ & (\all_features[5530]  | \all_features[5531]  | \all_features[5529] )));
  assign new_n17494_ = \all_features[5532]  & \all_features[5533] ;
  assign new_n17495_ = new_n17498_ & (new_n17496_ | \all_features[5532]  | \all_features[5533]  | ~new_n17497_);
  assign new_n17496_ = \all_features[5528]  & \all_features[5529] ;
  assign new_n17497_ = ~\all_features[5530]  & ~\all_features[5531] ;
  assign new_n17498_ = \all_features[5534]  & \all_features[5535] ;
  assign new_n17499_ = new_n17498_ & \all_features[5533]  & ((~new_n17500_ & \all_features[5530] ) | \all_features[5532]  | \all_features[5531] );
  assign new_n17500_ = ~\all_features[5528]  & ~\all_features[5529] ;
  assign new_n17501_ = ~new_n17502_ & ~\all_features[5535] ;
  assign new_n17502_ = \all_features[5533]  & \all_features[5534]  & (\all_features[5532]  | (\all_features[5530]  & \all_features[5531]  & \all_features[5529] ));
  assign new_n17503_ = ~\all_features[5535]  & (~\all_features[5534]  | ~new_n17504_ | ~new_n17496_ | ~new_n17494_);
  assign new_n17504_ = \all_features[5530]  & \all_features[5531] ;
  assign new_n17505_ = \all_features[5535]  & (\all_features[5534]  | (\all_features[5533]  & (\all_features[5532]  | ~new_n17497_ | ~new_n17500_)));
  assign new_n17506_ = \all_features[5535]  & (\all_features[5533]  | \all_features[5534]  | \all_features[5532] );
  assign new_n17507_ = ~new_n17503_ & (~new_n17506_ | (new_n17505_ & (~new_n17493_ | (~new_n17508_ & new_n17495_))));
  assign new_n17508_ = new_n17498_ & (\all_features[5533]  | (~new_n17497_ & \all_features[5532] ));
  assign new_n17509_ = ~new_n17513_ & ~new_n17510_ & ~new_n17512_;
  assign new_n17510_ = new_n17511_ & (~\all_features[5533]  | (~\all_features[5532]  & (~\all_features[5531]  | (~\all_features[5530]  & ~\all_features[5529] ))));
  assign new_n17511_ = ~\all_features[5534]  & ~\all_features[5535] ;
  assign new_n17512_ = new_n17511_ & (~\all_features[5531]  | ~new_n17494_ | (~\all_features[5530]  & ~new_n17496_));
  assign new_n17513_ = ~\all_features[5533]  & new_n17511_ & ((~\all_features[5530]  & new_n17500_) | ~\all_features[5532]  | ~\all_features[5531] );
  assign new_n17514_ = ~\all_features[5535]  & (~\all_features[5534]  | (~\all_features[5532]  & ~\all_features[5533]  & ~new_n17504_));
  assign new_n17515_ = ~\all_features[5535]  & (~\all_features[5534]  | (~\all_features[5533]  & (new_n17500_ | ~\all_features[5532]  | ~new_n17504_)));
  assign new_n17517_ = ~new_n17503_ & ~new_n17501_ & ~new_n17514_ & ~new_n17515_;
  assign new_n17518_ = ~new_n17519_ & ~new_n17513_ & ~new_n17510_ & ~new_n17512_;
  assign new_n17519_ = ~\all_features[5535]  & ~\all_features[5534]  & ~\all_features[5533]  & ~\all_features[5531]  & ~\all_features[5532] ;
  assign new_n17520_ = new_n17553_ & (new_n17521_ | (new_n17544_ & new_n17549_));
  assign new_n17521_ = ~new_n17543_ & ~new_n17542_ & ~new_n17541_ & ~new_n17522_ & ~new_n17539_;
  assign new_n17522_ = ~new_n17523_ & ~new_n17537_ & new_n17526_ & (~new_n17538_ | ~new_n17530_);
  assign new_n17523_ = ~\all_features[4399]  & (~\all_features[4398]  | new_n17524_);
  assign new_n17524_ = ~\all_features[4397]  & (new_n17525_ | ~\all_features[4395]  | ~\all_features[4396]  | ~\all_features[4394] );
  assign new_n17525_ = ~\all_features[4392]  & ~\all_features[4393] ;
  assign new_n17526_ = ~new_n17527_ & ~new_n17529_;
  assign new_n17527_ = ~new_n17528_ & ~\all_features[4399] ;
  assign new_n17528_ = \all_features[4397]  & \all_features[4398]  & (\all_features[4396]  | (\all_features[4394]  & \all_features[4395]  & \all_features[4393] ));
  assign new_n17529_ = ~\all_features[4399]  & (~\all_features[4398]  | (~\all_features[4397]  & ~\all_features[4396]  & (~\all_features[4395]  | ~\all_features[4394] )));
  assign new_n17530_ = new_n17536_ & new_n17531_ & new_n17533_;
  assign new_n17531_ = \all_features[4399]  & (\all_features[4398]  | (new_n17532_ & (\all_features[4394]  | \all_features[4395]  | \all_features[4393] )));
  assign new_n17532_ = \all_features[4396]  & \all_features[4397] ;
  assign new_n17533_ = \all_features[4398]  & \all_features[4399]  & (\all_features[4396]  | \all_features[4397]  | new_n17534_ | ~new_n17535_);
  assign new_n17534_ = \all_features[4392]  & \all_features[4393] ;
  assign new_n17535_ = ~\all_features[4394]  & ~\all_features[4395] ;
  assign new_n17536_ = \all_features[4399]  & (\all_features[4397]  | \all_features[4398]  | \all_features[4396] );
  assign new_n17537_ = ~\all_features[4399]  & (~new_n17532_ | ~\all_features[4394]  | ~\all_features[4395]  | ~\all_features[4398]  | ~new_n17534_);
  assign new_n17538_ = \all_features[4399]  & (\all_features[4398]  | (\all_features[4397]  & (\all_features[4396]  | ~new_n17535_ | ~new_n17525_)));
  assign new_n17539_ = new_n17540_ & (~\all_features[4395]  | ~new_n17532_ | (~\all_features[4394]  & ~new_n17534_));
  assign new_n17540_ = ~\all_features[4398]  & ~\all_features[4399] ;
  assign new_n17541_ = new_n17540_ & (~\all_features[4397]  | (~\all_features[4396]  & (~\all_features[4395]  | (~\all_features[4394]  & ~\all_features[4393] ))));
  assign new_n17542_ = ~\all_features[4397]  & new_n17540_ & ((~\all_features[4394]  & new_n17525_) | ~\all_features[4396]  | ~\all_features[4395] );
  assign new_n17543_ = ~\all_features[4399]  & ~\all_features[4398]  & ~\all_features[4397]  & ~\all_features[4395]  & ~\all_features[4396] ;
  assign new_n17544_ = ~new_n17543_ & ~new_n17542_ & (~new_n17548_ | (~new_n17545_ & ~new_n17523_ & ~new_n17529_));
  assign new_n17545_ = ~new_n17537_ & ~new_n17527_ & (~new_n17536_ | ~new_n17538_ | new_n17546_);
  assign new_n17546_ = new_n17531_ & new_n17533_ & (new_n17547_ | ~\all_features[4397]  | ~\all_features[4398]  | ~\all_features[4399] );
  assign new_n17547_ = ~\all_features[4395]  & ~\all_features[4396]  & (~\all_features[4394]  | new_n17525_);
  assign new_n17548_ = ~new_n17539_ & ~new_n17541_;
  assign new_n17549_ = ~new_n17550_ & ~new_n17543_;
  assign new_n17550_ = ~new_n17542_ & (new_n17541_ | (~new_n17539_ & (new_n17529_ | (~new_n17523_ & ~new_n17551_))));
  assign new_n17551_ = ~new_n17527_ & (new_n17537_ | (new_n17536_ & (~new_n17538_ | (~new_n17552_ & new_n17531_))));
  assign new_n17552_ = ~\all_features[4397]  & \all_features[4398]  & \all_features[4399]  & (\all_features[4396]  ? new_n17535_ : (new_n17534_ | ~new_n17535_));
  assign new_n17553_ = new_n17548_ & new_n17526_ & ~new_n17543_ & ~new_n17537_ & ~new_n17523_ & ~new_n17542_;
  assign new_n17554_ = ~new_n17555_ & new_n17582_;
  assign new_n17555_ = ~new_n17581_ & (~new_n17574_ | (~new_n17579_ & (new_n17572_ | new_n17580_ | ~new_n17556_)));
  assign new_n17556_ = ~new_n17568_ & ~new_n17566_ & ((~new_n17563_ & new_n17557_) | ~new_n17571_ | ~new_n17570_);
  assign new_n17557_ = \all_features[3751]  & \all_features[3750]  & ~new_n17560_ & new_n17558_;
  assign new_n17558_ = \all_features[3751]  & (\all_features[3750]  | (new_n17559_ & (\all_features[3746]  | \all_features[3747]  | \all_features[3745] )));
  assign new_n17559_ = \all_features[3748]  & \all_features[3749] ;
  assign new_n17560_ = new_n17562_ & ~\all_features[3749]  & ~new_n17561_ & ~\all_features[3748] ;
  assign new_n17561_ = \all_features[3744]  & \all_features[3745] ;
  assign new_n17562_ = ~\all_features[3746]  & ~\all_features[3747] ;
  assign new_n17563_ = \all_features[3751]  & \all_features[3750]  & ~new_n17564_ & \all_features[3749] ;
  assign new_n17564_ = ~\all_features[3747]  & ~\all_features[3748]  & (~\all_features[3746]  | new_n17565_);
  assign new_n17565_ = ~\all_features[3744]  & ~\all_features[3745] ;
  assign new_n17566_ = ~new_n17567_ & ~\all_features[3751] ;
  assign new_n17567_ = \all_features[3749]  & \all_features[3750]  & (\all_features[3748]  | (\all_features[3746]  & \all_features[3747]  & \all_features[3745] ));
  assign new_n17568_ = ~\all_features[3751]  & (~\all_features[3750]  | ~new_n17569_ | ~new_n17561_ | ~new_n17559_);
  assign new_n17569_ = \all_features[3746]  & \all_features[3747] ;
  assign new_n17570_ = \all_features[3751]  & (\all_features[3750]  | (\all_features[3749]  & (\all_features[3748]  | ~new_n17562_ | ~new_n17565_)));
  assign new_n17571_ = \all_features[3751]  & (\all_features[3749]  | \all_features[3750]  | \all_features[3748] );
  assign new_n17572_ = ~new_n17566_ & (new_n17568_ | (new_n17571_ & (~new_n17570_ | (~new_n17573_ & new_n17558_))));
  assign new_n17573_ = ~\all_features[3749]  & \all_features[3750]  & \all_features[3751]  & (\all_features[3748]  ? new_n17562_ : (new_n17561_ | ~new_n17562_));
  assign new_n17574_ = ~new_n17578_ & ~new_n17575_ & ~new_n17577_;
  assign new_n17575_ = new_n17576_ & (~\all_features[3749]  | (~\all_features[3748]  & (~\all_features[3747]  | (~\all_features[3746]  & ~\all_features[3745] ))));
  assign new_n17576_ = ~\all_features[3750]  & ~\all_features[3751] ;
  assign new_n17577_ = ~\all_features[3749]  & new_n17576_ & ((~\all_features[3746]  & new_n17565_) | ~\all_features[3748]  | ~\all_features[3747] );
  assign new_n17578_ = new_n17576_ & (~\all_features[3747]  | ~new_n17559_ | (~\all_features[3746]  & ~new_n17561_));
  assign new_n17579_ = ~\all_features[3751]  & (~\all_features[3750]  | (~\all_features[3748]  & ~\all_features[3749]  & ~new_n17569_));
  assign new_n17580_ = ~\all_features[3751]  & (~\all_features[3750]  | (~\all_features[3749]  & (new_n17565_ | ~\all_features[3748]  | ~new_n17569_)));
  assign new_n17581_ = ~\all_features[3751]  & ~\all_features[3750]  & ~\all_features[3749]  & ~\all_features[3747]  & ~\all_features[3748] ;
  assign new_n17582_ = new_n17575_ | ~new_n17585_ | ((new_n17566_ | ~new_n17586_) & (new_n17583_ | new_n17578_));
  assign new_n17583_ = new_n17584_ & (~new_n17557_ | ~new_n17570_ | ~new_n17571_);
  assign new_n17584_ = ~new_n17568_ & ~new_n17566_ & ~new_n17579_ & ~new_n17580_;
  assign new_n17585_ = ~new_n17577_ & ~new_n17581_;
  assign new_n17586_ = ~new_n17578_ & ~new_n17568_ & ~new_n17579_ & ~new_n17580_;
  assign new_n17587_ = new_n12730_ & new_n17588_;
  assign new_n17588_ = new_n17621_ & (new_n17619_ | ~new_n17589_);
  assign new_n17589_ = ~new_n17590_ & ~new_n17612_;
  assign new_n17590_ = ~new_n17611_ & (new_n17609_ | (~new_n17607_ & (new_n17610_ | (~new_n17591_ & ~new_n17606_))));
  assign new_n17591_ = ~new_n17600_ & (new_n17603_ | (~new_n17602_ & (~new_n17605_ | (~new_n17592_ & new_n17598_))));
  assign new_n17592_ = new_n17593_ & (\all_features[3741]  | ~new_n17596_ | (~new_n17597_ & ~\all_features[3740]  & new_n17595_) | (\all_features[3740]  & ~new_n17595_));
  assign new_n17593_ = \all_features[3743]  & (\all_features[3742]  | (new_n17594_ & (\all_features[3738]  | \all_features[3739]  | \all_features[3737] )));
  assign new_n17594_ = \all_features[3740]  & \all_features[3741] ;
  assign new_n17595_ = ~\all_features[3738]  & ~\all_features[3739] ;
  assign new_n17596_ = \all_features[3742]  & \all_features[3743] ;
  assign new_n17597_ = \all_features[3736]  & \all_features[3737] ;
  assign new_n17598_ = \all_features[3743]  & (\all_features[3742]  | (\all_features[3741]  & (\all_features[3740]  | ~new_n17599_ | ~new_n17595_)));
  assign new_n17599_ = ~\all_features[3736]  & ~\all_features[3737] ;
  assign new_n17600_ = ~\all_features[3743]  & (~\all_features[3742]  | (~\all_features[3741]  & (new_n17599_ | ~new_n17601_ | ~\all_features[3740] )));
  assign new_n17601_ = \all_features[3738]  & \all_features[3739] ;
  assign new_n17602_ = ~\all_features[3743]  & (~\all_features[3742]  | ~new_n17594_ | ~new_n17597_ | ~new_n17601_);
  assign new_n17603_ = ~new_n17604_ & ~\all_features[3743] ;
  assign new_n17604_ = \all_features[3741]  & \all_features[3742]  & (\all_features[3740]  | (\all_features[3738]  & \all_features[3739]  & \all_features[3737] ));
  assign new_n17605_ = \all_features[3743]  & (\all_features[3741]  | \all_features[3742]  | \all_features[3740] );
  assign new_n17606_ = ~\all_features[3743]  & (~\all_features[3742]  | (~\all_features[3740]  & ~\all_features[3741]  & ~new_n17601_));
  assign new_n17607_ = new_n17608_ & (~\all_features[3741]  | (~\all_features[3740]  & (~\all_features[3739]  | (~\all_features[3738]  & ~\all_features[3737] ))));
  assign new_n17608_ = ~\all_features[3742]  & ~\all_features[3743] ;
  assign new_n17609_ = ~\all_features[3741]  & new_n17608_ & ((~\all_features[3738]  & new_n17599_) | ~\all_features[3740]  | ~\all_features[3739] );
  assign new_n17610_ = new_n17608_ & (~\all_features[3739]  | ~new_n17594_ | (~\all_features[3738]  & ~new_n17597_));
  assign new_n17611_ = ~\all_features[3743]  & ~\all_features[3742]  & ~\all_features[3741]  & ~\all_features[3739]  & ~\all_features[3740] ;
  assign new_n17612_ = ~new_n17609_ & ~new_n17611_ & (~new_n17618_ | (~new_n17613_ & new_n17617_));
  assign new_n17613_ = new_n17614_ & ((~new_n17616_ & new_n17615_ & new_n17593_) | ~new_n17605_ | ~new_n17598_);
  assign new_n17614_ = ~new_n17602_ & ~new_n17603_;
  assign new_n17615_ = new_n17596_ & (new_n17597_ | \all_features[3740]  | \all_features[3741]  | ~new_n17595_);
  assign new_n17616_ = new_n17596_ & \all_features[3741]  & ((~new_n17599_ & \all_features[3738] ) | \all_features[3740]  | \all_features[3739] );
  assign new_n17617_ = ~new_n17606_ & ~new_n17600_;
  assign new_n17618_ = ~new_n17607_ & ~new_n17610_;
  assign new_n17619_ = ~new_n17611_ & ~new_n17610_ & ~new_n17609_ & ~new_n17620_ & ~new_n17607_;
  assign new_n17620_ = new_n17617_ & new_n17614_ & (~new_n17615_ | ~new_n17605_ | ~new_n17598_ | ~new_n17593_);
  assign new_n17621_ = new_n17618_ & new_n17622_ & ~new_n17609_ & ~new_n17603_ & ~new_n17606_ & ~new_n17600_;
  assign new_n17622_ = ~new_n17602_ & ~new_n17611_;
  assign new_n17623_ = (~new_n16234_ & new_n16263_) ? (new_n12049_ & new_n12081_) : new_n17624_;
  assign new_n17624_ = new_n17625_ & (~new_n17626_ | ~new_n12220_);
  assign new_n17625_ = ~new_n12198_ & ~new_n12226_;
  assign new_n17626_ = ~new_n17627_ & (\all_features[5259]  | \all_features[5260]  | \all_features[5261]  | \all_features[5262]  | \all_features[5263] );
  assign new_n17627_ = ~new_n12219_ & (new_n12218_ | (~new_n12216_ & (new_n12203_ | (~new_n12213_ & ~new_n17628_))));
  assign new_n17628_ = ~new_n12201_ & (new_n12205_ | (new_n12214_ & (~new_n12208_ | (~new_n17629_ & new_n12211_))));
  assign new_n17629_ = ~\all_features[5261]  & \all_features[5262]  & \all_features[5263]  & (\all_features[5260]  ? new_n12209_ : (new_n12207_ | ~new_n12209_));
  assign new_n17630_ = ~new_n12851_ & new_n17631_;
  assign new_n17631_ = ~new_n11551_ & ~new_n11573_;
  assign new_n17632_ = ~new_n17633_ & new_n17634_ & (new_n17454_ | (new_n17587_ & ~new_n17630_) | (new_n17623_ & new_n17630_));
  assign new_n17633_ = new_n17454_ & ~new_n17554_ & ~new_n17471_ & ~new_n17520_;
  assign new_n17634_ = ~new_n17471_ | ~new_n17454_ | (new_n17489_ ? ~new_n16611_ : new_n17635_);
  assign new_n17635_ = new_n17636_ & new_n17662_;
  assign new_n17636_ = ~new_n17637_ & ~new_n17659_;
  assign new_n17637_ = new_n17654_ & ~new_n17658_ & ~new_n17638_ & ~new_n17657_;
  assign new_n17638_ = new_n17639_ & ~new_n17652_ & (~new_n17647_ | ~new_n17653_ | ~new_n17650_ | ~new_n17651_);
  assign new_n17639_ = ~new_n17644_ & ~new_n17640_ & ~new_n17642_;
  assign new_n17640_ = ~new_n17641_ & ~\all_features[4655] ;
  assign new_n17641_ = \all_features[4653]  & \all_features[4654]  & (\all_features[4652]  | (\all_features[4650]  & \all_features[4651]  & \all_features[4649] ));
  assign new_n17642_ = ~\all_features[4655]  & (~\all_features[4654]  | (~\all_features[4652]  & ~\all_features[4653]  & ~new_n17643_));
  assign new_n17643_ = \all_features[4650]  & \all_features[4651] ;
  assign new_n17644_ = ~\all_features[4655]  & (~\all_features[4654]  | ~new_n17645_ | ~new_n17646_ | ~new_n17643_);
  assign new_n17645_ = \all_features[4652]  & \all_features[4653] ;
  assign new_n17646_ = \all_features[4648]  & \all_features[4649] ;
  assign new_n17647_ = \all_features[4655]  & (\all_features[4654]  | (\all_features[4653]  & (\all_features[4652]  | ~new_n17649_ | ~new_n17648_)));
  assign new_n17648_ = ~\all_features[4650]  & ~\all_features[4651] ;
  assign new_n17649_ = ~\all_features[4648]  & ~\all_features[4649] ;
  assign new_n17650_ = \all_features[4655]  & (\all_features[4654]  | (new_n17645_ & (\all_features[4650]  | \all_features[4651]  | \all_features[4649] )));
  assign new_n17651_ = \all_features[4654]  & \all_features[4655]  & (\all_features[4652]  | \all_features[4653]  | new_n17646_ | ~new_n17648_);
  assign new_n17652_ = ~\all_features[4655]  & (~\all_features[4654]  | (~\all_features[4653]  & (new_n17649_ | ~new_n17643_ | ~\all_features[4652] )));
  assign new_n17653_ = \all_features[4655]  & (\all_features[4653]  | \all_features[4654]  | \all_features[4652] );
  assign new_n17654_ = ~new_n17655_ & (\all_features[4651]  | \all_features[4652]  | \all_features[4653]  | \all_features[4654]  | \all_features[4655] );
  assign new_n17655_ = new_n17656_ & (~\all_features[4651]  | ~new_n17645_ | (~\all_features[4650]  & ~new_n17646_));
  assign new_n17656_ = ~\all_features[4654]  & ~\all_features[4655] ;
  assign new_n17657_ = new_n17656_ & (~\all_features[4653]  | (~\all_features[4652]  & (~\all_features[4651]  | (~\all_features[4650]  & ~\all_features[4649] ))));
  assign new_n17658_ = ~\all_features[4653]  & new_n17656_ & ((~\all_features[4650]  & new_n17649_) | ~\all_features[4652]  | ~\all_features[4651] );
  assign new_n17659_ = new_n17639_ & new_n17661_ & ~new_n17652_ & new_n17660_;
  assign new_n17660_ = ~new_n17658_ & (\all_features[4651]  | \all_features[4652]  | \all_features[4653]  | \all_features[4654]  | \all_features[4655] );
  assign new_n17661_ = ~new_n17657_ & ~new_n17655_;
  assign new_n17662_ = ~new_n17663_ & ~new_n17667_;
  assign new_n17663_ = ~new_n17664_ & (\all_features[4651]  | \all_features[4652]  | \all_features[4653]  | \all_features[4654]  | \all_features[4655] );
  assign new_n17664_ = ~new_n17658_ & (new_n17657_ | (~new_n17655_ & (new_n17642_ | (~new_n17652_ & ~new_n17665_))));
  assign new_n17665_ = ~new_n17640_ & (new_n17644_ | (new_n17653_ & (~new_n17647_ | (~new_n17666_ & new_n17650_))));
  assign new_n17666_ = ~\all_features[4653]  & \all_features[4654]  & \all_features[4655]  & (\all_features[4652]  ? new_n17648_ : (new_n17646_ | ~new_n17648_));
  assign new_n17667_ = new_n17660_ & (~new_n17661_ | (~new_n17668_ & ~new_n17652_ & ~new_n17642_));
  assign new_n17668_ = ~new_n17644_ & ~new_n17640_ & (~new_n17653_ | ~new_n17647_ | new_n17669_);
  assign new_n17669_ = new_n17650_ & new_n17651_ & (new_n17670_ | ~\all_features[4653]  | ~\all_features[4654]  | ~\all_features[4655] );
  assign new_n17670_ = ~\all_features[4651]  & ~\all_features[4652]  & (~\all_features[4650]  | new_n17649_);
  assign new_n17671_ = new_n17672_ & new_n17806_;
  assign new_n17672_ = new_n17673_ & (~new_n17805_ | ~new_n16527_) & (new_n17675_ ? new_n17767_ : new_n17764_);
  assign new_n17673_ = (~new_n17674_ | new_n17736_) & (~new_n17710_ | ~new_n17675_ | ~new_n7475_);
  assign new_n17674_ = ~new_n17709_ & ~new_n13134_ & ~new_n17675_;
  assign new_n17675_ = new_n17676_ & ~new_n17701_ & ~new_n17705_;
  assign new_n17676_ = ~new_n17677_ & ~new_n17699_;
  assign new_n17677_ = new_n17694_ & ~new_n17698_ & ~new_n17678_ & ~new_n17697_;
  assign new_n17678_ = new_n17679_ & (~new_n17692_ | ~new_n17693_ | ~new_n17689_ | ~new_n17691_);
  assign new_n17679_ = ~new_n17686_ & ~new_n17684_ & ~new_n17680_ & ~new_n17682_;
  assign new_n17680_ = ~\all_features[2327]  & (~\all_features[2326]  | (~\all_features[2324]  & ~\all_features[2325]  & ~new_n17681_));
  assign new_n17681_ = \all_features[2322]  & \all_features[2323] ;
  assign new_n17682_ = ~\all_features[2327]  & (~\all_features[2326]  | (~\all_features[2325]  & (new_n17683_ | ~new_n17681_ | ~\all_features[2324] )));
  assign new_n17683_ = ~\all_features[2320]  & ~\all_features[2321] ;
  assign new_n17684_ = ~new_n17685_ & ~\all_features[2327] ;
  assign new_n17685_ = \all_features[2325]  & \all_features[2326]  & (\all_features[2324]  | (\all_features[2322]  & \all_features[2323]  & \all_features[2321] ));
  assign new_n17686_ = ~\all_features[2327]  & (~\all_features[2326]  | ~new_n17687_ | ~new_n17688_ | ~new_n17681_);
  assign new_n17687_ = \all_features[2320]  & \all_features[2321] ;
  assign new_n17688_ = \all_features[2324]  & \all_features[2325] ;
  assign new_n17689_ = \all_features[2327]  & (\all_features[2326]  | (\all_features[2325]  & (\all_features[2324]  | ~new_n17690_ | ~new_n17683_)));
  assign new_n17690_ = ~\all_features[2322]  & ~\all_features[2323] ;
  assign new_n17691_ = \all_features[2327]  & (\all_features[2326]  | (new_n17688_ & (\all_features[2322]  | \all_features[2323]  | \all_features[2321] )));
  assign new_n17692_ = \all_features[2326]  & \all_features[2327]  & (\all_features[2324]  | \all_features[2325]  | new_n17687_ | ~new_n17690_);
  assign new_n17693_ = \all_features[2327]  & (\all_features[2325]  | \all_features[2326]  | \all_features[2324] );
  assign new_n17694_ = ~new_n17695_ & (\all_features[2323]  | \all_features[2324]  | \all_features[2325]  | \all_features[2326]  | \all_features[2327] );
  assign new_n17695_ = ~\all_features[2325]  & new_n17696_ & ((~\all_features[2322]  & new_n17683_) | ~\all_features[2324]  | ~\all_features[2323] );
  assign new_n17696_ = ~\all_features[2326]  & ~\all_features[2327] ;
  assign new_n17697_ = new_n17696_ & (~\all_features[2325]  | (~\all_features[2324]  & (~\all_features[2323]  | (~\all_features[2322]  & ~\all_features[2321] ))));
  assign new_n17698_ = new_n17696_ & (~\all_features[2323]  | ~new_n17688_ | (~\all_features[2322]  & ~new_n17687_));
  assign new_n17699_ = new_n17700_ & new_n17694_ & ~new_n17697_ & ~new_n17684_;
  assign new_n17700_ = ~new_n17686_ & ~new_n17682_ & ~new_n17698_ & ~new_n17680_;
  assign new_n17701_ = ~new_n17702_ & (\all_features[2323]  | \all_features[2324]  | \all_features[2325]  | \all_features[2326]  | \all_features[2327] );
  assign new_n17702_ = ~new_n17695_ & (new_n17697_ | (~new_n17698_ & (new_n17680_ | (~new_n17703_ & ~new_n17682_))));
  assign new_n17703_ = ~new_n17684_ & (new_n17686_ | (new_n17693_ & (~new_n17689_ | (~new_n17704_ & new_n17691_))));
  assign new_n17704_ = ~\all_features[2325]  & \all_features[2326]  & \all_features[2327]  & (\all_features[2324]  ? new_n17690_ : (new_n17687_ | ~new_n17690_));
  assign new_n17705_ = new_n17694_ & (new_n17698_ | new_n17697_ | (~new_n17706_ & ~new_n17680_ & ~new_n17682_));
  assign new_n17706_ = ~new_n17684_ & ~new_n17686_ & (~new_n17693_ | ~new_n17689_ | new_n17707_);
  assign new_n17707_ = new_n17691_ & new_n17692_ & (new_n17708_ | ~\all_features[2325]  | ~\all_features[2326]  | ~\all_features[2327] );
  assign new_n17708_ = ~\all_features[2323]  & ~\all_features[2324]  & (~\all_features[2322]  | new_n17683_);
  assign new_n17709_ = new_n16707_ & (new_n16709_ | new_n16680_);
  assign new_n17710_ = ~new_n17711_ & ~new_n17734_;
  assign new_n17711_ = new_n17729_ & ~new_n17733_ & ~new_n17712_ & ~new_n17732_;
  assign new_n17712_ = ~new_n17727_ & ~new_n17728_ & new_n17720_ & (~new_n17725_ | ~new_n17713_);
  assign new_n17713_ = new_n17719_ & new_n17714_ & new_n17716_;
  assign new_n17714_ = \all_features[5439]  & (\all_features[5438]  | (new_n17715_ & (\all_features[5434]  | \all_features[5435]  | \all_features[5433] )));
  assign new_n17715_ = \all_features[5436]  & \all_features[5437] ;
  assign new_n17716_ = \all_features[5438]  & \all_features[5439]  & (\all_features[5436]  | \all_features[5437]  | new_n17718_ | ~new_n17717_);
  assign new_n17717_ = ~\all_features[5434]  & ~\all_features[5435] ;
  assign new_n17718_ = \all_features[5432]  & \all_features[5433] ;
  assign new_n17719_ = \all_features[5439]  & (\all_features[5437]  | \all_features[5438]  | \all_features[5436] );
  assign new_n17720_ = ~new_n17721_ & ~new_n17723_;
  assign new_n17721_ = ~new_n17722_ & ~\all_features[5439] ;
  assign new_n17722_ = \all_features[5437]  & \all_features[5438]  & (\all_features[5436]  | (\all_features[5434]  & \all_features[5435]  & \all_features[5433] ));
  assign new_n17723_ = ~\all_features[5439]  & (~\all_features[5438]  | (~\all_features[5436]  & ~\all_features[5437]  & ~new_n17724_));
  assign new_n17724_ = \all_features[5434]  & \all_features[5435] ;
  assign new_n17725_ = \all_features[5439]  & (\all_features[5438]  | (\all_features[5437]  & (\all_features[5436]  | ~new_n17726_ | ~new_n17717_)));
  assign new_n17726_ = ~\all_features[5432]  & ~\all_features[5433] ;
  assign new_n17727_ = ~\all_features[5439]  & (~\all_features[5438]  | (~\all_features[5437]  & (new_n17726_ | ~new_n17724_ | ~\all_features[5436] )));
  assign new_n17728_ = ~\all_features[5439]  & (~\all_features[5438]  | ~new_n17715_ | ~new_n17718_ | ~new_n17724_);
  assign new_n17729_ = ~new_n17730_ & (\all_features[5435]  | \all_features[5436]  | \all_features[5437]  | \all_features[5438]  | \all_features[5439] );
  assign new_n17730_ = ~\all_features[5437]  & new_n17731_ & ((~\all_features[5434]  & new_n17726_) | ~\all_features[5436]  | ~\all_features[5435] );
  assign new_n17731_ = ~\all_features[5438]  & ~\all_features[5439] ;
  assign new_n17732_ = new_n17731_ & (~\all_features[5437]  | (~\all_features[5436]  & (~\all_features[5435]  | (~\all_features[5434]  & ~\all_features[5433] ))));
  assign new_n17733_ = new_n17731_ & (~\all_features[5435]  | ~new_n17715_ | (~\all_features[5434]  & ~new_n17718_));
  assign new_n17734_ = new_n17729_ & new_n17720_ & new_n17735_ & ~new_n17727_ & ~new_n17728_;
  assign new_n17735_ = ~new_n17732_ & ~new_n17733_;
  assign new_n17736_ = ~new_n17757_ & (new_n17752_ | new_n17756_ | ~new_n17737_ | (new_n17759_ & ~new_n17760_));
  assign new_n17737_ = ~new_n17756_ & ~new_n17755_ & ~new_n17754_ & ~new_n17738_ & ~new_n17752_;
  assign new_n17738_ = ~new_n17751_ & ~new_n17750_ & ~new_n17748_ & ~new_n17739_ & ~new_n17746_;
  assign new_n17739_ = \all_features[4015]  & \all_features[4014]  & ~new_n17744_ & new_n17742_;
  assign new_n17740_ = \all_features[4013]  & (\all_features[4010]  | \all_features[4011]  | \all_features[4012]  | ~new_n17741_);
  assign new_n17741_ = ~\all_features[4008]  & ~\all_features[4009] ;
  assign new_n17742_ = \all_features[4015]  & (\all_features[4014]  | (new_n17743_ & (\all_features[4010]  | \all_features[4011]  | \all_features[4009] )));
  assign new_n17743_ = \all_features[4012]  & \all_features[4013] ;
  assign new_n17744_ = ~\all_features[4013]  & ~\all_features[4012]  & ~\all_features[4011]  & ~new_n17745_ & ~\all_features[4010] ;
  assign new_n17745_ = \all_features[4008]  & \all_features[4009] ;
  assign new_n17746_ = ~new_n17747_ & ~\all_features[4015] ;
  assign new_n17747_ = \all_features[4013]  & \all_features[4014]  & (\all_features[4012]  | (\all_features[4010]  & \all_features[4011]  & \all_features[4009] ));
  assign new_n17748_ = ~\all_features[4015]  & (~\all_features[4014]  | ~new_n17745_ | ~new_n17743_ | ~new_n17749_);
  assign new_n17749_ = \all_features[4010]  & \all_features[4011] ;
  assign new_n17750_ = ~\all_features[4015]  & (~\all_features[4014]  | (~\all_features[4012]  & ~\all_features[4013]  & ~new_n17749_));
  assign new_n17751_ = ~\all_features[4015]  & (~\all_features[4014]  | (~\all_features[4013]  & (new_n17741_ | ~\all_features[4012]  | ~new_n17749_)));
  assign new_n17752_ = ~\all_features[4013]  & new_n17753_ & ((~\all_features[4010]  & new_n17741_) | ~\all_features[4012]  | ~\all_features[4011] );
  assign new_n17753_ = ~\all_features[4014]  & ~\all_features[4015] ;
  assign new_n17754_ = new_n17753_ & (~\all_features[4011]  | ~new_n17743_ | (~\all_features[4010]  & ~new_n17745_));
  assign new_n17755_ = new_n17753_ & (~\all_features[4013]  | (~\all_features[4012]  & (~\all_features[4011]  | (~\all_features[4010]  & ~\all_features[4009] ))));
  assign new_n17756_ = ~\all_features[4015]  & ~\all_features[4014]  & ~\all_features[4013]  & ~\all_features[4011]  & ~\all_features[4012] ;
  assign new_n17757_ = new_n17759_ & new_n17758_ & ~new_n17751_ & ~new_n17752_ & ~new_n17746_ & ~new_n17750_;
  assign new_n17758_ = ~new_n17748_ & ~new_n17756_;
  assign new_n17759_ = ~new_n17754_ & ~new_n17755_;
  assign new_n17760_ = ~new_n17750_ & ~new_n17751_ & ((~new_n17762_ & new_n17761_) | new_n17748_ | new_n17746_);
  assign new_n17761_ = \all_features[4015]  & (\all_features[4014]  | new_n17740_);
  assign new_n17762_ = ~new_n17744_ & new_n17742_ & \all_features[4014]  & \all_features[4015]  & (~\all_features[4013]  | new_n17763_);
  assign new_n17763_ = ~\all_features[4011]  & ~\all_features[4012]  & (~\all_features[4010]  | new_n17741_);
  assign new_n17764_ = new_n13134_ ? ~new_n17765_ : ~new_n17709_;
  assign new_n17765_ = ~new_n14416_ & (~new_n14394_ | ~new_n17766_);
  assign new_n17766_ = new_n14418_ & new_n14422_;
  assign new_n17767_ = (new_n17768_ | new_n17804_ | new_n17710_) & (new_n7475_ | ~new_n17769_ | ~new_n17710_);
  assign new_n17768_ = ~new_n11444_ & (~new_n11442_ | ~new_n11412_);
  assign new_n17769_ = ~new_n17802_ & (~new_n17800_ | ~new_n17770_);
  assign new_n17770_ = new_n17771_ & new_n17791_;
  assign new_n17771_ = ~new_n17790_ & (new_n17788_ | (~new_n17785_ & (new_n17787_ | (~new_n17772_ & ~new_n17789_))));
  assign new_n17772_ = ~new_n17783_ & (new_n17779_ | (~new_n17781_ & (~new_n17784_ | new_n17773_)));
  assign new_n17773_ = \all_features[2735]  & ((~new_n17778_ & ~\all_features[2733]  & \all_features[2734] ) | (~new_n17776_ & (\all_features[2734]  | (~new_n17774_ & \all_features[2733] ))));
  assign new_n17774_ = new_n17775_ & ~\all_features[2732]  & ~\all_features[2730]  & ~\all_features[2731] ;
  assign new_n17775_ = ~\all_features[2728]  & ~\all_features[2729] ;
  assign new_n17776_ = \all_features[2735]  & (\all_features[2734]  | (new_n17777_ & (\all_features[2730]  | \all_features[2731]  | \all_features[2729] )));
  assign new_n17777_ = \all_features[2732]  & \all_features[2733] ;
  assign new_n17778_ = (~\all_features[2730]  & ~\all_features[2731]  & ~\all_features[2732]  & (~\all_features[2729]  | ~\all_features[2728] )) | (\all_features[2732]  & (\all_features[2730]  | \all_features[2731] ));
  assign new_n17779_ = ~new_n17780_ & ~\all_features[2735] ;
  assign new_n17780_ = \all_features[2733]  & \all_features[2734]  & (\all_features[2732]  | (\all_features[2730]  & \all_features[2731]  & \all_features[2729] ));
  assign new_n17781_ = ~\all_features[2735]  & (~new_n17777_ | ~\all_features[2728]  | ~\all_features[2729]  | ~\all_features[2734]  | ~new_n17782_);
  assign new_n17782_ = \all_features[2730]  & \all_features[2731] ;
  assign new_n17783_ = ~\all_features[2735]  & (~\all_features[2734]  | (~\all_features[2733]  & (new_n17775_ | ~\all_features[2732]  | ~new_n17782_)));
  assign new_n17784_ = \all_features[2735]  & (\all_features[2733]  | \all_features[2734]  | \all_features[2732] );
  assign new_n17785_ = new_n17786_ & (~\all_features[2733]  | (~\all_features[2732]  & (~\all_features[2731]  | (~\all_features[2730]  & ~\all_features[2729] ))));
  assign new_n17786_ = ~\all_features[2734]  & ~\all_features[2735] ;
  assign new_n17787_ = new_n17786_ & (~new_n17777_ | ~\all_features[2731]  | (~\all_features[2730]  & (~\all_features[2728]  | ~\all_features[2729] )));
  assign new_n17788_ = ~\all_features[2733]  & new_n17786_ & ((~\all_features[2730]  & new_n17775_) | ~\all_features[2732]  | ~\all_features[2731] );
  assign new_n17789_ = ~\all_features[2735]  & (~\all_features[2734]  | (~\all_features[2732]  & ~\all_features[2733]  & ~new_n17782_));
  assign new_n17790_ = ~\all_features[2735]  & ~\all_features[2734]  & ~\all_features[2733]  & ~\all_features[2731]  & ~\all_features[2732] ;
  assign new_n17791_ = new_n17798_ & (~new_n17799_ | (~new_n17792_ & ~new_n17783_ & ~new_n17789_));
  assign new_n17792_ = ~new_n17779_ & ~new_n17781_ & (~new_n17793_ | (~new_n17796_ & new_n17794_));
  assign new_n17793_ = \all_features[2735]  & (\all_features[2734]  | (~new_n17774_ & \all_features[2733] ));
  assign new_n17794_ = \all_features[2735]  & \all_features[2734]  & ~new_n17795_ & new_n17776_;
  assign new_n17795_ = ~\all_features[2730]  & ~\all_features[2731]  & ~\all_features[2732]  & ~\all_features[2733]  & (~\all_features[2729]  | ~\all_features[2728] );
  assign new_n17796_ = \all_features[2735]  & \all_features[2734]  & ~new_n17797_ & \all_features[2733] ;
  assign new_n17797_ = ~\all_features[2731]  & ~\all_features[2732]  & (~\all_features[2730]  | new_n17775_);
  assign new_n17798_ = ~new_n17788_ & ~new_n17790_;
  assign new_n17799_ = ~new_n17785_ & ~new_n17787_;
  assign new_n17800_ = new_n17799_ & ~new_n17801_ & new_n17798_;
  assign new_n17801_ = ~new_n17779_ & ~new_n17781_ & ~new_n17783_ & ~new_n17789_ & (~new_n17794_ | ~new_n17793_);
  assign new_n17802_ = new_n17803_ & ~new_n17790_ & ~new_n17781_ & ~new_n17779_ & ~new_n17785_;
  assign new_n17803_ = ~new_n17789_ & ~new_n17788_ & ~new_n17783_ & ~new_n17787_;
  assign new_n17804_ = ~new_n14119_ & ~new_n14122_;
  assign new_n17805_ = new_n13134_ & ~new_n17675_ & ~new_n17765_;
  assign new_n17806_ = ~new_n17807_ & new_n17808_ & (~new_n17674_ | ~new_n17736_) & (~new_n17805_ | new_n16527_);
  assign new_n17807_ = ~new_n17710_ & new_n17804_ & new_n17675_ & (~new_n12791_ | ~new_n12761_);
  assign new_n17808_ = ~new_n17675_ | ((new_n17769_ | new_n7475_ | ~new_n17710_) & (new_n17804_ | ~new_n17768_ | new_n17710_));
  assign new_n17809_ = new_n17810_ ? (~new_n17890_ ^ new_n17971_) : (new_n17890_ ^ new_n17971_);
  assign new_n17810_ = ~new_n17854_ & ~new_n17811_ & (~new_n17816_ | (new_n17842_ & new_n17889_) | (new_n17847_ & ~new_n17889_));
  assign new_n17811_ = ~new_n17814_ & ~new_n17816_ & (new_n9308_ ? new_n17812_ : ~new_n17328_);
  assign new_n17812_ = ~new_n11516_ & new_n17813_;
  assign new_n17813_ = ~new_n11545_ & ~new_n11547_;
  assign new_n17814_ = ~new_n17815_ & new_n8411_;
  assign new_n17815_ = ~new_n8438_ & ~new_n8442_;
  assign new_n17816_ = new_n17817_ & new_n17840_;
  assign new_n17817_ = new_n17835_ & ~new_n17839_ & ~new_n17818_ & ~new_n17838_;
  assign new_n17818_ = ~new_n17833_ & ~new_n17834_ & new_n17826_ & (~new_n17831_ | ~new_n17819_);
  assign new_n17819_ = new_n17825_ & new_n17820_ & new_n17822_;
  assign new_n17820_ = \all_features[4815]  & (\all_features[4814]  | (new_n17821_ & (\all_features[4810]  | \all_features[4811]  | \all_features[4809] )));
  assign new_n17821_ = \all_features[4812]  & \all_features[4813] ;
  assign new_n17822_ = \all_features[4814]  & \all_features[4815]  & (\all_features[4812]  | \all_features[4813]  | new_n17824_ | ~new_n17823_);
  assign new_n17823_ = ~\all_features[4810]  & ~\all_features[4811] ;
  assign new_n17824_ = \all_features[4808]  & \all_features[4809] ;
  assign new_n17825_ = \all_features[4815]  & (\all_features[4813]  | \all_features[4814]  | \all_features[4812] );
  assign new_n17826_ = ~new_n17827_ & ~new_n17829_;
  assign new_n17827_ = ~new_n17828_ & ~\all_features[4815] ;
  assign new_n17828_ = \all_features[4813]  & \all_features[4814]  & (\all_features[4812]  | (\all_features[4810]  & \all_features[4811]  & \all_features[4809] ));
  assign new_n17829_ = ~\all_features[4815]  & (~\all_features[4814]  | (~\all_features[4812]  & ~\all_features[4813]  & ~new_n17830_));
  assign new_n17830_ = \all_features[4810]  & \all_features[4811] ;
  assign new_n17831_ = \all_features[4815]  & (\all_features[4814]  | (\all_features[4813]  & (\all_features[4812]  | ~new_n17832_ | ~new_n17823_)));
  assign new_n17832_ = ~\all_features[4808]  & ~\all_features[4809] ;
  assign new_n17833_ = ~\all_features[4815]  & (~\all_features[4814]  | (~\all_features[4813]  & (new_n17832_ | ~new_n17830_ | ~\all_features[4812] )));
  assign new_n17834_ = ~\all_features[4815]  & (~\all_features[4814]  | ~new_n17821_ | ~new_n17824_ | ~new_n17830_);
  assign new_n17835_ = ~new_n17836_ & (\all_features[4811]  | \all_features[4812]  | \all_features[4813]  | \all_features[4814]  | \all_features[4815] );
  assign new_n17836_ = ~\all_features[4813]  & new_n17837_ & ((~\all_features[4810]  & new_n17832_) | ~\all_features[4812]  | ~\all_features[4811] );
  assign new_n17837_ = ~\all_features[4814]  & ~\all_features[4815] ;
  assign new_n17838_ = new_n17837_ & (~\all_features[4813]  | (~\all_features[4812]  & (~\all_features[4811]  | (~\all_features[4810]  & ~\all_features[4809] ))));
  assign new_n17839_ = new_n17837_ & (~\all_features[4811]  | ~new_n17821_ | (~\all_features[4810]  & ~new_n17824_));
  assign new_n17840_ = new_n17835_ & new_n17826_ & new_n17841_ & ~new_n17833_ & ~new_n17834_;
  assign new_n17841_ = ~new_n17838_ & ~new_n17839_;
  assign new_n17842_ = (~new_n17846_ & ~new_n17843_) | (~new_n13838_ & new_n17843_ & (~new_n13840_ | new_n17845_));
  assign new_n17843_ = new_n13038_ & (new_n13015_ | new_n17844_);
  assign new_n17844_ = new_n14339_ & new_n14343_;
  assign new_n17845_ = ~new_n13809_ & ~new_n13830_;
  assign new_n17846_ = new_n16263_ & new_n16235_ & new_n16261_;
  assign new_n17847_ = new_n16479_ ? new_n17848_ : (new_n8619_ | (~new_n8621_ & new_n8596_));
  assign new_n17848_ = new_n15702_ & (new_n15676_ | ~new_n17849_);
  assign new_n17849_ = ~new_n15703_ & ~new_n17850_;
  assign new_n17850_ = ~new_n15696_ & (new_n15695_ | new_n17851_);
  assign new_n17851_ = ~new_n15691_ & (new_n15693_ | (~new_n15686_ & (new_n15687_ | (~new_n15679_ & ~new_n17852_))));
  assign new_n17852_ = ~new_n15681_ & (~new_n15701_ | (new_n15700_ & (~new_n15697_ | (~new_n17853_ & new_n15698_))));
  assign new_n17853_ = \all_features[2150]  & \all_features[2151]  & (\all_features[2149]  | (~new_n15699_ & \all_features[2148] ));
  assign new_n17854_ = new_n17814_ & ~new_n17855_ & ~new_n17816_;
  assign new_n17855_ = (new_n10024_ & (~new_n10027_ | new_n10002_)) ? ~new_n17856_ : new_n14436_;
  assign new_n17856_ = new_n17888_ & new_n17886_ & new_n17857_ & new_n17877_;
  assign new_n17857_ = ~new_n17876_ & (new_n17871_ | (~new_n17873_ & (new_n17874_ | (~new_n17858_ & ~new_n17875_))));
  assign new_n17858_ = ~new_n17865_ & (new_n17867_ | (~new_n17869_ & (~new_n17870_ | new_n17859_)));
  assign new_n17859_ = \all_features[1983]  & ((~new_n17864_ & ~\all_features[1981]  & \all_features[1982] ) | (~new_n17862_ & (\all_features[1982]  | (~new_n17860_ & \all_features[1981] ))));
  assign new_n17860_ = new_n17861_ & ~\all_features[1980]  & ~\all_features[1978]  & ~\all_features[1979] ;
  assign new_n17861_ = ~\all_features[1976]  & ~\all_features[1977] ;
  assign new_n17862_ = \all_features[1983]  & (\all_features[1982]  | (new_n17863_ & (\all_features[1978]  | \all_features[1979]  | \all_features[1977] )));
  assign new_n17863_ = \all_features[1980]  & \all_features[1981] ;
  assign new_n17864_ = (~\all_features[1978]  & ~\all_features[1979]  & ~\all_features[1980]  & (~\all_features[1977]  | ~\all_features[1976] )) | (\all_features[1980]  & (\all_features[1978]  | \all_features[1979] ));
  assign new_n17865_ = ~\all_features[1983]  & (~\all_features[1982]  | (~\all_features[1981]  & (new_n17861_ | ~new_n17866_ | ~\all_features[1980] )));
  assign new_n17866_ = \all_features[1978]  & \all_features[1979] ;
  assign new_n17867_ = ~new_n17868_ & ~\all_features[1983] ;
  assign new_n17868_ = \all_features[1981]  & \all_features[1982]  & (\all_features[1980]  | (\all_features[1978]  & \all_features[1979]  & \all_features[1977] ));
  assign new_n17869_ = ~\all_features[1983]  & (~new_n17866_ | ~\all_features[1976]  | ~\all_features[1977]  | ~\all_features[1982]  | ~new_n17863_);
  assign new_n17870_ = \all_features[1983]  & (\all_features[1981]  | \all_features[1982]  | \all_features[1980] );
  assign new_n17871_ = ~\all_features[1981]  & new_n17872_ & ((~\all_features[1978]  & new_n17861_) | ~\all_features[1980]  | ~\all_features[1979] );
  assign new_n17872_ = ~\all_features[1982]  & ~\all_features[1983] ;
  assign new_n17873_ = new_n17872_ & (~\all_features[1981]  | (~\all_features[1980]  & (~\all_features[1979]  | (~\all_features[1978]  & ~\all_features[1977] ))));
  assign new_n17874_ = new_n17872_ & (~new_n17863_ | ~\all_features[1979]  | (~\all_features[1978]  & (~\all_features[1976]  | ~\all_features[1977] )));
  assign new_n17875_ = ~\all_features[1983]  & (~\all_features[1982]  | (~\all_features[1980]  & ~\all_features[1981]  & ~new_n17866_));
  assign new_n17876_ = ~\all_features[1983]  & ~\all_features[1982]  & ~\all_features[1981]  & ~\all_features[1979]  & ~\all_features[1980] ;
  assign new_n17877_ = new_n17883_ & (~new_n17884_ | (new_n17885_ & (new_n17878_ | new_n17867_ | new_n17869_)));
  assign new_n17878_ = new_n17879_ & (~new_n17880_ | (~new_n17882_ & \all_features[1981]  & \all_features[1982]  & \all_features[1983] ));
  assign new_n17879_ = \all_features[1983]  & (\all_features[1982]  | (~new_n17860_ & \all_features[1981] ));
  assign new_n17880_ = \all_features[1983]  & \all_features[1982]  & ~new_n17881_ & new_n17862_;
  assign new_n17881_ = ~\all_features[1978]  & ~\all_features[1979]  & ~\all_features[1980]  & ~\all_features[1981]  & (~\all_features[1977]  | ~\all_features[1976] );
  assign new_n17882_ = ~\all_features[1979]  & ~\all_features[1980]  & (~\all_features[1978]  | new_n17861_);
  assign new_n17883_ = ~new_n17871_ & ~new_n17876_;
  assign new_n17884_ = ~new_n17873_ & ~new_n17874_;
  assign new_n17885_ = ~new_n17875_ & ~new_n17865_;
  assign new_n17886_ = new_n17884_ & ~new_n17887_ & new_n17883_;
  assign new_n17887_ = ~new_n17875_ & ~new_n17865_ & ~new_n17867_ & ~new_n17869_ & (~new_n17880_ | ~new_n17879_);
  assign new_n17888_ = new_n17885_ & new_n17884_ & ~new_n17876_ & ~new_n17869_ & ~new_n17871_ & ~new_n17867_;
  assign new_n17889_ = ~new_n6566_ & (~new_n6563_ | new_n6534_);
  assign new_n17890_ = ~new_n17897_ & (new_n17933_ | ((new_n17891_ | new_n17934_) & (~new_n17936_ | ~new_n17937_ | ~new_n17934_)));
  assign new_n17891_ = (new_n15167_ | ~new_n17896_ | new_n6766_) & (new_n14955_ | new_n14985_ | ~new_n17892_ | (new_n17896_ & ~new_n6766_));
  assign new_n17892_ = ~new_n14980_ & (new_n14979_ | (~new_n14978_ & (new_n14976_ | new_n17893_)));
  assign new_n17893_ = ~new_n14974_ & (new_n14964_ | (~new_n14966_ & (new_n14967_ | (~new_n17894_ & ~new_n14969_))));
  assign new_n17894_ = new_n14972_ & (~new_n14957_ | (new_n14971_ & (new_n17895_ | ~new_n14960_)));
  assign new_n17895_ = \all_features[4166]  & \all_features[4167]  & (\all_features[4165]  | (\all_features[4164]  & (\all_features[4163]  | \all_features[4162] )));
  assign new_n17896_ = ~new_n6738_ & ~new_n6760_;
  assign new_n17897_ = ~new_n17898_ & new_n17933_ & new_n17931_ & (new_n9932_ | (new_n9930_ & new_n9898_));
  assign new_n17898_ = ~new_n17899_ & new_n17927_;
  assign new_n17899_ = ~new_n17926_ & (new_n17919_ | new_n17922_ | new_n17924_ | new_n17925_ | new_n17900_);
  assign new_n17900_ = ~new_n17913_ & ~new_n17918_ & ((~new_n17901_ & new_n17910_) | new_n17917_ | new_n17915_);
  assign new_n17901_ = new_n17902_ & (new_n17908_ | ~\all_features[5053]  | ~\all_features[5054]  | ~\all_features[5055] );
  assign new_n17902_ = \all_features[5055]  & \all_features[5054]  & ~new_n17903_ & new_n17906_;
  assign new_n17903_ = new_n17904_ & ~\all_features[5053]  & ~new_n17905_ & ~\all_features[5052] ;
  assign new_n17904_ = ~\all_features[5050]  & ~\all_features[5051] ;
  assign new_n17905_ = \all_features[5048]  & \all_features[5049] ;
  assign new_n17906_ = \all_features[5055]  & (\all_features[5054]  | (new_n17907_ & (\all_features[5050]  | \all_features[5051]  | \all_features[5049] )));
  assign new_n17907_ = \all_features[5052]  & \all_features[5053] ;
  assign new_n17908_ = ~\all_features[5051]  & ~\all_features[5052]  & (~\all_features[5050]  | new_n17909_);
  assign new_n17909_ = ~\all_features[5048]  & ~\all_features[5049] ;
  assign new_n17910_ = new_n17911_ & new_n17912_;
  assign new_n17911_ = \all_features[5055]  & (\all_features[5054]  | (\all_features[5053]  & (\all_features[5052]  | ~new_n17909_ | ~new_n17904_)));
  assign new_n17912_ = \all_features[5055]  & (\all_features[5053]  | \all_features[5054]  | \all_features[5052] );
  assign new_n17913_ = ~\all_features[5055]  & (~\all_features[5054]  | (~\all_features[5053]  & (new_n17909_ | ~new_n17914_ | ~\all_features[5052] )));
  assign new_n17914_ = \all_features[5050]  & \all_features[5051] ;
  assign new_n17915_ = ~new_n17916_ & ~\all_features[5055] ;
  assign new_n17916_ = \all_features[5053]  & \all_features[5054]  & (\all_features[5052]  | (\all_features[5050]  & \all_features[5051]  & \all_features[5049] ));
  assign new_n17917_ = ~\all_features[5055]  & (~\all_features[5054]  | ~new_n17905_ | ~new_n17907_ | ~new_n17914_);
  assign new_n17918_ = ~\all_features[5055]  & (~\all_features[5054]  | (~\all_features[5052]  & ~\all_features[5053]  & ~new_n17914_));
  assign new_n17919_ = ~new_n17918_ & (new_n17913_ | (~new_n17915_ & (new_n17917_ | new_n17920_)));
  assign new_n17920_ = new_n17912_ & (~new_n17911_ | (~new_n17921_ & new_n17906_));
  assign new_n17921_ = ~\all_features[5053]  & \all_features[5054]  & \all_features[5055]  & (\all_features[5052]  ? new_n17904_ : (new_n17905_ | ~new_n17904_));
  assign new_n17922_ = new_n17923_ & (~\all_features[5053]  | (~\all_features[5052]  & (~\all_features[5051]  | (~\all_features[5050]  & ~\all_features[5049] ))));
  assign new_n17923_ = ~\all_features[5054]  & ~\all_features[5055] ;
  assign new_n17924_ = new_n17923_ & (~\all_features[5051]  | ~new_n17907_ | (~\all_features[5050]  & ~new_n17905_));
  assign new_n17925_ = ~\all_features[5053]  & new_n17923_ & ((~\all_features[5050]  & new_n17909_) | ~\all_features[5052]  | ~\all_features[5051] );
  assign new_n17926_ = ~\all_features[5055]  & ~\all_features[5054]  & ~\all_features[5053]  & ~\all_features[5051]  & ~\all_features[5052] ;
  assign new_n17927_ = new_n17922_ | ~new_n17929_ | ((new_n17915_ | ~new_n17930_) & (new_n17928_ | new_n17924_));
  assign new_n17928_ = ~new_n17913_ & ~new_n17915_ & ~new_n17917_ & ~new_n17918_ & (~new_n17910_ | ~new_n17902_);
  assign new_n17929_ = ~new_n17925_ & ~new_n17926_;
  assign new_n17930_ = ~new_n17924_ & ~new_n17918_ & ~new_n17913_ & ~new_n17917_;
  assign new_n17931_ = ~new_n10871_ & new_n17932_;
  assign new_n17932_ = ~new_n10861_ & ~new_n10868_;
  assign new_n17933_ = new_n13170_ & new_n13196_;
  assign new_n17934_ = ~new_n17935_ & ~new_n12001_;
  assign new_n17935_ = new_n12002_ & new_n11978_;
  assign new_n17936_ = new_n7602_ & (~new_n7627_ | ~new_n7631_);
  assign new_n17937_ = new_n17938_ & (~new_n17963_ | (~new_n17968_ & ~new_n17957_));
  assign new_n17938_ = ~new_n17939_ & ~new_n17961_;
  assign new_n17939_ = new_n17956_ & ~new_n17960_ & ~new_n17940_ & ~new_n17959_;
  assign new_n17940_ = new_n17944_ & (~new_n17953_ | ~new_n17955_ | ~new_n17941_ | ~new_n17952_);
  assign new_n17941_ = \all_features[3719]  & (\all_features[3718]  | new_n17942_);
  assign new_n17942_ = \all_features[3717]  & (\all_features[3714]  | \all_features[3715]  | \all_features[3716]  | ~new_n17943_);
  assign new_n17943_ = ~\all_features[3712]  & ~\all_features[3713] ;
  assign new_n17944_ = ~new_n17950_ & ~new_n17949_ & ~new_n17945_ & ~new_n17947_;
  assign new_n17945_ = ~\all_features[3719]  & (~\all_features[3718]  | (~\all_features[3717]  & (new_n17943_ | ~new_n17946_ | ~\all_features[3716] )));
  assign new_n17946_ = \all_features[3714]  & \all_features[3715] ;
  assign new_n17947_ = ~new_n17948_ & ~\all_features[3719] ;
  assign new_n17948_ = \all_features[3717]  & \all_features[3718]  & (\all_features[3716]  | (\all_features[3714]  & \all_features[3715]  & \all_features[3713] ));
  assign new_n17949_ = ~\all_features[3719]  & (~\all_features[3718]  | (~\all_features[3716]  & ~\all_features[3717]  & ~new_n17946_));
  assign new_n17950_ = ~\all_features[3719]  & (~new_n17946_ | ~\all_features[3712]  | ~\all_features[3713]  | ~\all_features[3718]  | ~new_n17951_);
  assign new_n17951_ = \all_features[3716]  & \all_features[3717] ;
  assign new_n17952_ = \all_features[3719]  & (\all_features[3718]  | (new_n17951_ & (\all_features[3714]  | \all_features[3715]  | \all_features[3713] )));
  assign new_n17953_ = \all_features[3719]  & ~new_n17954_ & \all_features[3718] ;
  assign new_n17954_ = ~\all_features[3714]  & ~\all_features[3715]  & ~\all_features[3716]  & ~\all_features[3717]  & (~\all_features[3713]  | ~\all_features[3712] );
  assign new_n17955_ = \all_features[3719]  & (\all_features[3717]  | \all_features[3718]  | \all_features[3716] );
  assign new_n17956_ = ~new_n17957_ & (\all_features[3715]  | \all_features[3716]  | \all_features[3717]  | \all_features[3718]  | \all_features[3719] );
  assign new_n17957_ = ~\all_features[3717]  & new_n17958_ & ((~\all_features[3714]  & new_n17943_) | ~\all_features[3716]  | ~\all_features[3715] );
  assign new_n17958_ = ~\all_features[3718]  & ~\all_features[3719] ;
  assign new_n17959_ = new_n17958_ & (~\all_features[3717]  | (~\all_features[3716]  & (~\all_features[3715]  | (~\all_features[3714]  & ~\all_features[3713] ))));
  assign new_n17960_ = new_n17958_ & (~new_n17951_ | ~\all_features[3715]  | (~\all_features[3714]  & (~\all_features[3712]  | ~\all_features[3713] )));
  assign new_n17961_ = new_n17962_ & new_n17956_ & ~new_n17947_ & ~new_n17959_;
  assign new_n17962_ = ~new_n17960_ & ~new_n17950_ & ~new_n17945_ & ~new_n17949_;
  assign new_n17963_ = new_n17964_ & (\all_features[3715]  | \all_features[3716]  | \all_features[3717]  | \all_features[3718]  | \all_features[3719] );
  assign new_n17964_ = new_n17956_ & (new_n17960_ | new_n17959_ | (~new_n17945_ & ~new_n17949_ & ~new_n17965_));
  assign new_n17965_ = ~new_n17950_ & ~new_n17947_ & (~new_n17955_ | new_n17966_ | ~new_n17941_);
  assign new_n17966_ = ~new_n17954_ & new_n17952_ & \all_features[3718]  & \all_features[3719]  & (~\all_features[3717]  | new_n17967_);
  assign new_n17967_ = ~\all_features[3715]  & ~\all_features[3716]  & (~\all_features[3714]  | new_n17943_);
  assign new_n17968_ = ~new_n17959_ & (new_n17960_ | (~new_n17949_ & (new_n17945_ | (~new_n17947_ & ~new_n17969_))));
  assign new_n17969_ = ~new_n17950_ & (~new_n17955_ | (new_n17941_ & (~new_n17952_ | (~new_n17970_ & new_n17953_))));
  assign new_n17970_ = \all_features[3718]  & \all_features[3719]  & (\all_features[3717]  | (\all_features[3716]  & (\all_features[3715]  | \all_features[3714] )));
  assign new_n17971_ = (new_n17972_ | ~new_n13099_ | new_n13130_) & (new_n18008_ | ~new_n13479_ | (new_n13099_ & ~new_n13130_));
  assign new_n17972_ = (~new_n17737_ & ~new_n17757_) ? ~new_n17974_ : new_n17973_;
  assign new_n17973_ = new_n17176_ & (new_n17154_ | ~new_n17177_);
  assign new_n17974_ = new_n17975_ & new_n17999_;
  assign new_n17975_ = ~new_n17976_ & ~new_n17998_;
  assign new_n17976_ = new_n17977_ & (~new_n17986_ | (new_n17996_ & new_n17997_ & new_n17993_ & new_n17995_));
  assign new_n17977_ = new_n17978_ & ~new_n17982_ & ~new_n17983_;
  assign new_n17978_ = ~new_n17979_ & (\all_features[5659]  | \all_features[5660]  | \all_features[5661]  | \all_features[5662]  | \all_features[5663] );
  assign new_n17979_ = ~\all_features[5661]  & new_n17981_ & ((~\all_features[5658]  & new_n17980_) | ~\all_features[5660]  | ~\all_features[5659] );
  assign new_n17980_ = ~\all_features[5656]  & ~\all_features[5657] ;
  assign new_n17981_ = ~\all_features[5662]  & ~\all_features[5663] ;
  assign new_n17982_ = new_n17981_ & (~\all_features[5661]  | (~\all_features[5660]  & (~\all_features[5659]  | (~\all_features[5658]  & ~\all_features[5657] ))));
  assign new_n17983_ = new_n17981_ & (~\all_features[5659]  | ~new_n17984_ | (~\all_features[5658]  & ~new_n17985_));
  assign new_n17984_ = \all_features[5660]  & \all_features[5661] ;
  assign new_n17985_ = \all_features[5656]  & \all_features[5657] ;
  assign new_n17986_ = ~new_n17992_ & ~new_n17991_ & ~new_n17987_ & ~new_n17989_;
  assign new_n17987_ = ~\all_features[5663]  & (~\all_features[5662]  | (~\all_features[5661]  & (new_n17980_ | ~new_n17988_ | ~\all_features[5660] )));
  assign new_n17988_ = \all_features[5658]  & \all_features[5659] ;
  assign new_n17989_ = ~new_n17990_ & ~\all_features[5663] ;
  assign new_n17990_ = \all_features[5661]  & \all_features[5662]  & (\all_features[5660]  | (\all_features[5658]  & \all_features[5659]  & \all_features[5657] ));
  assign new_n17991_ = ~\all_features[5663]  & (~\all_features[5662]  | ~new_n17984_ | ~new_n17985_ | ~new_n17988_);
  assign new_n17992_ = ~\all_features[5663]  & (~\all_features[5662]  | (~\all_features[5660]  & ~\all_features[5661]  & ~new_n17988_));
  assign new_n17993_ = \all_features[5663]  & (\all_features[5662]  | (\all_features[5661]  & (\all_features[5660]  | ~new_n17980_ | ~new_n17994_)));
  assign new_n17994_ = ~\all_features[5658]  & ~\all_features[5659] ;
  assign new_n17995_ = \all_features[5663]  & (\all_features[5662]  | (new_n17984_ & (\all_features[5658]  | \all_features[5659]  | \all_features[5657] )));
  assign new_n17996_ = \all_features[5662]  & \all_features[5663]  & (\all_features[5660]  | \all_features[5661]  | new_n17985_ | ~new_n17994_);
  assign new_n17997_ = \all_features[5663]  & (\all_features[5661]  | \all_features[5662]  | \all_features[5660] );
  assign new_n17998_ = new_n17977_ & new_n17986_;
  assign new_n17999_ = ~new_n18000_ & ~new_n18004_;
  assign new_n18000_ = new_n17978_ & (new_n17983_ | new_n17982_ | (~new_n17987_ & ~new_n17992_ & ~new_n18001_));
  assign new_n18001_ = ~new_n17991_ & ~new_n17989_ & (~new_n17997_ | ~new_n17993_ | new_n18002_);
  assign new_n18002_ = new_n17995_ & new_n17996_ & (new_n18003_ | ~\all_features[5661]  | ~\all_features[5662]  | ~\all_features[5663] );
  assign new_n18003_ = ~\all_features[5659]  & ~\all_features[5660]  & (~\all_features[5658]  | new_n17980_);
  assign new_n18004_ = ~new_n18005_ & (\all_features[5659]  | \all_features[5660]  | \all_features[5661]  | \all_features[5662]  | \all_features[5663] );
  assign new_n18005_ = ~new_n17979_ & (new_n17982_ | (~new_n17983_ & (new_n17992_ | (~new_n17987_ & ~new_n18006_))));
  assign new_n18006_ = ~new_n17989_ & (new_n17991_ | (new_n17997_ & (~new_n17993_ | (~new_n18007_ & new_n17995_))));
  assign new_n18007_ = ~\all_features[5661]  & \all_features[5662]  & \all_features[5663]  & (\all_features[5660]  ? new_n17994_ : (new_n17985_ | ~new_n17994_));
  assign new_n18008_ = ~new_n13506_ & ~new_n13510_;
  assign new_n18009_ = ~new_n18010_ & new_n18103_;
  assign new_n18010_ = new_n18011_ & new_n18090_ & (~new_n18098_ | (~new_n18099_ & new_n16101_) | (~new_n18101_ & ~new_n16101_));
  assign new_n18011_ = (~new_n18012_ | new_n18079_) & (new_n18015_ | (new_n18044_ ? ~new_n18040_ : ~new_n18080_));
  assign new_n18012_ = ~new_n18039_ & new_n18013_;
  assign new_n18013_ = ~new_n18014_ & new_n18015_;
  assign new_n18014_ = ~new_n8434_ & (~new_n8412_ | ~new_n8437_);
  assign new_n18015_ = ~new_n18035_ & (new_n18016_ | new_n18037_ | new_n18038_);
  assign new_n18016_ = ~new_n18034_ & new_n18029_ & (~new_n18019_ | ~new_n18023_) & (new_n18017_ | new_n18032_);
  assign new_n18017_ = ~new_n18027_ & ~new_n18018_ & ~new_n18025_;
  assign new_n18018_ = new_n18019_ & (~new_n18023_ | (~new_n18022_ & \all_features[5333]  & \all_features[5334]  & \all_features[5335] ));
  assign new_n18019_ = \all_features[5335]  & (\all_features[5334]  | (\all_features[5333]  & (\all_features[5332]  | ~new_n18021_ | ~new_n18020_)));
  assign new_n18020_ = ~\all_features[5328]  & ~\all_features[5329] ;
  assign new_n18021_ = ~\all_features[5330]  & ~\all_features[5331] ;
  assign new_n18022_ = ~\all_features[5331]  & ~\all_features[5332]  & (~\all_features[5330]  | new_n18020_);
  assign new_n18023_ = \all_features[5334]  & \all_features[5335]  & (\all_features[5332]  | \all_features[5333]  | new_n18024_ | ~new_n18021_);
  assign new_n18024_ = \all_features[5328]  & \all_features[5329] ;
  assign new_n18025_ = ~new_n18026_ & ~\all_features[5335] ;
  assign new_n18026_ = \all_features[5333]  & \all_features[5334]  & (\all_features[5332]  | (\all_features[5330]  & \all_features[5331]  & \all_features[5329] ));
  assign new_n18027_ = ~\all_features[5335]  & (~new_n18028_ | ~\all_features[5332]  | ~\all_features[5333]  | ~\all_features[5334]  | ~new_n18024_);
  assign new_n18028_ = \all_features[5330]  & \all_features[5331] ;
  assign new_n18029_ = ~new_n18033_ & ~new_n18032_ & ~new_n18027_ & ~new_n18025_ & ~new_n18030_;
  assign new_n18030_ = new_n18031_ & (~\all_features[5333]  | (~\all_features[5332]  & (~\all_features[5331]  | (~\all_features[5330]  & ~\all_features[5329] ))));
  assign new_n18031_ = ~\all_features[5334]  & ~\all_features[5335] ;
  assign new_n18032_ = ~\all_features[5335]  & (~\all_features[5334]  | (~\all_features[5332]  & ~\all_features[5333]  & ~new_n18028_));
  assign new_n18033_ = new_n18031_ & (~\all_features[5331]  | ~\all_features[5332]  | ~\all_features[5333]  | (~\all_features[5330]  & ~new_n18024_));
  assign new_n18034_ = ~\all_features[5335]  & (~\all_features[5334]  | (~\all_features[5333]  & (new_n18020_ | ~\all_features[5332]  | ~new_n18028_)));
  assign new_n18035_ = new_n18036_ & ~new_n18038_ & ~new_n18027_ & ~new_n18025_ & ~new_n18030_;
  assign new_n18036_ = ~new_n18033_ & ~new_n18037_ & ~new_n18034_ & ~new_n18032_;
  assign new_n18037_ = ~\all_features[5333]  & new_n18031_ & ((~\all_features[5330]  & new_n18020_) | ~\all_features[5332]  | ~\all_features[5331] );
  assign new_n18038_ = ~\all_features[5335]  & ~\all_features[5334]  & ~\all_features[5333]  & ~\all_features[5331]  & ~\all_features[5332] ;
  assign new_n18039_ = new_n12439_ & new_n12442_;
  assign new_n18040_ = ~new_n18041_ & (new_n17802_ | (~new_n18043_ & new_n17800_));
  assign new_n18041_ = new_n16744_ & ~new_n18042_ & new_n16712_;
  assign new_n18042_ = ~new_n16735_ & ~new_n16740_;
  assign new_n18043_ = ~new_n17771_ & ~new_n17791_;
  assign new_n18044_ = new_n18045_ & ~new_n18071_ & ~new_n18075_;
  assign new_n18045_ = ~new_n18046_ & ~new_n18069_;
  assign new_n18046_ = new_n18064_ & ~new_n18068_ & ~new_n18047_ & ~new_n18067_;
  assign new_n18047_ = ~new_n18060_ & ~new_n18062_ & new_n18055_ & (~new_n18063_ | ~new_n18048_);
  assign new_n18048_ = new_n18054_ & new_n18049_ & new_n18051_;
  assign new_n18049_ = \all_features[4207]  & (\all_features[4206]  | (new_n18050_ & (\all_features[4202]  | \all_features[4203]  | \all_features[4201] )));
  assign new_n18050_ = \all_features[4204]  & \all_features[4205] ;
  assign new_n18051_ = \all_features[4206]  & \all_features[4207]  & (\all_features[4204]  | \all_features[4205]  | new_n18052_ | ~new_n18053_);
  assign new_n18052_ = \all_features[4200]  & \all_features[4201] ;
  assign new_n18053_ = ~\all_features[4202]  & ~\all_features[4203] ;
  assign new_n18054_ = \all_features[4207]  & (\all_features[4205]  | \all_features[4206]  | \all_features[4204] );
  assign new_n18055_ = ~new_n18056_ & ~new_n18058_;
  assign new_n18056_ = ~\all_features[4207]  & (~\all_features[4206]  | (~\all_features[4204]  & ~\all_features[4205]  & ~new_n18057_));
  assign new_n18057_ = \all_features[4202]  & \all_features[4203] ;
  assign new_n18058_ = ~new_n18059_ & ~\all_features[4207] ;
  assign new_n18059_ = \all_features[4205]  & \all_features[4206]  & (\all_features[4204]  | (\all_features[4202]  & \all_features[4203]  & \all_features[4201] ));
  assign new_n18060_ = ~\all_features[4207]  & (~\all_features[4206]  | (~\all_features[4205]  & (new_n18061_ | ~new_n18057_ | ~\all_features[4204] )));
  assign new_n18061_ = ~\all_features[4200]  & ~\all_features[4201] ;
  assign new_n18062_ = ~\all_features[4207]  & (~\all_features[4206]  | ~new_n18052_ | ~new_n18050_ | ~new_n18057_);
  assign new_n18063_ = \all_features[4207]  & (\all_features[4206]  | (\all_features[4205]  & (\all_features[4204]  | ~new_n18053_ | ~new_n18061_)));
  assign new_n18064_ = ~new_n18065_ & (\all_features[4203]  | \all_features[4204]  | \all_features[4205]  | \all_features[4206]  | \all_features[4207] );
  assign new_n18065_ = ~\all_features[4205]  & new_n18066_ & ((~\all_features[4202]  & new_n18061_) | ~\all_features[4204]  | ~\all_features[4203] );
  assign new_n18066_ = ~\all_features[4206]  & ~\all_features[4207] ;
  assign new_n18067_ = new_n18066_ & (~\all_features[4205]  | (~\all_features[4204]  & (~\all_features[4203]  | (~\all_features[4202]  & ~\all_features[4201] ))));
  assign new_n18068_ = new_n18066_ & (~\all_features[4203]  | ~new_n18050_ | (~\all_features[4202]  & ~new_n18052_));
  assign new_n18069_ = new_n18064_ & new_n18055_ & new_n18070_ & ~new_n18060_ & ~new_n18062_;
  assign new_n18070_ = ~new_n18067_ & ~new_n18068_;
  assign new_n18071_ = ~new_n18072_ & (\all_features[4203]  | \all_features[4204]  | \all_features[4205]  | \all_features[4206]  | \all_features[4207] );
  assign new_n18072_ = ~new_n18065_ & (new_n18067_ | (~new_n18068_ & (new_n18056_ | (~new_n18073_ & ~new_n18060_))));
  assign new_n18073_ = ~new_n18058_ & (new_n18062_ | (new_n18054_ & (~new_n18063_ | (~new_n18074_ & new_n18049_))));
  assign new_n18074_ = ~\all_features[4205]  & \all_features[4206]  & \all_features[4207]  & (\all_features[4204]  ? new_n18053_ : (new_n18052_ | ~new_n18053_));
  assign new_n18075_ = new_n18064_ & (~new_n18070_ | (~new_n18076_ & ~new_n18056_ & ~new_n18060_));
  assign new_n18076_ = ~new_n18058_ & ~new_n18062_ & (~new_n18054_ | ~new_n18063_ | new_n18077_);
  assign new_n18077_ = new_n18049_ & new_n18051_ & (new_n18078_ | ~\all_features[4205]  | ~\all_features[4206]  | ~\all_features[4207] );
  assign new_n18078_ = ~\all_features[4203]  & ~\all_features[4204]  & (~\all_features[4202]  | new_n18061_);
  assign new_n18079_ = ~new_n17964_ & new_n17938_;
  assign new_n18080_ = ~new_n18081_ & new_n14786_;
  assign new_n18081_ = ~new_n18082_ & ~new_n18086_;
  assign new_n18082_ = ~new_n18083_ & (\all_features[4587]  | \all_features[4588]  | \all_features[4589]  | \all_features[4590]  | \all_features[4591] );
  assign new_n18083_ = ~new_n14806_ & (new_n14808_ | (~new_n14809_ & (new_n14799_ | (~new_n14803_ & ~new_n18084_))));
  assign new_n18084_ = ~new_n14797_ & (new_n14804_ | (new_n14795_ & (~new_n14801_ | (~new_n18085_ & new_n14790_))));
  assign new_n18085_ = ~\all_features[4589]  & \all_features[4590]  & \all_features[4591]  & (\all_features[4588]  ? new_n14793_ : (new_n14794_ | ~new_n14793_));
  assign new_n18086_ = new_n14805_ & (~new_n14811_ | (~new_n18087_ & ~new_n14799_ & ~new_n14803_));
  assign new_n18087_ = ~new_n14804_ & ~new_n14797_ & (~new_n14795_ | ~new_n14801_ | new_n18088_);
  assign new_n18088_ = new_n14790_ & new_n14792_ & (new_n18089_ | ~\all_features[4589]  | ~\all_features[4590]  | ~\all_features[4591] );
  assign new_n18089_ = ~\all_features[4587]  & ~\all_features[4588]  & (~\all_features[4586]  | new_n14802_);
  assign new_n18090_ = ~new_n18091_ & ((~new_n18093_ & new_n7221_) | ~new_n18039_ | ~new_n18013_);
  assign new_n18091_ = new_n18092_ & new_n18044_ & ~new_n18015_ & new_n18041_;
  assign new_n18092_ = new_n13503_ & (new_n13480_ | ~new_n18008_);
  assign new_n18093_ = ~new_n7194_ & new_n18094_;
  assign new_n18094_ = ~new_n7218_ & (new_n7217_ | (~new_n7216_ & (new_n7214_ | new_n18095_)));
  assign new_n18095_ = ~new_n7212_ & (new_n7210_ | (~new_n7196_ & (new_n7207_ | (~new_n7209_ & ~new_n18096_))));
  assign new_n18096_ = \all_features[1959]  & ((new_n18097_ & (\all_features[1958]  | \all_features[1957] )) | (~\all_features[1958]  & (\all_features[1957]  ? new_n7200_ : \all_features[1956] )));
  assign new_n18097_ = new_n7203_ & (\all_features[1957]  | ~new_n7206_ | (~new_n7205_ & ~\all_features[1956]  & new_n7201_) | (\all_features[1956]  & ~new_n7201_));
  assign new_n18098_ = new_n18014_ & new_n18015_;
  assign new_n18099_ = new_n18100_ & new_n8268_;
  assign new_n18100_ = ~new_n16412_ & ~new_n8295_;
  assign new_n18101_ = ~new_n18102_ & ~new_n11884_;
  assign new_n18102_ = new_n11861_ & new_n11887_;
  assign new_n18103_ = new_n18104_ & (~new_n18079_ | ~new_n18012_);
  assign new_n18104_ = new_n18105_ & (~new_n18098_ | (new_n18099_ & new_n16101_) | (new_n18101_ & ~new_n16101_));
  assign new_n18105_ = new_n18015_ | ((new_n18092_ | ~new_n18041_ | ~new_n18044_) & (new_n18080_ | new_n18044_));
  assign new_n18106_ = (new_n8268_ | ~new_n18109_ | (~new_n6355_ & new_n16279_)) & new_n18107_ & (~new_n18111_ | new_n6355_ | ~new_n16279_);
  assign new_n18107_ = ~new_n9163_ & (~new_n9159_ | ~new_n18108_);
  assign new_n18108_ = new_n9135_ & new_n9165_;
  assign new_n18109_ = new_n16909_ & new_n18110_;
  assign new_n18110_ = new_n13210_ & new_n13234_;
  assign new_n18111_ = new_n10001_ & new_n8854_;
  assign new_n18112_ = new_n18113_ ? (new_n18372_ ^ new_n18908_) : (~new_n18372_ ^ new_n18908_);
  assign new_n18113_ = new_n18114_ ? (~new_n18338_ ^ new_n18339_) : (new_n18338_ ^ new_n18339_);
  assign new_n18114_ = new_n18115_ ? (new_n18182_ ^ new_n18337_) : (~new_n18182_ ^ new_n18337_);
  assign new_n18115_ = ~new_n18116_ & new_n18179_;
  assign new_n18116_ = ~new_n18159_ & new_n18117_ & (~new_n18173_ | (~new_n18177_ & new_n18174_) | (new_n18175_ & ~new_n18174_));
  assign new_n18117_ = new_n11202_ | ((new_n18153_ | new_n18158_ | new_n10513_ | new_n16956_) & (new_n18118_ | ~new_n16956_));
  assign new_n18118_ = new_n8740_ ? new_n18119_ : ~new_n18152_;
  assign new_n18119_ = new_n18120_ & (new_n18138_ | (~new_n18149_ & ~new_n18137_));
  assign new_n18120_ = new_n18121_ & (~new_n18136_ | (new_n18132_ & (new_n18146_ | new_n18140_ | new_n18143_)));
  assign new_n18121_ = ~new_n18132_ | ~new_n18136_;
  assign new_n18123_ = \all_features[4191]  & (\all_features[4190]  | new_n18124_);
  assign new_n18124_ = \all_features[4189]  & (\all_features[4186]  | \all_features[4187]  | \all_features[4188]  | ~new_n18125_);
  assign new_n18125_ = ~\all_features[4184]  & ~\all_features[4185] ;
  assign new_n18126_ = \all_features[4191]  & ~new_n18127_ & \all_features[4190] ;
  assign new_n18127_ = ~\all_features[4189]  & ~\all_features[4188]  & ~\all_features[4187]  & ~new_n18128_ & ~\all_features[4186] ;
  assign new_n18128_ = \all_features[4184]  & \all_features[4185] ;
  assign new_n18129_ = \all_features[4191]  & (\all_features[4190]  | (new_n18130_ & (\all_features[4186]  | \all_features[4187]  | \all_features[4185] )));
  assign new_n18130_ = \all_features[4188]  & \all_features[4189] ;
  assign new_n18131_ = \all_features[4191]  & (\all_features[4189]  | \all_features[4190]  | \all_features[4188] );
  assign new_n18132_ = ~new_n18133_ & ~new_n18135_;
  assign new_n18133_ = new_n18134_ & (~\all_features[4189]  | (~\all_features[4188]  & (~\all_features[4187]  | (~\all_features[4186]  & ~\all_features[4185] ))));
  assign new_n18134_ = ~\all_features[4190]  & ~\all_features[4191] ;
  assign new_n18135_ = new_n18134_ & (~\all_features[4187]  | ~new_n18130_ | (~\all_features[4186]  & ~new_n18128_));
  assign new_n18136_ = ~new_n18137_ & ~new_n18138_;
  assign new_n18137_ = ~\all_features[4189]  & new_n18134_ & ((~\all_features[4186]  & new_n18125_) | ~\all_features[4188]  | ~\all_features[4187] );
  assign new_n18138_ = ~\all_features[4191]  & ~\all_features[4190]  & ~\all_features[4189]  & ~\all_features[4187]  & ~\all_features[4188] ;
  assign new_n18139_ = ~new_n18140_ & ~new_n18142_;
  assign new_n18140_ = ~\all_features[4191]  & (~\all_features[4190]  | (~\all_features[4188]  & ~\all_features[4189]  & ~new_n18141_));
  assign new_n18141_ = \all_features[4186]  & \all_features[4187] ;
  assign new_n18142_ = ~\all_features[4191]  & (~\all_features[4190]  | ~new_n18128_ | ~new_n18130_ | ~new_n18141_);
  assign new_n18143_ = ~\all_features[4191]  & (~\all_features[4190]  | (~\all_features[4189]  & (new_n18125_ | ~new_n18141_ | ~\all_features[4188] )));
  assign new_n18144_ = ~new_n18145_ & ~\all_features[4191] ;
  assign new_n18145_ = \all_features[4189]  & \all_features[4190]  & (\all_features[4188]  | (\all_features[4186]  & \all_features[4187]  & \all_features[4185] ));
  assign new_n18146_ = ~new_n18142_ & ~new_n18144_ & (~new_n18131_ | new_n18147_ | ~new_n18123_);
  assign new_n18147_ = ~new_n18127_ & new_n18129_ & \all_features[4190]  & \all_features[4191]  & (~\all_features[4189]  | new_n18148_);
  assign new_n18148_ = ~\all_features[4187]  & ~\all_features[4188]  & (~\all_features[4186]  | new_n18125_);
  assign new_n18149_ = ~new_n18133_ & (new_n18135_ | (~new_n18140_ & (new_n18143_ | (~new_n18150_ & ~new_n18144_))));
  assign new_n18150_ = ~new_n18142_ & (~new_n18131_ | (new_n18123_ & (~new_n18129_ | (~new_n18151_ & new_n18126_))));
  assign new_n18151_ = \all_features[4190]  & \all_features[4191]  & (\all_features[4189]  | (\all_features[4188]  & (\all_features[4187]  | \all_features[4186] )));
  assign new_n18152_ = ~new_n9835_ & new_n10637_;
  assign new_n18153_ = ~new_n18154_ & new_n13450_;
  assign new_n18154_ = ~new_n18155_ & (\all_features[3107]  | \all_features[3108]  | \all_features[3109]  | \all_features[3110]  | \all_features[3111] );
  assign new_n18155_ = ~new_n13472_ & (new_n13470_ | (~new_n13468_ & (new_n13473_ | (~new_n18156_ & ~new_n13474_))));
  assign new_n18156_ = ~new_n13464_ & (new_n13462_ | (new_n13466_ & (~new_n13461_ | (~new_n18157_ & new_n13454_))));
  assign new_n18157_ = ~\all_features[3109]  & \all_features[3110]  & \all_features[3111]  & (\all_features[3108]  ? new_n13460_ : (new_n13459_ | ~new_n13460_));
  assign new_n18158_ = new_n10491_ & new_n10516_;
  assign new_n18159_ = new_n18160_ & new_n18162_;
  assign new_n18160_ = (new_n16518_ & new_n18161_ & (new_n16515_ | (new_n16487_ & new_n16508_))) | (~new_n6389_ & ~new_n18161_);
  assign new_n18161_ = ~new_n8356_ & new_n12598_;
  assign new_n18162_ = ~new_n18163_ & new_n11202_;
  assign new_n18163_ = new_n12624_ & (new_n12601_ | new_n18164_);
  assign new_n18164_ = new_n18165_ & new_n18169_;
  assign new_n18165_ = ~new_n18166_ & (\all_features[4571]  | \all_features[4572]  | \all_features[4573]  | \all_features[4574]  | \all_features[4575] );
  assign new_n18166_ = ~new_n12620_ & (new_n12622_ | (~new_n12623_ & (new_n12613_ | (~new_n12617_ & ~new_n18167_))));
  assign new_n18167_ = ~new_n12611_ & (new_n12618_ | (new_n12609_ & (~new_n12615_ | (~new_n18168_ & new_n12604_))));
  assign new_n18168_ = ~\all_features[4573]  & \all_features[4574]  & \all_features[4575]  & (\all_features[4572]  ? new_n12607_ : (new_n12608_ | ~new_n12607_));
  assign new_n18169_ = new_n12619_ & (~new_n12625_ | (~new_n18170_ & ~new_n12613_ & ~new_n12617_));
  assign new_n18170_ = ~new_n12618_ & ~new_n12611_ & (~new_n12609_ | ~new_n12615_ | new_n18171_);
  assign new_n18171_ = new_n12604_ & new_n12606_ & (new_n18172_ | ~\all_features[4573]  | ~\all_features[4574]  | ~\all_features[4575] );
  assign new_n18172_ = ~\all_features[4571]  & ~\all_features[4572]  & (~\all_features[4570]  | new_n12616_);
  assign new_n18173_ = new_n11202_ & new_n18163_;
  assign new_n18174_ = ~new_n12049_ & ~new_n12081_;
  assign new_n18175_ = new_n7591_ & new_n18176_;
  assign new_n18176_ = ~new_n7376_ & ~new_n7396_;
  assign new_n18177_ = new_n18178_ & (~new_n12747_ | ~new_n12739_);
  assign new_n18178_ = ~new_n12338_ & ~new_n12753_;
  assign new_n18179_ = ~new_n18180_ & new_n18181_ & (~new_n18173_ | (new_n18177_ & new_n18174_) | (~new_n18175_ & ~new_n18174_));
  assign new_n18180_ = ~new_n18160_ & new_n18162_;
  assign new_n18181_ = new_n11202_ | (new_n16956_ ? (new_n8740_ ? ~new_n18119_ : new_n18152_) : ~new_n18153_);
  assign new_n18182_ = ~new_n18183_ & new_n18336_;
  assign new_n18183_ = ~new_n18327_ & ~new_n18325_ & new_n18184_ & (~new_n16658_ | ~new_n18335_);
  assign new_n18184_ = ~new_n18185_ & (~new_n18187_ | (~new_n18258_ & new_n18323_ & new_n18289_) | (~new_n18222_ & ~new_n18289_));
  assign new_n18185_ = new_n18186_ & new_n18193_;
  assign new_n18186_ = ~new_n18191_ & ~new_n18187_ & ~new_n18189_;
  assign new_n18187_ = ~new_n18188_ & new_n13348_;
  assign new_n18188_ = new_n12269_ & new_n12294_;
  assign new_n18189_ = ~new_n17218_ & new_n18190_;
  assign new_n18190_ = ~new_n17244_ & ~new_n17247_;
  assign new_n18191_ = new_n18192_ & new_n10801_;
  assign new_n18192_ = new_n10778_ & new_n10834_;
  assign new_n18193_ = new_n18221_ & (new_n18217_ | new_n18194_);
  assign new_n18194_ = new_n18215_ & ~new_n18195_ & new_n18211_;
  assign new_n18195_ = ~new_n18205_ & ~new_n18207_ & ~new_n18208_ & ~new_n18210_ & (~new_n18200_ | ~new_n18196_);
  assign new_n18196_ = \all_features[5327]  & (\all_features[5326]  | (~new_n18197_ & \all_features[5325] ));
  assign new_n18197_ = new_n18198_ & ~\all_features[5324]  & new_n18199_;
  assign new_n18198_ = ~\all_features[5320]  & ~\all_features[5321] ;
  assign new_n18199_ = ~\all_features[5322]  & ~\all_features[5323] ;
  assign new_n18200_ = \all_features[5327]  & \all_features[5326]  & ~new_n18203_ & new_n18201_;
  assign new_n18201_ = \all_features[5327]  & (\all_features[5326]  | (new_n18202_ & (\all_features[5322]  | \all_features[5323]  | \all_features[5321] )));
  assign new_n18202_ = \all_features[5324]  & \all_features[5325] ;
  assign new_n18203_ = new_n18199_ & ~\all_features[5325]  & ~new_n18204_ & ~\all_features[5324] ;
  assign new_n18204_ = \all_features[5320]  & \all_features[5321] ;
  assign new_n18205_ = ~\all_features[5327]  & (~\all_features[5326]  | (~\all_features[5324]  & ~\all_features[5325]  & ~new_n18206_));
  assign new_n18206_ = \all_features[5322]  & \all_features[5323] ;
  assign new_n18207_ = ~\all_features[5327]  & (~\all_features[5326]  | (~\all_features[5325]  & (new_n18198_ | ~\all_features[5324]  | ~new_n18206_)));
  assign new_n18208_ = ~new_n18209_ & ~\all_features[5327] ;
  assign new_n18209_ = \all_features[5325]  & \all_features[5326]  & (\all_features[5324]  | (\all_features[5322]  & \all_features[5323]  & \all_features[5321] ));
  assign new_n18210_ = ~\all_features[5327]  & (~\all_features[5326]  | ~new_n18206_ | ~new_n18204_ | ~new_n18202_);
  assign new_n18211_ = ~new_n18212_ & ~new_n18214_;
  assign new_n18212_ = new_n18213_ & (~\all_features[5323]  | ~new_n18202_ | (~\all_features[5322]  & ~new_n18204_));
  assign new_n18213_ = ~\all_features[5326]  & ~\all_features[5327] ;
  assign new_n18214_ = new_n18213_ & (~\all_features[5325]  | (~\all_features[5324]  & (~\all_features[5323]  | (~\all_features[5322]  & ~\all_features[5321] ))));
  assign new_n18215_ = ~new_n18216_ & (\all_features[5323]  | \all_features[5324]  | \all_features[5325]  | \all_features[5326]  | \all_features[5327] );
  assign new_n18216_ = ~\all_features[5325]  & new_n18213_ & ((~\all_features[5322]  & new_n18198_) | ~\all_features[5324]  | ~\all_features[5323] );
  assign new_n18217_ = new_n18215_ & (~new_n18211_ | (new_n18220_ & (new_n18218_ | new_n18208_ | new_n18210_)));
  assign new_n18218_ = new_n18196_ & (~new_n18200_ | (~new_n18219_ & \all_features[5325]  & \all_features[5326]  & \all_features[5327] ));
  assign new_n18219_ = ~\all_features[5323]  & ~\all_features[5324]  & (~\all_features[5322]  | new_n18198_);
  assign new_n18220_ = ~new_n18205_ & ~new_n18207_;
  assign new_n18221_ = new_n18211_ & new_n18220_ & new_n18215_ & ~new_n18208_ & ~new_n18210_;
  assign new_n18222_ = ~new_n14384_ & new_n18223_;
  assign new_n18223_ = new_n18224_ & ~new_n18253_ & ~new_n18256_;
  assign new_n18224_ = ~new_n18225_ & ~new_n18249_;
  assign new_n18225_ = new_n18240_ & (~new_n18245_ | (~new_n18243_ & ~new_n18226_ & ~new_n18248_));
  assign new_n18226_ = ~new_n18238_ & ~new_n18236_ & (~new_n18239_ | ~new_n18235_ | new_n18227_);
  assign new_n18227_ = new_n18228_ & new_n18230_ & (new_n18233_ | ~\all_features[3789]  | ~\all_features[3790]  | ~\all_features[3791] );
  assign new_n18228_ = \all_features[3791]  & (\all_features[3790]  | (new_n18229_ & (\all_features[3786]  | \all_features[3787]  | \all_features[3785] )));
  assign new_n18229_ = \all_features[3788]  & \all_features[3789] ;
  assign new_n18230_ = \all_features[3790]  & \all_features[3791]  & (\all_features[3788]  | \all_features[3789]  | new_n18232_ | ~new_n18231_);
  assign new_n18231_ = ~\all_features[3786]  & ~\all_features[3787] ;
  assign new_n18232_ = \all_features[3784]  & \all_features[3785] ;
  assign new_n18233_ = ~\all_features[3787]  & ~\all_features[3788]  & (~\all_features[3786]  | new_n18234_);
  assign new_n18234_ = ~\all_features[3784]  & ~\all_features[3785] ;
  assign new_n18235_ = \all_features[3791]  & (\all_features[3790]  | (\all_features[3789]  & (\all_features[3788]  | ~new_n18231_ | ~new_n18234_)));
  assign new_n18236_ = ~new_n18237_ & ~\all_features[3791] ;
  assign new_n18237_ = \all_features[3789]  & \all_features[3790]  & (\all_features[3788]  | (\all_features[3786]  & \all_features[3787]  & \all_features[3785] ));
  assign new_n18238_ = ~\all_features[3791]  & (~new_n18232_ | ~\all_features[3786]  | ~\all_features[3787]  | ~\all_features[3790]  | ~new_n18229_);
  assign new_n18239_ = \all_features[3791]  & (\all_features[3789]  | \all_features[3790]  | \all_features[3788] );
  assign new_n18240_ = ~new_n18241_ & (\all_features[3787]  | \all_features[3788]  | \all_features[3789]  | \all_features[3790]  | \all_features[3791] );
  assign new_n18241_ = ~\all_features[3789]  & new_n18242_ & ((~\all_features[3786]  & new_n18234_) | ~\all_features[3788]  | ~\all_features[3787] );
  assign new_n18242_ = ~\all_features[3790]  & ~\all_features[3791] ;
  assign new_n18243_ = ~\all_features[3791]  & (~\all_features[3790]  | new_n18244_);
  assign new_n18244_ = ~\all_features[3789]  & (new_n18234_ | ~\all_features[3787]  | ~\all_features[3788]  | ~\all_features[3786] );
  assign new_n18245_ = ~new_n18246_ & ~new_n18247_;
  assign new_n18246_ = new_n18242_ & (~\all_features[3787]  | ~new_n18229_ | (~new_n18232_ & ~\all_features[3786] ));
  assign new_n18247_ = new_n18242_ & (~\all_features[3789]  | (~\all_features[3788]  & (~\all_features[3787]  | (~\all_features[3786]  & ~\all_features[3785] ))));
  assign new_n18248_ = ~\all_features[3791]  & (~\all_features[3790]  | (~\all_features[3789]  & ~\all_features[3788]  & (~\all_features[3787]  | ~\all_features[3786] )));
  assign new_n18249_ = ~new_n18250_ & (\all_features[3787]  | \all_features[3788]  | \all_features[3789]  | \all_features[3790]  | \all_features[3791] );
  assign new_n18250_ = ~new_n18241_ & (new_n18247_ | (~new_n18246_ & (new_n18248_ | (~new_n18243_ & ~new_n18251_))));
  assign new_n18251_ = ~new_n18236_ & (new_n18238_ | (new_n18239_ & (~new_n18235_ | (~new_n18252_ & new_n18228_))));
  assign new_n18252_ = ~\all_features[3789]  & \all_features[3790]  & \all_features[3791]  & (\all_features[3788]  ? new_n18231_ : (new_n18232_ | ~new_n18231_));
  assign new_n18253_ = new_n18245_ & ~new_n18254_ & new_n18240_;
  assign new_n18254_ = ~new_n18248_ & ~new_n18238_ & ~new_n18236_ & ~new_n18243_ & ~new_n18255_;
  assign new_n18255_ = new_n18239_ & new_n18235_ & new_n18228_ & new_n18230_;
  assign new_n18256_ = new_n18240_ & new_n18257_ & ~new_n18236_ & ~new_n18247_;
  assign new_n18257_ = ~new_n18248_ & ~new_n18246_ & ~new_n18243_ & ~new_n18238_;
  assign new_n18258_ = new_n18259_ & new_n18288_;
  assign new_n18259_ = new_n18260_ & new_n18285_;
  assign new_n18260_ = new_n18283_ & (~new_n18271_ | (new_n18275_ & (~new_n18279_ | new_n18261_)));
  assign new_n18261_ = new_n18262_ & (~new_n18265_ | (~new_n18270_ & \all_features[4821]  & \all_features[4822]  & \all_features[4823] ));
  assign new_n18262_ = \all_features[4823]  & (\all_features[4822]  | (~new_n18263_ & \all_features[4821] ));
  assign new_n18263_ = new_n18264_ & ~\all_features[4820]  & ~\all_features[4818]  & ~\all_features[4819] ;
  assign new_n18264_ = ~\all_features[4816]  & ~\all_features[4817] ;
  assign new_n18265_ = \all_features[4823]  & \all_features[4822]  & ~new_n18268_ & new_n18266_;
  assign new_n18266_ = \all_features[4823]  & (\all_features[4822]  | (new_n18267_ & (\all_features[4818]  | \all_features[4819]  | \all_features[4817] )));
  assign new_n18267_ = \all_features[4820]  & \all_features[4821] ;
  assign new_n18268_ = ~\all_features[4821]  & ~\all_features[4820]  & ~\all_features[4819]  & ~new_n18269_ & ~\all_features[4818] ;
  assign new_n18269_ = \all_features[4816]  & \all_features[4817] ;
  assign new_n18270_ = ~\all_features[4819]  & ~\all_features[4820]  & (~\all_features[4818]  | new_n18264_);
  assign new_n18271_ = ~new_n18272_ & ~new_n18273_;
  assign new_n18272_ = ~\all_features[4822]  & ~\all_features[4823]  & (~\all_features[4819]  | ~new_n18267_ | (~\all_features[4818]  & ~new_n18269_));
  assign new_n18273_ = ~\all_features[4823]  & ~new_n18274_ & ~\all_features[4822] ;
  assign new_n18274_ = \all_features[4821]  & (\all_features[4820]  | (\all_features[4819]  & (\all_features[4818]  | \all_features[4817] )));
  assign new_n18275_ = ~new_n18276_ & ~new_n18278_;
  assign new_n18276_ = ~\all_features[4823]  & (~\all_features[4822]  | (~\all_features[4820]  & ~\all_features[4821]  & ~new_n18277_));
  assign new_n18277_ = \all_features[4818]  & \all_features[4819] ;
  assign new_n18278_ = ~\all_features[4823]  & (~\all_features[4822]  | (~\all_features[4821]  & (new_n18264_ | ~new_n18277_ | ~\all_features[4820] )));
  assign new_n18279_ = ~new_n18280_ & ~new_n18281_;
  assign new_n18280_ = ~\all_features[4823]  & (~\all_features[4822]  | ~new_n18269_ | ~new_n18267_ | ~new_n18277_);
  assign new_n18281_ = ~new_n18282_ & ~\all_features[4823] ;
  assign new_n18282_ = \all_features[4821]  & \all_features[4822]  & (\all_features[4820]  | (\all_features[4818]  & \all_features[4819]  & \all_features[4817] ));
  assign new_n18283_ = ~new_n18284_ | (\all_features[4819]  & \all_features[4820]  & (\all_features[4818]  | ~new_n18264_));
  assign new_n18284_ = ~\all_features[4823]  & ~\all_features[4821]  & ~\all_features[4822] ;
  assign new_n18285_ = new_n18286_ & (new_n18278_ | new_n18281_ | ~new_n18287_ | (new_n18265_ & new_n18262_));
  assign new_n18286_ = new_n18271_ & new_n18283_;
  assign new_n18287_ = ~new_n18276_ & ~new_n18280_;
  assign new_n18288_ = new_n18279_ & new_n18286_ & new_n18275_;
  assign new_n18289_ = new_n18321_ & (~new_n18290_ | (~new_n18317_ & (new_n18316_ | new_n18318_)));
  assign new_n18290_ = new_n18316_ | new_n18317_ | (~new_n18313_ & ~new_n18315_ & ~new_n18309_ & new_n18291_);
  assign new_n18291_ = ~new_n18307_ & ~new_n18308_ & new_n18299_ & (~new_n18304_ | ~new_n18292_);
  assign new_n18292_ = new_n18298_ & new_n18293_ & new_n18296_;
  assign new_n18293_ = \all_features[1039]  & ~new_n18294_ & \all_features[1038] ;
  assign new_n18294_ = ~\all_features[1037]  & ~\all_features[1036]  & ~\all_features[1035]  & ~new_n18295_ & ~\all_features[1034] ;
  assign new_n18295_ = \all_features[1032]  & \all_features[1033] ;
  assign new_n18296_ = \all_features[1039]  & (\all_features[1038]  | (new_n18297_ & (\all_features[1034]  | \all_features[1035]  | \all_features[1033] )));
  assign new_n18297_ = \all_features[1036]  & \all_features[1037] ;
  assign new_n18298_ = \all_features[1039]  & (\all_features[1037]  | \all_features[1038]  | \all_features[1036] );
  assign new_n18299_ = ~new_n18300_ & ~new_n18302_;
  assign new_n18300_ = ~new_n18301_ & ~\all_features[1039] ;
  assign new_n18301_ = \all_features[1037]  & \all_features[1038]  & (\all_features[1036]  | (\all_features[1034]  & \all_features[1035]  & \all_features[1033] ));
  assign new_n18302_ = ~\all_features[1039]  & (~\all_features[1038]  | (~\all_features[1036]  & ~\all_features[1037]  & ~new_n18303_));
  assign new_n18303_ = \all_features[1034]  & \all_features[1035] ;
  assign new_n18304_ = \all_features[1039]  & (\all_features[1038]  | new_n18305_);
  assign new_n18305_ = \all_features[1037]  & (\all_features[1034]  | \all_features[1035]  | \all_features[1036]  | ~new_n18306_);
  assign new_n18306_ = ~\all_features[1032]  & ~\all_features[1033] ;
  assign new_n18307_ = ~\all_features[1039]  & (~\all_features[1038]  | ~new_n18295_ | ~new_n18297_ | ~new_n18303_);
  assign new_n18308_ = ~\all_features[1039]  & (~\all_features[1038]  | (~\all_features[1037]  & (new_n18306_ | ~new_n18303_ | ~\all_features[1036] )));
  assign new_n18309_ = ~new_n18308_ & ~new_n18302_ & (new_n18300_ | new_n18307_ | new_n18310_);
  assign new_n18310_ = new_n18298_ & ~new_n18311_ & new_n18304_;
  assign new_n18311_ = ~new_n18294_ & new_n18296_ & \all_features[1038]  & \all_features[1039]  & (~\all_features[1037]  | new_n18312_);
  assign new_n18312_ = ~\all_features[1035]  & ~\all_features[1036]  & (~\all_features[1034]  | new_n18306_);
  assign new_n18313_ = new_n18314_ & (~\all_features[1035]  | ~new_n18297_ | (~\all_features[1034]  & ~new_n18295_));
  assign new_n18314_ = ~\all_features[1038]  & ~\all_features[1039] ;
  assign new_n18315_ = new_n18314_ & (~\all_features[1037]  | (~\all_features[1036]  & (~\all_features[1035]  | (~\all_features[1034]  & ~\all_features[1033] ))));
  assign new_n18316_ = ~\all_features[1037]  & new_n18314_ & ((~\all_features[1034]  & new_n18306_) | ~\all_features[1036]  | ~\all_features[1035] );
  assign new_n18317_ = ~\all_features[1039]  & ~\all_features[1038]  & ~\all_features[1037]  & ~\all_features[1035]  & ~\all_features[1036] ;
  assign new_n18318_ = ~new_n18315_ & (new_n18313_ | (~new_n18302_ & (new_n18308_ | (~new_n18319_ & ~new_n18300_))));
  assign new_n18319_ = ~new_n18307_ & (~new_n18298_ | (new_n18304_ & (~new_n18296_ | (~new_n18320_ & new_n18293_))));
  assign new_n18320_ = \all_features[1038]  & \all_features[1039]  & (\all_features[1037]  | (\all_features[1036]  & (\all_features[1035]  | \all_features[1034] )));
  assign new_n18321_ = new_n18299_ & new_n18322_ & ~new_n18308_ & ~new_n18316_ & ~new_n18313_ & ~new_n18315_;
  assign new_n18322_ = ~new_n18307_ & ~new_n18317_;
  assign new_n18323_ = new_n8298_ & new_n18324_;
  assign new_n18324_ = ~new_n8344_ & ~new_n8346_;
  assign new_n18325_ = ~new_n18187_ & ((~new_n18326_ & new_n11000_ & new_n18189_) | (~new_n10247_ & new_n18191_ & ~new_n18189_));
  assign new_n18326_ = new_n15195_ & (new_n15172_ | new_n15197_);
  assign new_n18327_ = ~new_n18289_ & new_n18187_ & (new_n18223_ ? new_n14384_ : (~new_n18334_ | new_n18328_));
  assign new_n18328_ = new_n8508_ & new_n18329_;
  assign new_n18329_ = ~new_n8514_ & (new_n8510_ | (~new_n8529_ & (new_n8528_ | (~new_n8524_ & ~new_n18330_))));
  assign new_n18330_ = ~new_n8526_ & (new_n8530_ | (~new_n8532_ & (~new_n18333_ | new_n18331_)));
  assign new_n18331_ = \all_features[3087]  & ((~new_n18332_ & ~\all_features[3085]  & \all_features[3086] ) | (~new_n8519_ & (\all_features[3086]  | (~new_n8517_ & \all_features[3085] ))));
  assign new_n18332_ = (~\all_features[3082]  & ~\all_features[3083]  & ~\all_features[3084]  & (~\all_features[3081]  | ~\all_features[3080] )) | (\all_features[3084]  & (\all_features[3082]  | \all_features[3083] ));
  assign new_n18333_ = \all_features[3087]  & (\all_features[3085]  | \all_features[3086]  | \all_features[3084] );
  assign new_n18334_ = ~new_n8533_ & ~new_n8535_;
  assign new_n18335_ = new_n18326_ & ~new_n18187_ & new_n18189_;
  assign new_n18336_ = (new_n16658_ | ~new_n18335_) & (new_n18193_ | ~new_n18186_);
  assign new_n18337_ = ~new_n17672_ & new_n17806_;
  assign new_n18338_ = new_n17147_ & new_n17286_;
  assign new_n18339_ = new_n18107_ & (~new_n9583_ | (new_n18340_ & (~new_n18368_ | ~new_n18364_)));
  assign new_n18340_ = new_n18363_ | ~new_n18361_ | ((new_n18352_ | new_n18350_) & (new_n18358_ | ~new_n18341_));
  assign new_n18341_ = new_n18342_ & ~new_n18348_ & ~new_n18350_;
  assign new_n18342_ = ~new_n18343_ & ~new_n18347_;
  assign new_n18343_ = ~\all_features[839]  & (~\all_features[838]  | ~new_n18344_ | ~new_n18345_ | ~new_n18346_);
  assign new_n18344_ = \all_features[834]  & \all_features[835] ;
  assign new_n18345_ = \all_features[832]  & \all_features[833] ;
  assign new_n18346_ = \all_features[836]  & \all_features[837] ;
  assign new_n18347_ = ~\all_features[839]  & (~\all_features[838]  | (~\all_features[836]  & ~\all_features[837]  & ~new_n18344_));
  assign new_n18348_ = ~\all_features[839]  & (~\all_features[838]  | (~\all_features[837]  & (new_n18349_ | ~new_n18344_ | ~\all_features[836] )));
  assign new_n18349_ = ~\all_features[832]  & ~\all_features[833] ;
  assign new_n18350_ = new_n18351_ & (~\all_features[835]  | ~new_n18346_ | (~\all_features[834]  & ~new_n18345_));
  assign new_n18351_ = ~\all_features[838]  & ~\all_features[839] ;
  assign new_n18352_ = ~new_n18358_ & ~new_n18348_ & new_n18342_ & (~new_n18360_ | ~new_n18353_);
  assign new_n18353_ = new_n18357_ & new_n18354_ & new_n18355_;
  assign new_n18354_ = \all_features[839]  & (\all_features[838]  | (new_n18346_ & (\all_features[834]  | \all_features[835]  | \all_features[833] )));
  assign new_n18355_ = \all_features[838]  & \all_features[839]  & (\all_features[836]  | \all_features[837]  | new_n18345_ | ~new_n18356_);
  assign new_n18356_ = ~\all_features[834]  & ~\all_features[835] ;
  assign new_n18357_ = \all_features[839]  & (\all_features[837]  | \all_features[838]  | \all_features[836] );
  assign new_n18358_ = ~new_n18359_ & ~\all_features[839] ;
  assign new_n18359_ = \all_features[837]  & \all_features[838]  & (\all_features[836]  | (\all_features[834]  & \all_features[835]  & \all_features[833] ));
  assign new_n18360_ = \all_features[839]  & (\all_features[838]  | (\all_features[837]  & (\all_features[836]  | ~new_n18356_ | ~new_n18349_)));
  assign new_n18361_ = ~new_n18362_ & (\all_features[835]  | \all_features[836]  | \all_features[837]  | \all_features[838]  | \all_features[839] );
  assign new_n18362_ = ~\all_features[837]  & new_n18351_ & ((~\all_features[834]  & new_n18349_) | ~\all_features[836]  | ~\all_features[835] );
  assign new_n18363_ = new_n18351_ & (~\all_features[837]  | (~\all_features[836]  & (~\all_features[835]  | (~\all_features[834]  & ~\all_features[833] ))));
  assign new_n18364_ = new_n18361_ & (new_n18350_ | new_n18363_ | (~new_n18365_ & ~new_n18348_ & ~new_n18347_));
  assign new_n18365_ = ~new_n18358_ & ~new_n18343_ & (~new_n18357_ | ~new_n18360_ | new_n18366_);
  assign new_n18366_ = new_n18354_ & new_n18355_ & (new_n18367_ | ~\all_features[837]  | ~\all_features[838]  | ~\all_features[839] );
  assign new_n18367_ = ~\all_features[835]  & ~\all_features[836]  & (~\all_features[834]  | new_n18349_);
  assign new_n18368_ = ~new_n18369_ & (\all_features[835]  | \all_features[836]  | \all_features[837]  | \all_features[838]  | \all_features[839] );
  assign new_n18369_ = ~new_n18362_ & (new_n18363_ | (~new_n18350_ & (new_n18347_ | (~new_n18348_ & ~new_n18370_))));
  assign new_n18370_ = ~new_n18358_ & (new_n18343_ | (new_n18357_ & (~new_n18360_ | (~new_n18371_ & new_n18354_))));
  assign new_n18371_ = ~\all_features[837]  & \all_features[838]  & \all_features[839]  & (\all_features[836]  ? new_n18356_ : (new_n18345_ | ~new_n18356_));
  assign new_n18372_ = new_n18338_ ? (new_n18373_ ^ new_n18664_) : (~new_n18373_ ^ new_n18664_);
  assign new_n18373_ = new_n18374_ ^ new_n18570_;
  assign new_n18374_ = ~new_n18375_ & new_n18544_;
  assign new_n18375_ = new_n18376_ & (~new_n18477_ | new_n18455_);
  assign new_n18376_ = new_n18383_ & (~new_n9649_ | ~new_n18377_) & (~new_n18420_ | ~new_n18382_);
  assign new_n18377_ = new_n18378_ & new_n18380_;
  assign new_n18378_ = ~new_n10247_ & ~new_n18379_;
  assign new_n18379_ = ~new_n13733_ & ~new_n17001_ & ~new_n13709_;
  assign new_n18380_ = ~new_n15556_ & new_n18381_;
  assign new_n18381_ = ~new_n15577_ & new_n15918_;
  assign new_n18382_ = ~new_n18380_ & new_n18378_;
  assign new_n18383_ = (~new_n18394_ | ~new_n18384_) & (new_n18393_ | ~new_n18392_ | (~new_n18412_ & ~new_n18396_));
  assign new_n18384_ = new_n18385_ & new_n18391_;
  assign new_n18385_ = new_n18386_ & ~new_n16261_ & ~new_n16263_;
  assign new_n18386_ = ~new_n16235_ & (new_n16257_ | (~new_n16256_ & (new_n16254_ | new_n18387_)));
  assign new_n18387_ = ~new_n16252_ & (new_n16248_ | (~new_n16250_ & (new_n16258_ | (~new_n18388_ & ~new_n16260_))));
  assign new_n18388_ = ~new_n18389_ & \all_features[2775]  & (\all_features[2774]  | \all_features[2773]  | \all_features[2772] );
  assign new_n18389_ = \all_features[2775]  & ((~new_n18390_ & ~\all_features[2773]  & \all_features[2774] ) | (~new_n16242_ & (\all_features[2774]  | (~new_n16238_ & \all_features[2773] ))));
  assign new_n18390_ = (\all_features[2772]  & ~new_n16240_) | (~new_n16245_ & ~\all_features[2772]  & new_n16240_);
  assign new_n18391_ = ~new_n17258_ & new_n18379_;
  assign new_n18392_ = new_n17258_ & new_n18379_;
  assign new_n18393_ = ~new_n12834_ & ~new_n17256_ & ~new_n12825_;
  assign new_n18394_ = new_n10648_ & new_n18395_;
  assign new_n18395_ = ~new_n10677_ & ~new_n10679_;
  assign new_n18396_ = new_n18401_ & new_n18397_ & ~new_n18411_ & ~new_n18410_ & ~new_n18407_ & ~new_n18409_;
  assign new_n18397_ = ~new_n18398_ & (\all_features[2971]  | \all_features[2972]  | \all_features[2973]  | \all_features[2974]  | \all_features[2975] );
  assign new_n18398_ = ~\all_features[2973]  & new_n18399_ & ((~\all_features[2970]  & new_n18400_) | ~\all_features[2972]  | ~\all_features[2971] );
  assign new_n18399_ = ~\all_features[2974]  & ~\all_features[2975] ;
  assign new_n18400_ = ~\all_features[2968]  & ~\all_features[2969] ;
  assign new_n18401_ = ~new_n18402_ & ~new_n18406_;
  assign new_n18402_ = ~\all_features[2975]  & (~\all_features[2974]  | ~new_n18403_ | ~new_n18404_ | ~new_n18405_);
  assign new_n18403_ = \all_features[2970]  & \all_features[2971] ;
  assign new_n18404_ = \all_features[2968]  & \all_features[2969] ;
  assign new_n18405_ = \all_features[2972]  & \all_features[2973] ;
  assign new_n18406_ = ~\all_features[2975]  & (~\all_features[2974]  | (~\all_features[2972]  & ~\all_features[2973]  & ~new_n18403_));
  assign new_n18407_ = ~new_n18408_ & ~\all_features[2975] ;
  assign new_n18408_ = \all_features[2973]  & \all_features[2974]  & (\all_features[2972]  | (\all_features[2970]  & \all_features[2971]  & \all_features[2969] ));
  assign new_n18409_ = new_n18399_ & (~\all_features[2973]  | (~\all_features[2972]  & (~\all_features[2971]  | (~\all_features[2970]  & ~\all_features[2969] ))));
  assign new_n18410_ = ~\all_features[2975]  & (~\all_features[2974]  | (~\all_features[2973]  & (new_n18400_ | ~new_n18403_ | ~\all_features[2972] )));
  assign new_n18411_ = new_n18399_ & (~\all_features[2971]  | ~new_n18405_ | (~\all_features[2970]  & ~new_n18404_));
  assign new_n18412_ = new_n18397_ & new_n18419_ & (new_n18413_ | new_n18407_ | new_n18410_ | ~new_n18401_);
  assign new_n18413_ = new_n18418_ & new_n18417_ & new_n18414_ & new_n18416_;
  assign new_n18414_ = \all_features[2975]  & (\all_features[2974]  | (\all_features[2973]  & (\all_features[2972]  | ~new_n18415_ | ~new_n18400_)));
  assign new_n18415_ = ~\all_features[2970]  & ~\all_features[2971] ;
  assign new_n18416_ = \all_features[2975]  & (\all_features[2974]  | (new_n18405_ & (\all_features[2970]  | \all_features[2971]  | \all_features[2969] )));
  assign new_n18417_ = \all_features[2974]  & \all_features[2975]  & (\all_features[2972]  | \all_features[2973]  | new_n18404_ | ~new_n18415_);
  assign new_n18418_ = \all_features[2975]  & (\all_features[2973]  | \all_features[2974]  | \all_features[2972] );
  assign new_n18419_ = ~new_n18409_ & ~new_n18411_;
  assign new_n18420_ = new_n18421_ & ~new_n18447_ & ~new_n18451_;
  assign new_n18421_ = ~new_n18422_ & ~new_n18444_;
  assign new_n18422_ = new_n18439_ & ~new_n18443_ & ~new_n18423_ & ~new_n18442_;
  assign new_n18423_ = new_n18424_ & ~new_n18432_ & (~new_n18437_ | ~new_n18438_ | ~new_n18434_ | ~new_n18436_);
  assign new_n18424_ = ~new_n18429_ & ~new_n18425_ & ~new_n18427_;
  assign new_n18425_ = ~\all_features[4775]  & (~\all_features[4774]  | (~\all_features[4772]  & ~\all_features[4773]  & ~new_n18426_));
  assign new_n18426_ = \all_features[4770]  & \all_features[4771] ;
  assign new_n18427_ = ~new_n18428_ & ~\all_features[4775] ;
  assign new_n18428_ = \all_features[4773]  & \all_features[4774]  & (\all_features[4772]  | (\all_features[4770]  & \all_features[4771]  & \all_features[4769] ));
  assign new_n18429_ = ~\all_features[4775]  & (~\all_features[4774]  | ~new_n18430_ | ~new_n18431_ | ~new_n18426_);
  assign new_n18430_ = \all_features[4768]  & \all_features[4769] ;
  assign new_n18431_ = \all_features[4772]  & \all_features[4773] ;
  assign new_n18432_ = ~\all_features[4775]  & (~\all_features[4774]  | (~\all_features[4773]  & (new_n18433_ | ~new_n18426_ | ~\all_features[4772] )));
  assign new_n18433_ = ~\all_features[4768]  & ~\all_features[4769] ;
  assign new_n18434_ = \all_features[4775]  & (\all_features[4774]  | (\all_features[4773]  & (\all_features[4772]  | ~new_n18435_ | ~new_n18433_)));
  assign new_n18435_ = ~\all_features[4770]  & ~\all_features[4771] ;
  assign new_n18436_ = \all_features[4775]  & (\all_features[4774]  | (new_n18431_ & (\all_features[4770]  | \all_features[4771]  | \all_features[4769] )));
  assign new_n18437_ = \all_features[4774]  & \all_features[4775]  & (\all_features[4772]  | \all_features[4773]  | new_n18430_ | ~new_n18435_);
  assign new_n18438_ = \all_features[4775]  & (\all_features[4773]  | \all_features[4774]  | \all_features[4772] );
  assign new_n18439_ = ~new_n18440_ & (\all_features[4771]  | \all_features[4772]  | \all_features[4773]  | \all_features[4774]  | \all_features[4775] );
  assign new_n18440_ = new_n18441_ & (~\all_features[4771]  | ~new_n18431_ | (~\all_features[4770]  & ~new_n18430_));
  assign new_n18441_ = ~\all_features[4774]  & ~\all_features[4775] ;
  assign new_n18442_ = ~\all_features[4773]  & new_n18441_ & ((~\all_features[4770]  & new_n18433_) | ~\all_features[4772]  | ~\all_features[4771] );
  assign new_n18443_ = new_n18441_ & (~\all_features[4773]  | (~\all_features[4772]  & (~\all_features[4771]  | (~\all_features[4770]  & ~\all_features[4769] ))));
  assign new_n18444_ = new_n18424_ & new_n18446_ & ~new_n18432_ & new_n18445_;
  assign new_n18445_ = ~new_n18442_ & (\all_features[4771]  | \all_features[4772]  | \all_features[4773]  | \all_features[4774]  | \all_features[4775] );
  assign new_n18446_ = ~new_n18443_ & ~new_n18440_;
  assign new_n18447_ = ~new_n18448_ & (\all_features[4771]  | \all_features[4772]  | \all_features[4773]  | \all_features[4774]  | \all_features[4775] );
  assign new_n18448_ = ~new_n18442_ & (new_n18443_ | (~new_n18440_ & (new_n18425_ | (~new_n18449_ & ~new_n18432_))));
  assign new_n18449_ = ~new_n18427_ & (new_n18429_ | (new_n18438_ & (~new_n18434_ | (~new_n18450_ & new_n18436_))));
  assign new_n18450_ = ~\all_features[4773]  & \all_features[4774]  & \all_features[4775]  & (\all_features[4772]  ? new_n18435_ : (new_n18430_ | ~new_n18435_));
  assign new_n18451_ = new_n18445_ & (~new_n18446_ | (~new_n18452_ & ~new_n18425_ & ~new_n18432_));
  assign new_n18452_ = ~new_n18427_ & ~new_n18429_ & (~new_n18438_ | ~new_n18434_ | new_n18453_);
  assign new_n18453_ = new_n18436_ & new_n18437_ & (new_n18454_ | ~\all_features[4773]  | ~\all_features[4774]  | ~\all_features[4775] );
  assign new_n18454_ = ~\all_features[4771]  & ~\all_features[4772]  & (~\all_features[4770]  | new_n18433_);
  assign new_n18455_ = (new_n18420_ | ~new_n18382_) & (new_n18394_ | ~new_n18384_) & (new_n14953_ | ~new_n18456_);
  assign new_n18456_ = ~new_n18458_ & new_n18457_;
  assign new_n18457_ = ~new_n18379_ & new_n10247_;
  assign new_n18458_ = new_n18459_ & new_n18469_;
  assign new_n18459_ = ~new_n18460_ & ~new_n11704_;
  assign new_n18460_ = new_n11705_ & new_n18468_ & (new_n18461_ | new_n11716_ | new_n11719_ | ~new_n11710_);
  assign new_n18461_ = new_n18467_ & new_n18466_ & new_n18462_ & new_n18464_;
  assign new_n18462_ = \all_features[3543]  & (\all_features[3542]  | new_n18463_);
  assign new_n18463_ = \all_features[3541]  & (\all_features[3538]  | \all_features[3539]  | \all_features[3540]  | ~new_n11708_);
  assign new_n18464_ = \all_features[3543]  & ~new_n18465_ & \all_features[3542] ;
  assign new_n18465_ = ~\all_features[3541]  & ~\all_features[3540]  & ~\all_features[3539]  & ~new_n11713_ & ~\all_features[3538] ;
  assign new_n18466_ = \all_features[3543]  & (\all_features[3542]  | (new_n11714_ & (\all_features[3538]  | \all_features[3539]  | \all_features[3537] )));
  assign new_n18467_ = \all_features[3543]  & (\all_features[3541]  | \all_features[3542]  | \all_features[3540] );
  assign new_n18468_ = ~new_n11718_ & ~new_n11720_;
  assign new_n18469_ = ~new_n18470_ & (new_n11709_ | (~new_n18474_ & ~new_n11706_));
  assign new_n18470_ = new_n11705_ & (~new_n18468_ | (~new_n18471_ & ~new_n11719_ & ~new_n11715_));
  assign new_n18471_ = ~new_n11711_ & ~new_n11716_ & (~new_n18467_ | new_n18472_ | ~new_n18462_);
  assign new_n18472_ = ~new_n18465_ & new_n18466_ & \all_features[3542]  & \all_features[3543]  & (~\all_features[3541]  | new_n18473_);
  assign new_n18473_ = ~\all_features[3539]  & ~\all_features[3540]  & (~\all_features[3538]  | new_n11708_);
  assign new_n18474_ = ~new_n11718_ & (new_n11720_ | (~new_n11715_ & (new_n11719_ | (~new_n11716_ & ~new_n18475_))));
  assign new_n18475_ = ~new_n11711_ & (~new_n18467_ | (new_n18462_ & (~new_n18466_ | (~new_n18476_ & new_n18464_))));
  assign new_n18476_ = \all_features[3542]  & \all_features[3543]  & (\all_features[3541]  | (\all_features[3540]  & (\all_features[3539]  | \all_features[3538] )));
  assign new_n18477_ = (new_n18511_ | ~new_n18479_) & (~new_n18478_ | ~new_n18480_);
  assign new_n18478_ = ~new_n18385_ & new_n18391_;
  assign new_n18479_ = new_n18392_ & new_n18393_;
  assign new_n18480_ = new_n18510_ & (new_n18507_ | new_n18481_);
  assign new_n18481_ = new_n18501_ & (~new_n18497_ | (new_n18493_ & (new_n18482_ | new_n18504_ | new_n18506_)));
  assign new_n18482_ = new_n18491_ & new_n18492_ & (~new_n18488_ | ~new_n18486_ | new_n18483_);
  assign new_n18483_ = \all_features[5103]  & \all_features[5102]  & ~new_n18484_ & \all_features[5101] ;
  assign new_n18484_ = ~\all_features[5099]  & ~\all_features[5100]  & (~\all_features[5098]  | new_n18485_);
  assign new_n18485_ = ~\all_features[5096]  & ~\all_features[5097] ;
  assign new_n18486_ = \all_features[5103]  & (\all_features[5102]  | (new_n18487_ & (\all_features[5098]  | \all_features[5099]  | \all_features[5097] )));
  assign new_n18487_ = \all_features[5100]  & \all_features[5101] ;
  assign new_n18488_ = \all_features[5102]  & \all_features[5103]  & (\all_features[5100]  | \all_features[5101]  | new_n18489_ | ~new_n18490_);
  assign new_n18489_ = \all_features[5096]  & \all_features[5097] ;
  assign new_n18490_ = ~\all_features[5098]  & ~\all_features[5099] ;
  assign new_n18491_ = \all_features[5103]  & (\all_features[5102]  | (\all_features[5101]  & (\all_features[5100]  | ~new_n18490_ | ~new_n18485_)));
  assign new_n18492_ = \all_features[5103]  & (\all_features[5101]  | \all_features[5102]  | \all_features[5100] );
  assign new_n18493_ = ~new_n18494_ & ~new_n18496_;
  assign new_n18494_ = ~\all_features[5103]  & (~\all_features[5102]  | (~\all_features[5100]  & ~\all_features[5101]  & ~new_n18495_));
  assign new_n18495_ = \all_features[5098]  & \all_features[5099] ;
  assign new_n18496_ = ~\all_features[5103]  & (~\all_features[5102]  | (~\all_features[5101]  & (new_n18485_ | ~\all_features[5100]  | ~new_n18495_)));
  assign new_n18497_ = ~new_n18498_ & ~new_n18500_;
  assign new_n18498_ = new_n18499_ & (~\all_features[5101]  | (~\all_features[5100]  & (~\all_features[5099]  | (~\all_features[5098]  & ~\all_features[5097] ))));
  assign new_n18499_ = ~\all_features[5102]  & ~\all_features[5103] ;
  assign new_n18500_ = new_n18499_ & (~\all_features[5099]  | ~new_n18487_ | (~\all_features[5098]  & ~new_n18489_));
  assign new_n18501_ = ~new_n18502_ & ~new_n18503_;
  assign new_n18502_ = ~\all_features[5101]  & new_n18499_ & ((~\all_features[5098]  & new_n18485_) | ~\all_features[5100]  | ~\all_features[5099] );
  assign new_n18503_ = ~\all_features[5103]  & ~\all_features[5102]  & ~\all_features[5101]  & ~\all_features[5099]  & ~\all_features[5100] ;
  assign new_n18504_ = ~new_n18505_ & ~\all_features[5103] ;
  assign new_n18505_ = \all_features[5101]  & \all_features[5102]  & (\all_features[5100]  | (\all_features[5098]  & \all_features[5099]  & \all_features[5097] ));
  assign new_n18506_ = ~\all_features[5103]  & (~\all_features[5102]  | ~new_n18495_ | ~new_n18489_ | ~new_n18487_);
  assign new_n18507_ = new_n18501_ & ~new_n18508_ & new_n18497_;
  assign new_n18508_ = new_n18509_ & (~new_n18491_ | ~new_n18492_ | ~new_n18486_ | ~new_n18488_);
  assign new_n18509_ = ~new_n18506_ & ~new_n18504_ & ~new_n18494_ & ~new_n18496_;
  assign new_n18510_ = new_n18497_ & new_n18493_ & ~new_n18503_ & ~new_n18506_ & ~new_n18504_ & ~new_n18502_;
  assign new_n18511_ = ~new_n18512_ & new_n18539_;
  assign new_n18512_ = ~new_n18538_ & (~new_n18531_ | (~new_n18536_ & (new_n18529_ | new_n18537_ | ~new_n18513_)));
  assign new_n18513_ = ~new_n18525_ & ~new_n18523_ & ((~new_n18520_ & new_n18514_) | ~new_n18528_ | ~new_n18527_);
  assign new_n18514_ = \all_features[4519]  & \all_features[4518]  & ~new_n18517_ & new_n18515_;
  assign new_n18515_ = \all_features[4519]  & (\all_features[4518]  | (new_n18516_ & (\all_features[4514]  | \all_features[4515]  | \all_features[4513] )));
  assign new_n18516_ = \all_features[4516]  & \all_features[4517] ;
  assign new_n18517_ = new_n18519_ & ~\all_features[4517]  & ~new_n18518_ & ~\all_features[4516] ;
  assign new_n18518_ = \all_features[4512]  & \all_features[4513] ;
  assign new_n18519_ = ~\all_features[4514]  & ~\all_features[4515] ;
  assign new_n18520_ = \all_features[4519]  & \all_features[4518]  & ~new_n18521_ & \all_features[4517] ;
  assign new_n18521_ = ~\all_features[4515]  & ~\all_features[4516]  & (~\all_features[4514]  | new_n18522_);
  assign new_n18522_ = ~\all_features[4512]  & ~\all_features[4513] ;
  assign new_n18523_ = ~new_n18524_ & ~\all_features[4519] ;
  assign new_n18524_ = \all_features[4517]  & \all_features[4518]  & (\all_features[4516]  | (\all_features[4514]  & \all_features[4515]  & \all_features[4513] ));
  assign new_n18525_ = ~\all_features[4519]  & (~\all_features[4518]  | ~new_n18526_ | ~new_n18518_ | ~new_n18516_);
  assign new_n18526_ = \all_features[4514]  & \all_features[4515] ;
  assign new_n18527_ = \all_features[4519]  & (\all_features[4518]  | (\all_features[4517]  & (\all_features[4516]  | ~new_n18519_ | ~new_n18522_)));
  assign new_n18528_ = \all_features[4519]  & (\all_features[4517]  | \all_features[4518]  | \all_features[4516] );
  assign new_n18529_ = ~new_n18523_ & (new_n18525_ | (new_n18528_ & (~new_n18527_ | (~new_n18530_ & new_n18515_))));
  assign new_n18530_ = ~\all_features[4517]  & \all_features[4518]  & \all_features[4519]  & (\all_features[4516]  ? new_n18519_ : (new_n18518_ | ~new_n18519_));
  assign new_n18531_ = ~new_n18535_ & ~new_n18532_ & ~new_n18534_;
  assign new_n18532_ = new_n18533_ & (~\all_features[4517]  | (~\all_features[4516]  & (~\all_features[4515]  | (~\all_features[4514]  & ~\all_features[4513] ))));
  assign new_n18533_ = ~\all_features[4518]  & ~\all_features[4519] ;
  assign new_n18534_ = ~\all_features[4517]  & new_n18533_ & ((~\all_features[4514]  & new_n18522_) | ~\all_features[4516]  | ~\all_features[4515] );
  assign new_n18535_ = new_n18533_ & (~\all_features[4515]  | ~new_n18516_ | (~\all_features[4514]  & ~new_n18518_));
  assign new_n18536_ = ~\all_features[4519]  & (~\all_features[4518]  | (~\all_features[4516]  & ~\all_features[4517]  & ~new_n18526_));
  assign new_n18537_ = ~\all_features[4519]  & (~\all_features[4518]  | (~\all_features[4517]  & (new_n18522_ | ~\all_features[4516]  | ~new_n18526_)));
  assign new_n18538_ = ~\all_features[4519]  & ~\all_features[4518]  & ~\all_features[4517]  & ~\all_features[4515]  & ~\all_features[4516] ;
  assign new_n18539_ = new_n18532_ | ~new_n18542_ | ((new_n18523_ | ~new_n18543_) & (new_n18540_ | new_n18535_));
  assign new_n18540_ = new_n18541_ & (~new_n18514_ | ~new_n18527_ | ~new_n18528_);
  assign new_n18541_ = ~new_n18525_ & ~new_n18523_ & ~new_n18536_ & ~new_n18537_;
  assign new_n18542_ = ~new_n18534_ & ~new_n18538_;
  assign new_n18543_ = ~new_n18535_ & ~new_n18525_ & ~new_n18536_ & ~new_n18537_;
  assign new_n18544_ = new_n18545_ & new_n18546_ & (~new_n18511_ | ~new_n18479_);
  assign new_n18545_ = (~new_n14953_ | ~new_n18456_) & (new_n9649_ | ~new_n18377_);
  assign new_n18546_ = (~new_n18478_ | new_n18480_) & (~new_n18458_ | ~new_n18457_ | ~new_n18547_);
  assign new_n18547_ = new_n18548_ & new_n18568_;
  assign new_n18548_ = new_n18563_ & ~new_n18567_ & ~new_n18549_ & ~new_n18565_;
  assign new_n18549_ = ~new_n18561_ & new_n18550_ & (~new_n18559_ | ~new_n18558_);
  assign new_n18550_ = ~new_n18555_ & ~new_n18551_ & ~new_n18553_;
  assign new_n18551_ = ~new_n18552_ & ~\all_features[2959] ;
  assign new_n18552_ = \all_features[2957]  & \all_features[2958]  & (\all_features[2956]  | (\all_features[2954]  & \all_features[2955]  & \all_features[2953] ));
  assign new_n18553_ = ~\all_features[2959]  & (~\all_features[2958]  | (~\all_features[2956]  & ~\all_features[2957]  & ~new_n18554_));
  assign new_n18554_ = \all_features[2954]  & \all_features[2955] ;
  assign new_n18555_ = ~\all_features[2959]  & (~\all_features[2958]  | ~new_n18556_ | ~new_n18557_ | ~new_n18554_);
  assign new_n18556_ = \all_features[2956]  & \all_features[2957] ;
  assign new_n18557_ = \all_features[2952]  & \all_features[2953] ;
  assign new_n18558_ = \all_features[2959]  & (\all_features[2958]  | (new_n18556_ & (\all_features[2954]  | \all_features[2955]  | \all_features[2953] )));
  assign new_n18559_ = new_n18560_ & (new_n18557_ | \all_features[2954]  | \all_features[2955]  | \all_features[2956]  | \all_features[2957] );
  assign new_n18560_ = \all_features[2958]  & \all_features[2959] ;
  assign new_n18561_ = ~\all_features[2959]  & (~\all_features[2958]  | (~\all_features[2957]  & (new_n18562_ | ~\all_features[2956]  | ~new_n18554_)));
  assign new_n18562_ = ~\all_features[2952]  & ~\all_features[2953] ;
  assign new_n18563_ = \all_features[2957]  | \all_features[2958]  | \all_features[2959]  | (\all_features[2956]  & \all_features[2955]  & ~new_n18564_);
  assign new_n18564_ = ~\all_features[2954]  & new_n18562_;
  assign new_n18565_ = ~\all_features[2959]  & ~new_n18566_ & ~\all_features[2958] ;
  assign new_n18566_ = \all_features[2957]  & (\all_features[2956]  | (\all_features[2955]  & (\all_features[2954]  | \all_features[2953] )));
  assign new_n18567_ = ~\all_features[2958]  & ~\all_features[2959]  & (~\all_features[2955]  | ~new_n18556_ | (~\all_features[2954]  & ~new_n18557_));
  assign new_n18568_ = new_n18550_ & new_n18569_ & ~new_n18561_ & new_n18563_;
  assign new_n18569_ = ~new_n18565_ & ~new_n18567_;
  assign new_n18570_ = ~new_n18571_ & new_n18591_;
  assign new_n18571_ = new_n18572_ & (~new_n18574_ | ~new_n18590_ | new_n18588_ | new_n18576_);
  assign new_n18572_ = ~new_n18573_ & (new_n18574_ | new_n18582_ | new_n17927_ | ~new_n18580_);
  assign new_n18573_ = ~new_n18578_ & new_n18576_ & new_n18574_ & (new_n6662_ | (new_n16999_ & new_n6640_));
  assign new_n18574_ = new_n10839_ & new_n18575_;
  assign new_n18575_ = ~new_n10871_ & ~new_n10868_;
  assign new_n18576_ = new_n11061_ & new_n18577_;
  assign new_n18577_ = ~new_n6569_ & ~new_n6591_;
  assign new_n18578_ = new_n9346_ & new_n18579_;
  assign new_n18579_ = ~new_n9376_ & ~new_n9379_;
  assign new_n18580_ = ~new_n16316_ & new_n18581_;
  assign new_n18581_ = ~new_n16305_ & ~new_n16313_;
  assign new_n18582_ = ~new_n10127_ & ~new_n18583_ & ~new_n10100_ & ~new_n10125_;
  assign new_n18583_ = ~new_n10102_ & (new_n10105_ | (~new_n10117_ & (new_n10116_ | (~new_n18584_ & ~new_n10119_))));
  assign new_n18584_ = ~new_n10121_ & (new_n10123_ | (~new_n10122_ & (~new_n18587_ | new_n18585_)));
  assign new_n18585_ = \all_features[1031]  & ((~new_n18586_ & ~\all_features[1029]  & \all_features[1030] ) | (~new_n10111_ & (\all_features[1030]  | (~new_n10109_ & \all_features[1029] ))));
  assign new_n18586_ = (~\all_features[1026]  & ~\all_features[1027]  & ~\all_features[1028]  & (~\all_features[1025]  | ~\all_features[1024] )) | (\all_features[1028]  & (\all_features[1026]  | \all_features[1027] ));
  assign new_n18587_ = \all_features[1031]  & (\all_features[1029]  | \all_features[1030]  | \all_features[1028] );
  assign new_n18588_ = new_n18589_ & ~new_n7767_ & ~new_n7769_;
  assign new_n18589_ = ~new_n7738_ & ~new_n7760_;
  assign new_n18590_ = ~new_n7835_ & new_n12756_;
  assign new_n18591_ = new_n18595_ & (~new_n18574_ | (new_n18592_ & (new_n18576_ | ~new_n18588_ | ~new_n18590_)));
  assign new_n18592_ = (~new_n18593_ | ~new_n18576_) & (new_n18594_ | new_n18590_ | new_n18576_);
  assign new_n18593_ = new_n7517_ & new_n18578_ & ~new_n7547_ & ~new_n7550_;
  assign new_n18594_ = ~new_n8915_ & new_n8923_;
  assign new_n18595_ = new_n18574_ | (new_n18582_ ? (new_n12802_ ? new_n18632_ : new_n18634_) : new_n18596_);
  assign new_n18596_ = (new_n18580_ | new_n17927_) & (~new_n18597_ | ~new_n18626_ | ~new_n17927_);
  assign new_n18597_ = ~new_n18598_ & ~new_n18619_;
  assign new_n18598_ = ~new_n18599_ & (\all_features[1723]  | \all_features[1724]  | \all_features[1725]  | \all_features[1726]  | \all_features[1727] );
  assign new_n18599_ = ~new_n18613_ & (new_n18615_ | (~new_n18616_ & (new_n18617_ | (~new_n18600_ & ~new_n18618_))));
  assign new_n18600_ = ~new_n18601_ & (new_n18603_ | (new_n18612_ & (~new_n18607_ | (~new_n18611_ & new_n18610_))));
  assign new_n18601_ = ~new_n18602_ & ~\all_features[1727] ;
  assign new_n18602_ = \all_features[1725]  & \all_features[1726]  & (\all_features[1724]  | (\all_features[1722]  & \all_features[1723]  & \all_features[1721] ));
  assign new_n18603_ = ~\all_features[1727]  & (~\all_features[1726]  | ~new_n18604_ | ~new_n18605_ | ~new_n18606_);
  assign new_n18604_ = \all_features[1720]  & \all_features[1721] ;
  assign new_n18605_ = \all_features[1724]  & \all_features[1725] ;
  assign new_n18606_ = \all_features[1722]  & \all_features[1723] ;
  assign new_n18607_ = \all_features[1727]  & (\all_features[1726]  | (\all_features[1725]  & (\all_features[1724]  | ~new_n18609_ | ~new_n18608_)));
  assign new_n18608_ = ~\all_features[1720]  & ~\all_features[1721] ;
  assign new_n18609_ = ~\all_features[1722]  & ~\all_features[1723] ;
  assign new_n18610_ = \all_features[1727]  & (\all_features[1726]  | (new_n18605_ & (\all_features[1722]  | \all_features[1723]  | \all_features[1721] )));
  assign new_n18611_ = ~\all_features[1725]  & \all_features[1726]  & \all_features[1727]  & (\all_features[1724]  ? new_n18609_ : (new_n18604_ | ~new_n18609_));
  assign new_n18612_ = \all_features[1727]  & (\all_features[1725]  | \all_features[1726]  | \all_features[1724] );
  assign new_n18613_ = ~\all_features[1725]  & new_n18614_ & ((~\all_features[1722]  & new_n18608_) | ~\all_features[1724]  | ~\all_features[1723] );
  assign new_n18614_ = ~\all_features[1726]  & ~\all_features[1727] ;
  assign new_n18615_ = new_n18614_ & (~\all_features[1725]  | (~\all_features[1724]  & (~\all_features[1723]  | (~\all_features[1722]  & ~\all_features[1721] ))));
  assign new_n18616_ = new_n18614_ & (~\all_features[1723]  | ~new_n18605_ | (~\all_features[1722]  & ~new_n18604_));
  assign new_n18617_ = ~\all_features[1727]  & (~\all_features[1726]  | (~\all_features[1724]  & ~\all_features[1725]  & ~new_n18606_));
  assign new_n18618_ = ~\all_features[1727]  & (~\all_features[1726]  | (~\all_features[1725]  & (new_n18608_ | ~new_n18606_ | ~\all_features[1724] )));
  assign new_n18619_ = new_n18624_ & (~new_n18625_ | (~new_n18620_ & ~new_n18617_ & ~new_n18618_));
  assign new_n18620_ = ~new_n18601_ & ~new_n18603_ & (~new_n18612_ | ~new_n18607_ | new_n18621_);
  assign new_n18621_ = new_n18610_ & new_n18622_ & (new_n18623_ | ~\all_features[1725]  | ~\all_features[1726]  | ~\all_features[1727] );
  assign new_n18622_ = \all_features[1726]  & \all_features[1727]  & (\all_features[1724]  | \all_features[1725]  | new_n18604_ | ~new_n18609_);
  assign new_n18623_ = ~\all_features[1723]  & ~\all_features[1724]  & (~\all_features[1722]  | new_n18608_);
  assign new_n18624_ = ~new_n18613_ & (\all_features[1723]  | \all_features[1724]  | \all_features[1725]  | \all_features[1726]  | \all_features[1727] );
  assign new_n18625_ = ~new_n18615_ & ~new_n18616_;
  assign new_n18626_ = ~new_n18627_ & ~new_n18631_;
  assign new_n18627_ = new_n18624_ & ~new_n18616_ & ~new_n18628_ & ~new_n18615_;
  assign new_n18628_ = ~new_n18618_ & ~new_n18603_ & new_n18630_ & (~new_n18607_ | ~new_n18629_);
  assign new_n18629_ = new_n18612_ & new_n18610_ & new_n18622_;
  assign new_n18630_ = ~new_n18617_ & ~new_n18601_;
  assign new_n18631_ = new_n18625_ & new_n18624_ & new_n18630_ & ~new_n18618_ & ~new_n18603_;
  assign new_n18632_ = new_n18633_ & new_n8097_;
  assign new_n18633_ = new_n8083_ & new_n8094_;
  assign new_n18634_ = new_n18662_ & new_n18661_ & (new_n18660_ | (~new_n18635_ & ~new_n18663_));
  assign new_n18635_ = new_n18653_ & (new_n18659_ | (~new_n18658_ & new_n18648_ & (new_n18651_ | new_n18636_)));
  assign new_n18636_ = ~new_n18640_ & (~new_n18646_ | (new_n18637_ & (~new_n18643_ | (~new_n18647_ & new_n18644_))));
  assign new_n18637_ = \all_features[4679]  & (\all_features[4678]  | new_n18638_);
  assign new_n18638_ = \all_features[4677]  & (\all_features[4674]  | \all_features[4675]  | \all_features[4676]  | ~new_n18639_);
  assign new_n18639_ = ~\all_features[4672]  & ~\all_features[4673] ;
  assign new_n18640_ = ~\all_features[4679]  & (~new_n18642_ | ~\all_features[4672]  | ~\all_features[4673]  | ~\all_features[4678]  | ~new_n18641_);
  assign new_n18641_ = \all_features[4674]  & \all_features[4675] ;
  assign new_n18642_ = \all_features[4676]  & \all_features[4677] ;
  assign new_n18643_ = \all_features[4679]  & (\all_features[4678]  | (new_n18642_ & (\all_features[4674]  | \all_features[4675]  | \all_features[4673] )));
  assign new_n18644_ = \all_features[4679]  & ~new_n18645_ & \all_features[4678] ;
  assign new_n18645_ = ~\all_features[4674]  & ~\all_features[4675]  & ~\all_features[4676]  & ~\all_features[4677]  & (~\all_features[4673]  | ~\all_features[4672] );
  assign new_n18646_ = \all_features[4679]  & (\all_features[4677]  | \all_features[4678]  | \all_features[4676] );
  assign new_n18647_ = \all_features[4678]  & \all_features[4679]  & (\all_features[4677]  | (\all_features[4676]  & (\all_features[4675]  | \all_features[4674] )));
  assign new_n18648_ = ~new_n18640_ & ~new_n18651_ & (~new_n18646_ | new_n18649_ | ~new_n18637_);
  assign new_n18649_ = ~new_n18645_ & new_n18643_ & \all_features[4678]  & \all_features[4679]  & (~\all_features[4677]  | new_n18650_);
  assign new_n18650_ = ~\all_features[4675]  & ~\all_features[4676]  & (~\all_features[4674]  | new_n18639_);
  assign new_n18651_ = ~new_n18652_ & ~\all_features[4679] ;
  assign new_n18652_ = \all_features[4677]  & \all_features[4678]  & (\all_features[4676]  | (\all_features[4674]  & \all_features[4675]  & \all_features[4673] ));
  assign new_n18653_ = ~new_n18657_ & ~new_n18654_ & ~new_n18656_;
  assign new_n18654_ = new_n18655_ & (~\all_features[4677]  | (~\all_features[4676]  & (~\all_features[4675]  | (~\all_features[4674]  & ~\all_features[4673] ))));
  assign new_n18655_ = ~\all_features[4678]  & ~\all_features[4679] ;
  assign new_n18656_ = new_n18655_ & (~new_n18642_ | ~\all_features[4675]  | (~\all_features[4674]  & (~\all_features[4672]  | ~\all_features[4673] )));
  assign new_n18657_ = ~\all_features[4677]  & new_n18655_ & ((~\all_features[4674]  & new_n18639_) | ~\all_features[4676]  | ~\all_features[4675] );
  assign new_n18658_ = ~\all_features[4679]  & (~\all_features[4678]  | (~\all_features[4677]  & (new_n18639_ | ~\all_features[4676]  | ~new_n18641_)));
  assign new_n18659_ = ~\all_features[4679]  & (~\all_features[4678]  | (~\all_features[4676]  & ~\all_features[4677]  & ~new_n18641_));
  assign new_n18660_ = new_n18646_ & new_n18644_ & new_n18637_ & new_n18643_;
  assign new_n18661_ = ~new_n18640_ & ~new_n18659_ & ~new_n18658_ & ~new_n18651_;
  assign new_n18662_ = ~new_n18663_ & ~new_n18657_ & ~new_n18654_ & ~new_n18656_;
  assign new_n18663_ = ~\all_features[4679]  & ~\all_features[4678]  & ~\all_features[4677]  & ~\all_features[4675]  & ~\all_features[4676] ;
  assign new_n18664_ = new_n18665_ ? (new_n18790_ ^ new_n18852_) : (~new_n18790_ ^ new_n18852_);
  assign new_n18665_ = ~new_n18787_ & new_n18666_;
  assign new_n18666_ = new_n18667_ & (new_n8739_ | (new_n18753_ & (new_n12870_ | new_n14725_ | ~new_n18786_)));
  assign new_n18667_ = new_n18668_ & (~new_n18749_ | (new_n18750_ & new_n18751_) | (new_n12398_ & ~new_n18751_));
  assign new_n18668_ = new_n18706_ | ~new_n8739_ | (new_n18739_ ? new_n18669_ : (~new_n18744_ & new_n18740_));
  assign new_n18669_ = new_n18670_ & new_n18701_;
  assign new_n18670_ = ~new_n18671_ & ~new_n18691_;
  assign new_n18671_ = (new_n18672_ | (new_n18690_ & (~\all_features[5307]  | ~\all_features[5308]  | (~\all_features[5306]  & new_n18676_)))) & (~new_n18690_ | \all_features[5307]  | \all_features[5308] );
  assign new_n18672_ = ~new_n18683_ & (new_n18685_ | (~new_n18686_ & (new_n18687_ | (~new_n18673_ & ~new_n18688_))));
  assign new_n18673_ = ~new_n18681_ & (~\all_features[5311]  | new_n18674_ | (~\all_features[5308]  & ~\all_features[5309]  & ~\all_features[5310] ));
  assign new_n18674_ = \all_features[5311]  & ((~new_n18677_ & ~\all_features[5309]  & \all_features[5310] ) | (~new_n18679_ & (\all_features[5310]  | (~new_n18675_ & \all_features[5309] ))));
  assign new_n18675_ = new_n18676_ & ~\all_features[5308]  & ~\all_features[5306]  & ~\all_features[5307] ;
  assign new_n18676_ = ~\all_features[5304]  & ~\all_features[5305] ;
  assign new_n18677_ = (\all_features[5308]  & (\all_features[5306]  | \all_features[5307] )) | (~new_n18678_ & ~\all_features[5306]  & ~\all_features[5307]  & ~\all_features[5308] );
  assign new_n18678_ = \all_features[5304]  & \all_features[5305] ;
  assign new_n18679_ = \all_features[5311]  & (\all_features[5310]  | (new_n18680_ & (\all_features[5306]  | \all_features[5307]  | \all_features[5305] )));
  assign new_n18680_ = \all_features[5308]  & \all_features[5309] ;
  assign new_n18681_ = ~\all_features[5311]  & (~\all_features[5310]  | ~new_n18678_ | ~new_n18680_ | ~new_n18682_);
  assign new_n18682_ = \all_features[5306]  & \all_features[5307] ;
  assign new_n18683_ = ~\all_features[5311]  & ~new_n18684_ & ~\all_features[5310] ;
  assign new_n18684_ = \all_features[5309]  & (\all_features[5308]  | (\all_features[5307]  & (\all_features[5306]  | \all_features[5305] )));
  assign new_n18685_ = ~\all_features[5310]  & ~\all_features[5311]  & (~\all_features[5307]  | ~new_n18680_ | (~\all_features[5306]  & ~new_n18678_));
  assign new_n18686_ = ~\all_features[5311]  & (~\all_features[5310]  | (~\all_features[5308]  & ~\all_features[5309]  & ~new_n18682_));
  assign new_n18687_ = ~\all_features[5311]  & (~\all_features[5310]  | (~\all_features[5309]  & (new_n18676_ | ~new_n18682_ | ~\all_features[5308] )));
  assign new_n18688_ = ~new_n18689_ & ~\all_features[5311] ;
  assign new_n18689_ = \all_features[5309]  & \all_features[5310]  & (\all_features[5308]  | (\all_features[5306]  & \all_features[5307]  & \all_features[5305] ));
  assign new_n18690_ = ~\all_features[5311]  & ~\all_features[5309]  & ~\all_features[5310] ;
  assign new_n18691_ = new_n18700_ & (~new_n18697_ | (new_n18698_ & (~new_n18699_ | new_n18692_)));
  assign new_n18692_ = new_n18693_ & (~new_n18694_ | (~new_n18696_ & \all_features[5309]  & \all_features[5310]  & \all_features[5311] ));
  assign new_n18693_ = \all_features[5311]  & (\all_features[5310]  | (~new_n18675_ & \all_features[5309] ));
  assign new_n18694_ = \all_features[5311]  & \all_features[5310]  & ~new_n18695_ & new_n18679_;
  assign new_n18695_ = ~\all_features[5309]  & ~\all_features[5308]  & ~\all_features[5307]  & ~new_n18678_ & ~\all_features[5306] ;
  assign new_n18696_ = ~\all_features[5307]  & ~\all_features[5308]  & (~\all_features[5306]  | new_n18676_);
  assign new_n18697_ = ~new_n18683_ & ~new_n18685_;
  assign new_n18698_ = ~new_n18686_ & ~new_n18687_;
  assign new_n18699_ = ~new_n18688_ & ~new_n18681_;
  assign new_n18700_ = ~new_n18690_ | (\all_features[5307]  & \all_features[5308]  & (\all_features[5306]  | ~new_n18676_));
  assign new_n18701_ = ~new_n18702_ & ~new_n18705_;
  assign new_n18702_ = new_n18703_ & (new_n18687_ | new_n18688_ | ~new_n18704_ | (new_n18694_ & new_n18693_));
  assign new_n18703_ = new_n18697_ & new_n18700_;
  assign new_n18704_ = ~new_n18686_ & ~new_n18681_;
  assign new_n18705_ = new_n18699_ & new_n18703_ & new_n18698_;
  assign new_n18706_ = ~new_n18707_ & new_n18734_;
  assign new_n18707_ = ~new_n18733_ & (~new_n18726_ | (~new_n18731_ & (new_n18724_ | new_n18732_ | ~new_n18708_)));
  assign new_n18708_ = ~new_n18720_ & ~new_n18718_ & ((~new_n18715_ & new_n18709_) | ~new_n18723_ | ~new_n18722_);
  assign new_n18709_ = \all_features[5111]  & \all_features[5110]  & ~new_n18712_ & new_n18710_;
  assign new_n18710_ = \all_features[5111]  & (\all_features[5110]  | (new_n18711_ & (\all_features[5106]  | \all_features[5107]  | \all_features[5105] )));
  assign new_n18711_ = \all_features[5108]  & \all_features[5109] ;
  assign new_n18712_ = new_n18714_ & ~\all_features[5109]  & ~new_n18713_ & ~\all_features[5108] ;
  assign new_n18713_ = \all_features[5104]  & \all_features[5105] ;
  assign new_n18714_ = ~\all_features[5106]  & ~\all_features[5107] ;
  assign new_n18715_ = \all_features[5111]  & \all_features[5110]  & ~new_n18716_ & \all_features[5109] ;
  assign new_n18716_ = ~\all_features[5107]  & ~\all_features[5108]  & (~\all_features[5106]  | new_n18717_);
  assign new_n18717_ = ~\all_features[5104]  & ~\all_features[5105] ;
  assign new_n18718_ = ~new_n18719_ & ~\all_features[5111] ;
  assign new_n18719_ = \all_features[5109]  & \all_features[5110]  & (\all_features[5108]  | (\all_features[5106]  & \all_features[5107]  & \all_features[5105] ));
  assign new_n18720_ = ~\all_features[5111]  & (~\all_features[5110]  | ~new_n18721_ | ~new_n18713_ | ~new_n18711_);
  assign new_n18721_ = \all_features[5106]  & \all_features[5107] ;
  assign new_n18722_ = \all_features[5111]  & (\all_features[5110]  | (\all_features[5109]  & (\all_features[5108]  | ~new_n18714_ | ~new_n18717_)));
  assign new_n18723_ = \all_features[5111]  & (\all_features[5109]  | \all_features[5110]  | \all_features[5108] );
  assign new_n18724_ = ~new_n18718_ & (new_n18720_ | (new_n18723_ & (~new_n18722_ | (~new_n18725_ & new_n18710_))));
  assign new_n18725_ = ~\all_features[5109]  & \all_features[5110]  & \all_features[5111]  & (\all_features[5108]  ? new_n18714_ : (new_n18713_ | ~new_n18714_));
  assign new_n18726_ = ~new_n18730_ & ~new_n18727_ & ~new_n18729_;
  assign new_n18727_ = new_n18728_ & (~\all_features[5109]  | (~\all_features[5108]  & (~\all_features[5107]  | (~\all_features[5106]  & ~\all_features[5105] ))));
  assign new_n18728_ = ~\all_features[5110]  & ~\all_features[5111] ;
  assign new_n18729_ = ~\all_features[5109]  & new_n18728_ & ((~\all_features[5106]  & new_n18717_) | ~\all_features[5108]  | ~\all_features[5107] );
  assign new_n18730_ = new_n18728_ & (~\all_features[5107]  | ~new_n18711_ | (~\all_features[5106]  & ~new_n18713_));
  assign new_n18731_ = ~\all_features[5111]  & (~\all_features[5110]  | (~\all_features[5108]  & ~\all_features[5109]  & ~new_n18721_));
  assign new_n18732_ = ~\all_features[5111]  & (~\all_features[5110]  | (~\all_features[5109]  & (new_n18717_ | ~\all_features[5108]  | ~new_n18721_)));
  assign new_n18733_ = ~\all_features[5111]  & ~\all_features[5110]  & ~\all_features[5109]  & ~\all_features[5107]  & ~\all_features[5108] ;
  assign new_n18734_ = new_n18727_ | ~new_n18737_ | ((new_n18718_ | ~new_n18738_) & (new_n18735_ | new_n18730_));
  assign new_n18735_ = new_n18736_ & (~new_n18709_ | ~new_n18722_ | ~new_n18723_);
  assign new_n18736_ = ~new_n18720_ & ~new_n18718_ & ~new_n18731_ & ~new_n18732_;
  assign new_n18737_ = ~new_n18729_ & ~new_n18733_;
  assign new_n18738_ = ~new_n18730_ & ~new_n18720_ & ~new_n18731_ & ~new_n18732_;
  assign new_n18739_ = new_n17619_ & new_n17621_;
  assign new_n18740_ = ~new_n17284_ & ~new_n17262_ & (~new_n17278_ | (~new_n18741_ & ~new_n17282_ & ~new_n17283_));
  assign new_n18741_ = ~new_n17272_ & ~new_n17277_ & (new_n17276_ | new_n17274_ | new_n18742_);
  assign new_n18742_ = new_n17264_ & (~new_n17267_ | (~new_n18743_ & \all_features[3765]  & \all_features[3766]  & \all_features[3767] ));
  assign new_n18743_ = ~\all_features[3763]  & ~\all_features[3764]  & (~\all_features[3762]  | new_n17266_);
  assign new_n18744_ = ~new_n17281_ & (new_n17279_ | (~new_n17282_ & (new_n17283_ | (~new_n18745_ & ~new_n17277_))));
  assign new_n18745_ = ~new_n17272_ & (new_n17274_ | (~new_n17276_ & (~new_n18748_ | new_n18746_)));
  assign new_n18746_ = \all_features[3767]  & ((~new_n18747_ & ~\all_features[3765]  & \all_features[3766] ) | (~new_n17268_ & (\all_features[3766]  | (~new_n17265_ & \all_features[3765] ))));
  assign new_n18747_ = (\all_features[3764]  & (\all_features[3762]  | \all_features[3763] )) | (~new_n17271_ & ~\all_features[3762]  & ~\all_features[3763]  & ~\all_features[3764] );
  assign new_n18748_ = \all_features[3767]  & (\all_features[3765]  | \all_features[3766]  | \all_features[3764] );
  assign new_n18749_ = new_n18706_ & new_n8739_;
  assign new_n18750_ = new_n9583_ & ~new_n10527_ & ~new_n10531_;
  assign new_n18751_ = ~new_n11887_ & new_n18752_;
  assign new_n18752_ = ~new_n11861_ & ~new_n11884_;
  assign new_n18753_ = (new_n14469_ | new_n18755_ | ~new_n14725_) & (~new_n12870_ | ~new_n18754_ | new_n14725_);
  assign new_n18754_ = new_n12737_ & new_n16652_;
  assign new_n18755_ = new_n18774_ & (new_n18778_ | ~new_n18776_ | (~new_n18782_ & (~new_n18783_ | ~new_n18756_)));
  assign new_n18756_ = ~new_n18768_ & ~new_n18770_ & (new_n18773_ | new_n18771_ | new_n18757_);
  assign new_n18757_ = new_n18767_ & ~new_n18758_ & new_n18766_;
  assign new_n18758_ = new_n18759_ & new_n18761_ & (new_n18764_ | ~\all_features[973]  | ~\all_features[974]  | ~\all_features[975] );
  assign new_n18759_ = \all_features[975]  & (\all_features[974]  | (new_n18760_ & (\all_features[970]  | \all_features[971]  | \all_features[969] )));
  assign new_n18760_ = \all_features[972]  & \all_features[973] ;
  assign new_n18761_ = \all_features[974]  & \all_features[975]  & (\all_features[972]  | \all_features[973]  | new_n18762_ | ~new_n18763_);
  assign new_n18762_ = \all_features[968]  & \all_features[969] ;
  assign new_n18763_ = ~\all_features[970]  & ~\all_features[971] ;
  assign new_n18764_ = ~\all_features[971]  & ~\all_features[972]  & (~\all_features[970]  | new_n18765_);
  assign new_n18765_ = ~\all_features[968]  & ~\all_features[969] ;
  assign new_n18766_ = \all_features[975]  & (\all_features[974]  | (\all_features[973]  & (\all_features[972]  | ~new_n18763_ | ~new_n18765_)));
  assign new_n18767_ = \all_features[975]  & (\all_features[973]  | \all_features[974]  | \all_features[972] );
  assign new_n18768_ = ~\all_features[975]  & (~\all_features[974]  | (~\all_features[972]  & ~\all_features[973]  & ~new_n18769_));
  assign new_n18769_ = \all_features[970]  & \all_features[971] ;
  assign new_n18770_ = ~\all_features[975]  & (~\all_features[974]  | (~\all_features[973]  & (new_n18765_ | ~\all_features[972]  | ~new_n18769_)));
  assign new_n18771_ = ~new_n18772_ & ~\all_features[975] ;
  assign new_n18772_ = \all_features[973]  & \all_features[974]  & (\all_features[972]  | (\all_features[970]  & \all_features[971]  & \all_features[969] ));
  assign new_n18773_ = ~\all_features[975]  & (~\all_features[974]  | ~new_n18762_ | ~new_n18760_ | ~new_n18769_);
  assign new_n18774_ = new_n18782_ | ~new_n18775_;
  assign new_n18775_ = ~new_n18778_ & new_n18776_;
  assign new_n18776_ = \all_features[973]  | \all_features[974]  | \all_features[975]  | (\all_features[972]  & \all_features[971]  & ~new_n18777_);
  assign new_n18777_ = ~\all_features[970]  & new_n18765_;
  assign new_n18778_ = ~\all_features[975]  & ~new_n18779_ & ~\all_features[974] ;
  assign new_n18779_ = \all_features[973]  & (\all_features[972]  | (\all_features[971]  & (\all_features[970]  | \all_features[969] )));
  assign new_n18780_ = ~new_n18768_ & ~new_n18773_;
  assign new_n18782_ = ~\all_features[974]  & ~\all_features[975]  & (~\all_features[971]  | ~new_n18760_ | (~\all_features[970]  & ~new_n18762_));
  assign new_n18783_ = ~new_n18768_ & (new_n18770_ | (~new_n18784_ & ~new_n18771_));
  assign new_n18784_ = ~new_n18773_ & (~new_n18767_ | (new_n18766_ & (~new_n18759_ | (~new_n18785_ & new_n18761_))));
  assign new_n18785_ = \all_features[974]  & \all_features[975]  & (\all_features[973]  | (~new_n18763_ & \all_features[972] ));
  assign new_n18786_ = ~new_n14338_ & new_n13014_;
  assign new_n18787_ = ~new_n18789_ & (new_n18788_ | new_n8739_) & (new_n18706_ | ~new_n18669_ | ~new_n18739_ | ~new_n8739_);
  assign new_n18788_ = (~new_n18223_ | ~new_n18755_ | ~new_n14725_) & (new_n14725_ | (new_n12870_ ? new_n18754_ : new_n18786_));
  assign new_n18789_ = new_n18749_ & (new_n18751_ ? new_n18750_ : new_n12398_);
  assign new_n18790_ = ~new_n18791_ & new_n18848_;
  assign new_n18791_ = ~new_n18811_ & ~new_n18792_ & new_n18799_ & (~new_n18814_ | ~new_n18813_);
  assign new_n18792_ = new_n18793_ & (new_n18797_ ? ~new_n18796_ : new_n12374_);
  assign new_n18793_ = ~new_n16775_ & new_n18794_;
  assign new_n18794_ = ~new_n18795_ & new_n6949_;
  assign new_n18795_ = new_n6921_ & new_n6945_;
  assign new_n18796_ = ~new_n15554_ & ~new_n15587_;
  assign new_n18797_ = ~new_n11301_ & (~new_n11274_ | new_n18798_);
  assign new_n18798_ = ~new_n11297_ & ~new_n13768_;
  assign new_n18799_ = (~new_n18801_ | new_n10343_) & (~new_n6879_ | ~new_n18803_ | ~new_n18800_);
  assign new_n18800_ = new_n16775_ & new_n8923_;
  assign new_n18801_ = new_n16775_ & ~new_n8923_ & new_n18802_;
  assign new_n18802_ = new_n17636_ & (~new_n17667_ | ~new_n17663_);
  assign new_n18803_ = ~new_n11000_ & (new_n18804_ | new_n11015_ | ~new_n11016_);
  assign new_n18804_ = new_n18810_ & (new_n11009_ | (~new_n11002_ & new_n18805_ & (new_n11005_ | new_n18808_)));
  assign new_n18805_ = ~new_n11005_ & ~new_n11007_ & (~new_n11022_ | ~new_n11017_ | new_n18806_);
  assign new_n18806_ = new_n11019_ & ~new_n18807_ & new_n11020_;
  assign new_n18807_ = new_n11021_ & \all_features[2741]  & ((~new_n11004_ & \all_features[2738] ) | \all_features[2740]  | \all_features[2739] );
  assign new_n18808_ = ~new_n11007_ & (~new_n11022_ | (new_n11017_ & (~new_n11019_ | (~new_n18809_ & new_n11020_))));
  assign new_n18809_ = new_n11021_ & (\all_features[2741]  | (~new_n11018_ & \all_features[2740] ));
  assign new_n18810_ = ~new_n11014_ & ~new_n11011_ & ~new_n11013_;
  assign new_n18811_ = new_n16775_ & ((~new_n8740_ & ~new_n18802_ & ~new_n8923_) | (~new_n6879_ & ~new_n18812_ & new_n8923_));
  assign new_n18812_ = ~new_n6732_ & ~new_n6734_;
  assign new_n18813_ = ~new_n16775_ & ~new_n18794_;
  assign new_n18814_ = new_n18815_ & (new_n18256_ | (new_n18225_ & new_n18249_ & new_n18253_));
  assign new_n18815_ = ~new_n18816_ & new_n18843_;
  assign new_n18816_ = ~new_n18842_ & (~new_n18835_ | (~new_n18840_ & (new_n18833_ | new_n18841_ | ~new_n18817_)));
  assign new_n18817_ = ~new_n18829_ & ~new_n18827_ & ((~new_n18824_ & new_n18818_) | ~new_n18832_ | ~new_n18831_);
  assign new_n18818_ = \all_features[5119]  & \all_features[5118]  & ~new_n18821_ & new_n18819_;
  assign new_n18819_ = \all_features[5119]  & (\all_features[5118]  | (new_n18820_ & (\all_features[5114]  | \all_features[5115]  | \all_features[5113] )));
  assign new_n18820_ = \all_features[5116]  & \all_features[5117] ;
  assign new_n18821_ = new_n18823_ & ~\all_features[5117]  & ~new_n18822_ & ~\all_features[5116] ;
  assign new_n18822_ = \all_features[5112]  & \all_features[5113] ;
  assign new_n18823_ = ~\all_features[5114]  & ~\all_features[5115] ;
  assign new_n18824_ = \all_features[5119]  & \all_features[5118]  & ~new_n18825_ & \all_features[5117] ;
  assign new_n18825_ = ~\all_features[5115]  & ~\all_features[5116]  & (~\all_features[5114]  | new_n18826_);
  assign new_n18826_ = ~\all_features[5112]  & ~\all_features[5113] ;
  assign new_n18827_ = ~new_n18828_ & ~\all_features[5119] ;
  assign new_n18828_ = \all_features[5117]  & \all_features[5118]  & (\all_features[5116]  | (\all_features[5114]  & \all_features[5115]  & \all_features[5113] ));
  assign new_n18829_ = ~\all_features[5119]  & (~\all_features[5118]  | ~new_n18830_ | ~new_n18822_ | ~new_n18820_);
  assign new_n18830_ = \all_features[5114]  & \all_features[5115] ;
  assign new_n18831_ = \all_features[5119]  & (\all_features[5118]  | (\all_features[5117]  & (\all_features[5116]  | ~new_n18823_ | ~new_n18826_)));
  assign new_n18832_ = \all_features[5119]  & (\all_features[5117]  | \all_features[5118]  | \all_features[5116] );
  assign new_n18833_ = ~new_n18827_ & (new_n18829_ | (new_n18832_ & (~new_n18831_ | (~new_n18834_ & new_n18819_))));
  assign new_n18834_ = ~\all_features[5117]  & \all_features[5118]  & \all_features[5119]  & (\all_features[5116]  ? new_n18823_ : (new_n18822_ | ~new_n18823_));
  assign new_n18835_ = ~new_n18839_ & ~new_n18836_ & ~new_n18838_;
  assign new_n18836_ = new_n18837_ & (~\all_features[5117]  | (~\all_features[5116]  & (~\all_features[5115]  | (~\all_features[5114]  & ~\all_features[5113] ))));
  assign new_n18837_ = ~\all_features[5118]  & ~\all_features[5119] ;
  assign new_n18838_ = ~\all_features[5117]  & new_n18837_ & ((~\all_features[5114]  & new_n18826_) | ~\all_features[5116]  | ~\all_features[5115] );
  assign new_n18839_ = new_n18837_ & (~\all_features[5115]  | ~new_n18820_ | (~\all_features[5114]  & ~new_n18822_));
  assign new_n18840_ = ~\all_features[5119]  & (~\all_features[5118]  | (~\all_features[5116]  & ~\all_features[5117]  & ~new_n18830_));
  assign new_n18841_ = ~\all_features[5119]  & (~\all_features[5118]  | (~\all_features[5117]  & (new_n18826_ | ~\all_features[5116]  | ~new_n18830_)));
  assign new_n18842_ = ~\all_features[5119]  & ~\all_features[5118]  & ~\all_features[5117]  & ~\all_features[5115]  & ~\all_features[5116] ;
  assign new_n18843_ = new_n18836_ | ~new_n18846_ | ((new_n18827_ | ~new_n18847_) & (new_n18844_ | new_n18839_));
  assign new_n18844_ = new_n18845_ & (~new_n18818_ | ~new_n18831_ | ~new_n18832_);
  assign new_n18845_ = ~new_n18829_ & ~new_n18827_ & ~new_n18840_ & ~new_n18841_;
  assign new_n18846_ = ~new_n18838_ & ~new_n18842_;
  assign new_n18847_ = ~new_n18839_ & ~new_n18829_ & ~new_n18840_ & ~new_n18841_;
  assign new_n18848_ = ~new_n18849_ & new_n18850_ & (new_n18851_ | new_n18814_ | ~new_n18813_);
  assign new_n18849_ = new_n18793_ & (new_n18797_ ? new_n18796_ : ~new_n12374_);
  assign new_n18850_ = (~new_n10343_ | ~new_n18801_) & (~new_n18800_ | (new_n6879_ ? new_n18803_ : ~new_n18812_));
  assign new_n18851_ = ~new_n18815_ & new_n15441_ & (new_n15437_ | (new_n15409_ & new_n15433_));
  assign new_n18852_ = ~new_n18904_ & new_n18853_;
  assign new_n18853_ = ~new_n18900_ & new_n18854_ & (~new_n18901_ | (new_n8776_ & new_n18902_) | (new_n16106_ & ~new_n18902_));
  assign new_n18854_ = (~new_n10241_ | ~new_n18892_ | (~new_n18891_ & ~new_n18856_)) & (~new_n18855_ | new_n18899_ | new_n18892_);
  assign new_n18855_ = ~new_n7600_ & ~new_n18751_;
  assign new_n18856_ = new_n15167_ & new_n18857_;
  assign new_n18857_ = ~new_n18858_ & new_n18887_;
  assign new_n18858_ = new_n18881_ & (new_n18886_ | new_n18859_);
  assign new_n18859_ = ~new_n18879_ & ~new_n18873_ & ~new_n18860_ & ~new_n18880_ & (new_n18875_ | new_n18877_);
  assign new_n18860_ = new_n18872_ & (~new_n18870_ | (~new_n18861_ & new_n18864_));
  assign new_n18861_ = \all_features[5095]  & \all_features[5094]  & ~new_n18862_ & \all_features[5093] ;
  assign new_n18862_ = ~\all_features[5091]  & ~\all_features[5092]  & (~\all_features[5090]  | new_n18863_);
  assign new_n18863_ = ~\all_features[5088]  & ~\all_features[5089] ;
  assign new_n18864_ = new_n18865_ & \all_features[5094]  & \all_features[5095]  & (~new_n18869_ | ~new_n18868_ | new_n18867_);
  assign new_n18865_ = \all_features[5095]  & (\all_features[5094]  | (new_n18866_ & (\all_features[5090]  | \all_features[5091]  | \all_features[5089] )));
  assign new_n18866_ = \all_features[5092]  & \all_features[5093] ;
  assign new_n18867_ = \all_features[5088]  & \all_features[5089] ;
  assign new_n18868_ = ~\all_features[5092]  & ~\all_features[5093] ;
  assign new_n18869_ = ~\all_features[5090]  & ~\all_features[5091] ;
  assign new_n18870_ = \all_features[5095]  & (\all_features[5094]  | (~new_n18868_ & new_n18871_));
  assign new_n18871_ = \all_features[5093]  & (\all_features[5092]  | ~new_n18869_ | ~new_n18863_);
  assign new_n18872_ = ~new_n18873_ & ~new_n18875_;
  assign new_n18873_ = ~new_n18874_ & ~\all_features[5095] ;
  assign new_n18874_ = \all_features[5093]  & \all_features[5094]  & (\all_features[5092]  | (\all_features[5090]  & \all_features[5091]  & \all_features[5089] ));
  assign new_n18875_ = ~\all_features[5095]  & (~\all_features[5094]  | ~new_n18867_ | ~new_n18866_ | ~new_n18876_);
  assign new_n18876_ = \all_features[5090]  & \all_features[5091] ;
  assign new_n18877_ = \all_features[5095]  & ((~new_n18878_ & \all_features[5094]  & new_n18865_) | (~new_n18868_ & ((~new_n18878_ & new_n18865_) | (~new_n18871_ & ~\all_features[5094] ))));
  assign new_n18878_ = ~\all_features[5093]  & \all_features[5094]  & \all_features[5095]  & (\all_features[5092]  ? new_n18869_ : (new_n18867_ | ~new_n18869_));
  assign new_n18879_ = ~\all_features[5095]  & (~\all_features[5094]  | (~\all_features[5093]  & (new_n18863_ | ~\all_features[5092]  | ~new_n18876_)));
  assign new_n18880_ = ~\all_features[5095]  & (~\all_features[5094]  | (~new_n18876_ & new_n18868_));
  assign new_n18881_ = ~new_n18884_ & new_n18882_;
  assign new_n18882_ = \all_features[5093]  | \all_features[5094]  | \all_features[5095]  | (\all_features[5092]  & \all_features[5091]  & ~new_n18883_);
  assign new_n18883_ = ~\all_features[5090]  & new_n18863_;
  assign new_n18884_ = ~\all_features[5095]  & ~new_n18885_ & ~\all_features[5094] ;
  assign new_n18885_ = \all_features[5093]  & (\all_features[5092]  | (\all_features[5091]  & (\all_features[5090]  | \all_features[5089] )));
  assign new_n18886_ = ~\all_features[5094]  & ~\all_features[5095]  & (~\all_features[5091]  | ~new_n18866_ | (~\all_features[5090]  & ~new_n18867_));
  assign new_n18887_ = ~new_n18888_ & ~new_n18890_;
  assign new_n18888_ = new_n18882_ & ~new_n18884_ & ~new_n18889_ & ~new_n18886_;
  assign new_n18889_ = ~new_n18879_ & ~new_n18873_ & ~new_n18875_ & ~new_n18880_ & (~new_n18870_ | ~new_n18864_);
  assign new_n18890_ = new_n18881_ & new_n18872_ & ~new_n18880_ & ~new_n18886_ & ~new_n18879_;
  assign new_n18891_ = ~new_n15167_ & ~\all_features[3342]  & ~\all_features[3343]  & (~\all_features[3341]  | (~\all_features[3339]  & ~\all_features[3340] ));
  assign new_n18892_ = new_n18893_ & new_n18894_;
  assign new_n18893_ = ~new_n12762_ & ~new_n12791_;
  assign new_n18894_ = ~new_n12784_ & ~new_n18895_;
  assign new_n18895_ = ~new_n18896_ & (\all_features[4339]  | \all_features[4340]  | \all_features[4341]  | \all_features[4342]  | \all_features[4343] );
  assign new_n18896_ = ~new_n12780_ & (new_n12782_ | (~new_n12783_ & (new_n12773_ | (~new_n12765_ & ~new_n18897_))));
  assign new_n18897_ = ~new_n12768_ & (new_n12770_ | (new_n12778_ & (~new_n12774_ | (~new_n18898_ & new_n12776_))));
  assign new_n18898_ = ~\all_features[4341]  & \all_features[4342]  & \all_features[4343]  & (\all_features[4340]  ? new_n12775_ : (new_n12772_ | ~new_n12775_));
  assign new_n18899_ = ~new_n9548_ & ~new_n7475_;
  assign new_n18900_ = ~new_n18892_ & ((new_n15022_ & new_n18578_ & new_n18899_) | (~new_n14426_ & new_n7600_ & ~new_n18899_));
  assign new_n18901_ = ~new_n10241_ & new_n18892_;
  assign new_n18902_ = new_n18903_ & new_n15864_;
  assign new_n18903_ = ~new_n11239_ & ~new_n11260_;
  assign new_n18904_ = ~new_n18905_ & new_n18906_ & ((new_n15022_ & new_n18578_) | ~new_n18899_ | new_n18892_);
  assign new_n18905_ = new_n18902_ & new_n18901_ & new_n8776_;
  assign new_n18906_ = (new_n18907_ | ~new_n18892_) & (new_n18899_ | new_n18892_ | (new_n7600_ ? ~new_n14426_ : ~new_n18751_));
  assign new_n18907_ = (new_n18857_ | ~new_n15167_ | ~new_n10241_) & (new_n18902_ | ~new_n16106_ | new_n10241_);
  assign new_n18908_ = ~new_n18909_ & new_n18955_;
  assign new_n18909_ = ~new_n18910_ & (~new_n18755_ | (~new_n18917_ & new_n18954_ & new_n18919_) | (new_n18915_ & ~new_n18919_));
  assign new_n18910_ = ~new_n18755_ & new_n18189_ & (new_n18913_ ? ~new_n18914_ : ~new_n18911_);
  assign new_n18911_ = new_n12491_ & new_n18912_;
  assign new_n18912_ = ~new_n12523_ & ~new_n12525_;
  assign new_n18913_ = ~new_n15599_ & new_n15628_;
  assign new_n18914_ = ~new_n12006_ & (~new_n16653_ | ~new_n12030_);
  assign new_n18915_ = ~new_n13475_ & new_n18916_;
  assign new_n18916_ = ~new_n16345_ & new_n10001_;
  assign new_n18917_ = ~new_n13808_ & new_n18918_;
  assign new_n18918_ = ~new_n13838_ & ~new_n13840_;
  assign new_n18919_ = new_n18950_ & new_n18920_ & new_n18941_;
  assign new_n18920_ = ~new_n18921_ & (\all_features[1259]  | \all_features[1260]  | \all_features[1261]  | \all_features[1262]  | \all_features[1263] );
  assign new_n18921_ = ~new_n18935_ & (new_n18937_ | (~new_n18938_ & (new_n18939_ | (~new_n18922_ & ~new_n18940_))));
  assign new_n18922_ = ~new_n18923_ & (new_n18925_ | (new_n18934_ & (~new_n18929_ | (~new_n18933_ & new_n18932_))));
  assign new_n18923_ = ~new_n18924_ & ~\all_features[1263] ;
  assign new_n18924_ = \all_features[1261]  & \all_features[1262]  & (\all_features[1260]  | (\all_features[1258]  & \all_features[1259]  & \all_features[1257] ));
  assign new_n18925_ = ~\all_features[1263]  & (~\all_features[1262]  | ~new_n18926_ | ~new_n18927_ | ~new_n18928_);
  assign new_n18926_ = \all_features[1256]  & \all_features[1257] ;
  assign new_n18927_ = \all_features[1260]  & \all_features[1261] ;
  assign new_n18928_ = \all_features[1258]  & \all_features[1259] ;
  assign new_n18929_ = \all_features[1263]  & (\all_features[1262]  | (\all_features[1261]  & (\all_features[1260]  | ~new_n18931_ | ~new_n18930_)));
  assign new_n18930_ = ~\all_features[1256]  & ~\all_features[1257] ;
  assign new_n18931_ = ~\all_features[1258]  & ~\all_features[1259] ;
  assign new_n18932_ = \all_features[1263]  & (\all_features[1262]  | (new_n18927_ & (\all_features[1258]  | \all_features[1259]  | \all_features[1257] )));
  assign new_n18933_ = ~\all_features[1261]  & \all_features[1262]  & \all_features[1263]  & (\all_features[1260]  ? new_n18931_ : (new_n18926_ | ~new_n18931_));
  assign new_n18934_ = \all_features[1263]  & (\all_features[1261]  | \all_features[1262]  | \all_features[1260] );
  assign new_n18935_ = ~\all_features[1261]  & new_n18936_ & ((~\all_features[1258]  & new_n18930_) | ~\all_features[1260]  | ~\all_features[1259] );
  assign new_n18936_ = ~\all_features[1262]  & ~\all_features[1263] ;
  assign new_n18937_ = new_n18936_ & (~\all_features[1261]  | (~\all_features[1260]  & (~\all_features[1259]  | (~\all_features[1258]  & ~\all_features[1257] ))));
  assign new_n18938_ = new_n18936_ & (~\all_features[1259]  | ~new_n18927_ | (~\all_features[1258]  & ~new_n18926_));
  assign new_n18939_ = ~\all_features[1263]  & (~\all_features[1262]  | (~\all_features[1260]  & ~\all_features[1261]  & ~new_n18928_));
  assign new_n18940_ = ~\all_features[1263]  & (~\all_features[1262]  | (~\all_features[1261]  & (new_n18930_ | ~new_n18928_ | ~\all_features[1260] )));
  assign new_n18941_ = new_n18949_ & (~new_n18947_ | (~new_n18942_ & new_n18948_));
  assign new_n18942_ = new_n18945_ & ((~new_n18943_ & new_n18932_ & new_n18946_) | ~new_n18934_ | ~new_n18929_);
  assign new_n18943_ = \all_features[1263]  & \all_features[1262]  & ~new_n18944_ & \all_features[1261] ;
  assign new_n18944_ = ~\all_features[1259]  & ~\all_features[1260]  & (~\all_features[1258]  | new_n18930_);
  assign new_n18945_ = ~new_n18923_ & ~new_n18925_;
  assign new_n18946_ = \all_features[1262]  & \all_features[1263]  & (\all_features[1260]  | \all_features[1261]  | new_n18926_ | ~new_n18931_);
  assign new_n18947_ = ~new_n18937_ & ~new_n18938_;
  assign new_n18948_ = ~new_n18939_ & ~new_n18940_;
  assign new_n18949_ = ~new_n18935_ & (\all_features[1259]  | \all_features[1260]  | \all_features[1261]  | \all_features[1262]  | \all_features[1263] );
  assign new_n18950_ = new_n18951_ & new_n18953_;
  assign new_n18951_ = new_n18947_ & new_n18949_ & (~new_n18945_ | ~new_n18948_ | (new_n18952_ & new_n18929_));
  assign new_n18952_ = new_n18934_ & new_n18932_ & new_n18946_;
  assign new_n18953_ = new_n18949_ & new_n18947_ & ~new_n18925_ & ~new_n18923_ & ~new_n18939_ & ~new_n18940_;
  assign new_n18954_ = ~new_n15628_ & ~new_n16144_ & ~new_n15600_ & ~new_n15623_;
  assign new_n18955_ = new_n18755_ ? ((new_n18917_ | ~new_n18954_ | ~new_n18919_) & (~new_n18915_ | new_n18919_)) : new_n18956_;
  assign new_n18956_ = new_n18189_ & (~new_n18914_ | ~new_n18913_);
  assign new_n18957_ = ~new_n18958_ & new_n19028_;
  assign new_n18958_ = ~new_n18959_ & ~new_n18987_ & ~new_n19022_ & (new_n18395_ | new_n19026_ | ~new_n19025_);
  assign new_n18959_ = new_n18960_ & (new_n15867_ ? new_n7162_ : new_n18961_);
  assign new_n18960_ = ~new_n9869_ & new_n17675_;
  assign new_n18961_ = ~new_n18962_ & ~new_n18985_;
  assign new_n18962_ = new_n18980_ & ~new_n18984_ & ~new_n18963_ & ~new_n18983_;
  assign new_n18963_ = ~new_n18978_ & ~new_n18979_ & new_n18971_ & (~new_n18976_ | ~new_n18964_);
  assign new_n18964_ = new_n18970_ & new_n18965_ & new_n18967_;
  assign new_n18965_ = \all_features[2847]  & (\all_features[2846]  | (new_n18966_ & (\all_features[2842]  | \all_features[2843]  | \all_features[2841] )));
  assign new_n18966_ = \all_features[2844]  & \all_features[2845] ;
  assign new_n18967_ = \all_features[2846]  & \all_features[2847]  & (\all_features[2844]  | \all_features[2845]  | new_n18969_ | ~new_n18968_);
  assign new_n18968_ = ~\all_features[2842]  & ~\all_features[2843] ;
  assign new_n18969_ = \all_features[2840]  & \all_features[2841] ;
  assign new_n18970_ = \all_features[2847]  & (\all_features[2845]  | \all_features[2846]  | \all_features[2844] );
  assign new_n18971_ = ~new_n18972_ & ~new_n18974_;
  assign new_n18972_ = ~new_n18973_ & ~\all_features[2847] ;
  assign new_n18973_ = \all_features[2845]  & \all_features[2846]  & (\all_features[2844]  | (\all_features[2842]  & \all_features[2843]  & \all_features[2841] ));
  assign new_n18974_ = ~\all_features[2847]  & (~\all_features[2846]  | (~\all_features[2844]  & ~\all_features[2845]  & ~new_n18975_));
  assign new_n18975_ = \all_features[2842]  & \all_features[2843] ;
  assign new_n18976_ = \all_features[2847]  & (\all_features[2846]  | (\all_features[2845]  & (\all_features[2844]  | ~new_n18977_ | ~new_n18968_)));
  assign new_n18977_ = ~\all_features[2840]  & ~\all_features[2841] ;
  assign new_n18978_ = ~\all_features[2847]  & (~\all_features[2846]  | (~\all_features[2845]  & (new_n18977_ | ~new_n18975_ | ~\all_features[2844] )));
  assign new_n18979_ = ~\all_features[2847]  & (~\all_features[2846]  | ~new_n18966_ | ~new_n18969_ | ~new_n18975_);
  assign new_n18980_ = ~new_n18981_ & (\all_features[2843]  | \all_features[2844]  | \all_features[2845]  | \all_features[2846]  | \all_features[2847] );
  assign new_n18981_ = ~\all_features[2845]  & new_n18982_ & ((~\all_features[2842]  & new_n18977_) | ~\all_features[2844]  | ~\all_features[2843] );
  assign new_n18982_ = ~\all_features[2846]  & ~\all_features[2847] ;
  assign new_n18983_ = new_n18982_ & (~\all_features[2845]  | (~\all_features[2844]  & (~\all_features[2843]  | (~\all_features[2842]  & ~\all_features[2841] ))));
  assign new_n18984_ = new_n18982_ & (~\all_features[2843]  | ~new_n18966_ | (~\all_features[2842]  & ~new_n18969_));
  assign new_n18985_ = new_n18980_ & new_n18971_ & new_n18986_ & ~new_n18978_ & ~new_n18979_;
  assign new_n18986_ = ~new_n18983_ & ~new_n18984_;
  assign new_n18987_ = new_n18988_ & (new_n18989_ ? new_n8267_ : new_n13134_);
  assign new_n18988_ = new_n9869_ & new_n17675_;
  assign new_n18989_ = ~new_n19018_ & new_n18990_;
  assign new_n18990_ = ~new_n18991_ & ~new_n19017_;
  assign new_n18991_ = new_n19004_ & (~new_n18992_ | (new_n19015_ & new_n19016_ & new_n19012_ & new_n19013_));
  assign new_n18992_ = new_n18993_ & new_n19000_;
  assign new_n18993_ = ~new_n18994_ & ~new_n18996_;
  assign new_n18994_ = ~new_n18995_ & ~\all_features[2527] ;
  assign new_n18995_ = \all_features[2525]  & \all_features[2526]  & (\all_features[2524]  | (\all_features[2522]  & \all_features[2523]  & \all_features[2521] ));
  assign new_n18996_ = ~\all_features[2527]  & (~\all_features[2526]  | ~new_n18997_ | ~new_n18998_ | ~new_n18999_);
  assign new_n18997_ = \all_features[2524]  & \all_features[2525] ;
  assign new_n18998_ = \all_features[2520]  & \all_features[2521] ;
  assign new_n18999_ = \all_features[2522]  & \all_features[2523] ;
  assign new_n19000_ = ~new_n19001_ & ~new_n19002_;
  assign new_n19001_ = ~\all_features[2527]  & (~\all_features[2526]  | (~\all_features[2524]  & ~\all_features[2525]  & ~new_n18999_));
  assign new_n19002_ = ~\all_features[2527]  & (~\all_features[2526]  | (~\all_features[2525]  & (new_n19003_ | ~new_n18999_ | ~\all_features[2524] )));
  assign new_n19003_ = ~\all_features[2520]  & ~\all_features[2521] ;
  assign new_n19004_ = new_n19005_ & new_n19009_;
  assign new_n19005_ = ~new_n19006_ & ~new_n19008_;
  assign new_n19006_ = new_n19007_ & (~\all_features[2525]  | (~\all_features[2524]  & (~\all_features[2523]  | (~\all_features[2522]  & ~\all_features[2521] ))));
  assign new_n19007_ = ~\all_features[2526]  & ~\all_features[2527] ;
  assign new_n19008_ = new_n19007_ & (~\all_features[2523]  | ~new_n18997_ | (~\all_features[2522]  & ~new_n18998_));
  assign new_n19009_ = ~new_n19010_ & ~new_n19011_;
  assign new_n19010_ = ~\all_features[2525]  & new_n19007_ & ((~\all_features[2522]  & new_n19003_) | ~\all_features[2524]  | ~\all_features[2523] );
  assign new_n19011_ = ~\all_features[2527]  & ~\all_features[2526]  & ~\all_features[2525]  & ~\all_features[2523]  & ~\all_features[2524] ;
  assign new_n19012_ = \all_features[2527]  & (\all_features[2526]  | (new_n18997_ & (\all_features[2522]  | \all_features[2523]  | \all_features[2521] )));
  assign new_n19013_ = \all_features[2526]  & \all_features[2527]  & (\all_features[2524]  | \all_features[2525]  | new_n18998_ | ~new_n19014_);
  assign new_n19014_ = ~\all_features[2522]  & ~\all_features[2523] ;
  assign new_n19015_ = \all_features[2527]  & (\all_features[2526]  | (\all_features[2525]  & (\all_features[2524]  | ~new_n19014_ | ~new_n19003_)));
  assign new_n19016_ = \all_features[2527]  & (\all_features[2525]  | \all_features[2526]  | \all_features[2524] );
  assign new_n19017_ = new_n18992_ & new_n19004_;
  assign new_n19018_ = new_n19009_ & (~new_n19005_ | (~new_n19019_ & new_n19000_));
  assign new_n19019_ = new_n18993_ & ((~new_n19020_ & new_n19013_ & new_n19012_) | ~new_n19016_ | ~new_n19015_);
  assign new_n19020_ = \all_features[2527]  & \all_features[2526]  & ~new_n19021_ & \all_features[2525] ;
  assign new_n19021_ = ~\all_features[2523]  & ~\all_features[2524]  & (~\all_features[2522]  | new_n19003_);
  assign new_n19022_ = ~new_n17675_ & ((new_n8201_ & new_n18395_ & new_n19024_) | (~new_n19023_ & new_n18574_ & ~new_n19024_));
  assign new_n19023_ = new_n17659_ & (new_n17637_ | ~new_n17662_);
  assign new_n19024_ = ~new_n6953_ & (~new_n6950_ | new_n6920_);
  assign new_n19025_ = ~new_n17675_ & new_n19024_;
  assign new_n19026_ = new_n12525_ & new_n19027_ & new_n12523_;
  assign new_n19027_ = new_n12492_ & new_n12514_;
  assign new_n19028_ = ~new_n19030_ & new_n19029_ & (~new_n18960_ | (new_n7162_ & new_n15867_) | (new_n18961_ & ~new_n15867_));
  assign new_n19029_ = (new_n18989_ | new_n13134_ | ~new_n18988_) & (new_n8201_ | ~new_n19025_ | ~new_n18395_);
  assign new_n19030_ = ~new_n17675_ & ~new_n19024_ & (new_n19023_ ? ~new_n8667_ : ~new_n18574_);
  assign new_n19031_ = new_n19032_ ? (~new_n19502_ ^ new_n19593_) : (new_n19502_ ^ new_n19593_);
  assign new_n19032_ = new_n19033_ ? (~new_n19334_ ^ new_n19419_) : (new_n19334_ ^ new_n19419_);
  assign new_n19033_ = new_n19034_ ? (~new_n19133_ ^ new_n17671_) : (new_n19133_ ^ new_n17671_);
  assign new_n19034_ = ~new_n19035_ & new_n19131_;
  assign new_n19035_ = ~new_n19093_ & new_n19036_ & (~new_n19054_ | ~new_n19055_) & (~new_n19092_ | ~new_n19129_);
  assign new_n19036_ = (new_n19058_ | ~new_n19037_) & (~new_n19056_ | ~new_n19091_) & (new_n19089_ | ~new_n19053_);
  assign new_n19037_ = new_n19038_ & new_n19048_;
  assign new_n19038_ = new_n19039_ & new_n19047_;
  assign new_n19039_ = ~new_n19040_ & new_n19046_;
  assign new_n19040_ = new_n19041_ & new_n10805_;
  assign new_n19041_ = (new_n19042_ | (new_n10829_ & (~\all_features[1659]  | ~\all_features[1660]  | (~\all_features[1658]  & new_n10809_)))) & (~new_n10829_ | \all_features[1659]  | \all_features[1660] );
  assign new_n19042_ = ~new_n10818_ & (new_n10817_ | (~new_n10821_ & (new_n10823_ | (~new_n19043_ & ~new_n10826_))));
  assign new_n19043_ = ~new_n10825_ & (~\all_features[1663]  | new_n19044_ | (~\all_features[1660]  & ~\all_features[1661]  & ~\all_features[1662] ));
  assign new_n19044_ = \all_features[1663]  & ((~new_n19045_ & ~\all_features[1661]  & \all_features[1662] ) | (~new_n10811_ & (\all_features[1662]  | (~new_n10808_ & \all_features[1661] ))));
  assign new_n19045_ = (\all_features[1660]  & (\all_features[1658]  | \all_features[1659] )) | (~new_n10814_ & ~\all_features[1658]  & ~\all_features[1659]  & ~\all_features[1660] );
  assign new_n19046_ = ~new_n10830_ & ~new_n10833_;
  assign new_n19047_ = new_n13038_ & (new_n14339_ | new_n13015_);
  assign new_n19048_ = new_n11373_ & (~new_n19049_ | ~new_n11629_);
  assign new_n19049_ = ~new_n19050_ & (\all_features[3075]  | \all_features[3076]  | \all_features[3077]  | \all_features[3078]  | \all_features[3079] );
  assign new_n19050_ = ~new_n7044_ & (new_n7047_ | (~new_n7048_ & (new_n7057_ | (~new_n7052_ & ~new_n19051_))));
  assign new_n19051_ = ~new_n7054_ & (new_n7056_ | (new_n7062_ & (~new_n7058_ | (~new_n19052_ & new_n7060_))));
  assign new_n19052_ = ~\all_features[3077]  & \all_features[3078]  & \all_features[3079]  & (\all_features[3076]  ? new_n7059_ : (new_n7050_ | ~new_n7059_));
  assign new_n19053_ = ~new_n19055_ & new_n19054_;
  assign new_n19054_ = ~new_n19039_ & new_n19047_;
  assign new_n19055_ = new_n15485_ & new_n11096_;
  assign new_n19056_ = ~new_n19047_ & ~new_n19057_ & ~new_n17625_;
  assign new_n19057_ = new_n13921_ & (new_n13918_ | ~new_n13888_);
  assign new_n19058_ = ~new_n19085_ & new_n19059_;
  assign new_n19059_ = ~new_n19060_ & ~new_n19083_;
  assign new_n19060_ = new_n19080_ & ~new_n19061_ & new_n19077_;
  assign new_n19061_ = ~new_n19076_ & ~new_n19074_ & ~new_n19073_ & ~new_n19062_ & ~new_n19065_;
  assign new_n19062_ = ~\all_features[4111]  & (~\all_features[4110]  | new_n19063_);
  assign new_n19063_ = ~\all_features[4109]  & (new_n19064_ | ~\all_features[4107]  | ~\all_features[4108]  | ~\all_features[4106] );
  assign new_n19064_ = ~\all_features[4104]  & ~\all_features[4105] ;
  assign new_n19065_ = new_n19072_ & new_n19071_ & new_n19066_ & new_n19068_;
  assign new_n19066_ = \all_features[4111]  & (\all_features[4110]  | (new_n19067_ & (\all_features[4106]  | \all_features[4107]  | \all_features[4105] )));
  assign new_n19067_ = \all_features[4108]  & \all_features[4109] ;
  assign new_n19068_ = \all_features[4110]  & \all_features[4111]  & (\all_features[4108]  | \all_features[4109]  | new_n19070_ | ~new_n19069_);
  assign new_n19069_ = ~\all_features[4106]  & ~\all_features[4107] ;
  assign new_n19070_ = \all_features[4104]  & \all_features[4105] ;
  assign new_n19071_ = \all_features[4111]  & (\all_features[4110]  | (\all_features[4109]  & (\all_features[4108]  | ~new_n19069_ | ~new_n19064_)));
  assign new_n19072_ = \all_features[4111]  & (\all_features[4109]  | \all_features[4110]  | \all_features[4108] );
  assign new_n19073_ = ~\all_features[4111]  & (~new_n19070_ | ~\all_features[4106]  | ~\all_features[4107]  | ~\all_features[4110]  | ~new_n19067_);
  assign new_n19074_ = ~new_n19075_ & ~\all_features[4111] ;
  assign new_n19075_ = \all_features[4109]  & \all_features[4110]  & (\all_features[4108]  | (\all_features[4106]  & \all_features[4107]  & \all_features[4105] ));
  assign new_n19076_ = ~\all_features[4111]  & (~\all_features[4110]  | (~\all_features[4109]  & ~\all_features[4108]  & (~\all_features[4107]  | ~\all_features[4106] )));
  assign new_n19077_ = ~new_n19078_ & (\all_features[4107]  | \all_features[4108]  | \all_features[4109]  | \all_features[4110]  | \all_features[4111] );
  assign new_n19078_ = ~\all_features[4109]  & new_n19079_ & ((~\all_features[4106]  & new_n19064_) | ~\all_features[4108]  | ~\all_features[4107] );
  assign new_n19079_ = ~\all_features[4110]  & ~\all_features[4111] ;
  assign new_n19080_ = ~new_n19081_ & ~new_n19082_;
  assign new_n19081_ = new_n19079_ & (~\all_features[4107]  | ~new_n19067_ | (~new_n19070_ & ~\all_features[4106] ));
  assign new_n19082_ = new_n19079_ & (~\all_features[4109]  | (~\all_features[4108]  & (~\all_features[4107]  | (~\all_features[4106]  & ~\all_features[4105] ))));
  assign new_n19083_ = new_n19077_ & new_n19084_ & ~new_n19074_ & ~new_n19082_;
  assign new_n19084_ = ~new_n19076_ & ~new_n19081_ & ~new_n19062_ & ~new_n19073_;
  assign new_n19085_ = new_n19077_ & (~new_n19080_ | (~new_n19062_ & ~new_n19086_ & ~new_n19076_));
  assign new_n19086_ = ~new_n19074_ & ~new_n19073_ & (~new_n19072_ | ~new_n19071_ | new_n19087_);
  assign new_n19087_ = new_n19066_ & new_n19068_ & (new_n19088_ | ~\all_features[4109]  | ~\all_features[4110]  | ~\all_features[4111] );
  assign new_n19088_ = ~\all_features[4107]  & ~\all_features[4108]  & (~\all_features[4106]  | new_n19064_);
  assign new_n19089_ = ~new_n19090_ & ~new_n15702_;
  assign new_n19090_ = new_n15703_ & new_n15676_;
  assign new_n19091_ = new_n14723_ & (new_n14720_ | ~new_n14691_);
  assign new_n19092_ = ~new_n19048_ & new_n19038_;
  assign new_n19093_ = ~new_n19047_ & (new_n19057_ ? (new_n19095_ | ~new_n19094_) : new_n17625_);
  assign new_n19094_ = new_n14493_ & (new_n14471_ | ~new_n14494_);
  assign new_n19095_ = ~new_n19127_ & ~new_n19096_ & ~new_n19125_;
  assign new_n19096_ = new_n19097_ & new_n19118_;
  assign new_n19097_ = ~new_n19098_ & (\all_features[5443]  | \all_features[5444]  | \all_features[5445]  | \all_features[5446]  | \all_features[5447] );
  assign new_n19098_ = ~new_n19112_ & (new_n19114_ | (~new_n19115_ & (new_n19116_ | (~new_n19099_ & ~new_n19117_))));
  assign new_n19099_ = ~new_n19100_ & (new_n19102_ | (new_n19111_ & (~new_n19106_ | (~new_n19110_ & new_n19109_))));
  assign new_n19100_ = ~new_n19101_ & ~\all_features[5447] ;
  assign new_n19101_ = \all_features[5445]  & \all_features[5446]  & (\all_features[5444]  | (\all_features[5442]  & \all_features[5443]  & \all_features[5441] ));
  assign new_n19102_ = ~\all_features[5447]  & (~\all_features[5446]  | ~new_n19103_ | ~new_n19104_ | ~new_n19105_);
  assign new_n19103_ = \all_features[5440]  & \all_features[5441] ;
  assign new_n19104_ = \all_features[5444]  & \all_features[5445] ;
  assign new_n19105_ = \all_features[5442]  & \all_features[5443] ;
  assign new_n19106_ = \all_features[5447]  & (\all_features[5446]  | (\all_features[5445]  & (\all_features[5444]  | ~new_n19108_ | ~new_n19107_)));
  assign new_n19107_ = ~\all_features[5440]  & ~\all_features[5441] ;
  assign new_n19108_ = ~\all_features[5442]  & ~\all_features[5443] ;
  assign new_n19109_ = \all_features[5447]  & (\all_features[5446]  | (new_n19104_ & (\all_features[5442]  | \all_features[5443]  | \all_features[5441] )));
  assign new_n19110_ = ~\all_features[5445]  & \all_features[5446]  & \all_features[5447]  & (\all_features[5444]  ? new_n19108_ : (new_n19103_ | ~new_n19108_));
  assign new_n19111_ = \all_features[5447]  & (\all_features[5445]  | \all_features[5446]  | \all_features[5444] );
  assign new_n19112_ = ~\all_features[5445]  & new_n19113_ & ((~\all_features[5442]  & new_n19107_) | ~\all_features[5444]  | ~\all_features[5443] );
  assign new_n19113_ = ~\all_features[5446]  & ~\all_features[5447] ;
  assign new_n19114_ = new_n19113_ & (~\all_features[5445]  | (~\all_features[5444]  & (~\all_features[5443]  | (~\all_features[5442]  & ~\all_features[5441] ))));
  assign new_n19115_ = new_n19113_ & (~\all_features[5443]  | ~new_n19104_ | (~\all_features[5442]  & ~new_n19103_));
  assign new_n19116_ = ~\all_features[5447]  & (~\all_features[5446]  | (~\all_features[5444]  & ~\all_features[5445]  & ~new_n19105_));
  assign new_n19117_ = ~\all_features[5447]  & (~\all_features[5446]  | (~\all_features[5445]  & (new_n19107_ | ~new_n19105_ | ~\all_features[5444] )));
  assign new_n19118_ = new_n19123_ & (~new_n19124_ | (~new_n19119_ & ~new_n19116_ & ~new_n19117_));
  assign new_n19119_ = ~new_n19100_ & ~new_n19102_ & (~new_n19111_ | ~new_n19106_ | new_n19120_);
  assign new_n19120_ = new_n19109_ & new_n19121_ & (new_n19122_ | ~\all_features[5445]  | ~\all_features[5446]  | ~\all_features[5447] );
  assign new_n19121_ = \all_features[5446]  & \all_features[5447]  & (\all_features[5444]  | \all_features[5445]  | new_n19103_ | ~new_n19108_);
  assign new_n19122_ = ~\all_features[5443]  & ~\all_features[5444]  & (~\all_features[5442]  | new_n19107_);
  assign new_n19123_ = ~new_n19112_ & (\all_features[5443]  | \all_features[5444]  | \all_features[5445]  | \all_features[5446]  | \all_features[5447] );
  assign new_n19124_ = ~new_n19114_ & ~new_n19115_;
  assign new_n19125_ = new_n19126_ & new_n19123_ & ~new_n19100_ & ~new_n19117_ & ~new_n19114_ & ~new_n19115_;
  assign new_n19126_ = ~new_n19116_ & ~new_n19102_;
  assign new_n19127_ = new_n19123_ & new_n19124_ & (new_n19128_ | new_n19117_ | new_n19100_ | ~new_n19126_);
  assign new_n19128_ = new_n19111_ & new_n19121_ & new_n19106_ & new_n19109_;
  assign new_n19129_ = new_n19130_ & new_n7732_;
  assign new_n19130_ = new_n7701_ & new_n7722_;
  assign new_n19131_ = new_n19132_ & (new_n19091_ | ~new_n19056_) & (~new_n19058_ | ~new_n19037_);
  assign new_n19132_ = (new_n19129_ | ~new_n19092_) & (~new_n19053_ | ~new_n19089_);
  assign new_n19133_ = new_n19134_ ? (new_n19155_ ^ new_n19242_) : (~new_n19155_ ^ new_n19242_);
  assign new_n19134_ = ~new_n19135_ & new_n19151_;
  assign new_n19135_ = new_n17217_ ? new_n19136_ : (new_n19147_ ? new_n19140_ : ~new_n19149_);
  assign new_n19136_ = ~new_n19137_ & (~new_n14294_ | new_n19138_);
  assign new_n19137_ = new_n10833_ & (new_n10830_ | new_n19040_);
  assign new_n19138_ = new_n11788_ & new_n19139_ & new_n11784_;
  assign new_n19139_ = new_n11758_ & new_n11781_;
  assign new_n19140_ = new_n9998_ ? ~new_n15477_ : ~new_n19141_;
  assign new_n19141_ = new_n8475_ & (new_n8447_ | ~new_n19142_);
  assign new_n19142_ = ~new_n8471_ & (new_n8470_ | (~new_n8469_ & (new_n8467_ | new_n19143_)));
  assign new_n19143_ = ~new_n8465_ & (new_n8458_ | (~new_n8460_ & (new_n8461_ | (~new_n19144_ & ~new_n8463_))));
  assign new_n19144_ = ~new_n19145_ & \all_features[2511]  & (\all_features[2510]  | \all_features[2509]  | \all_features[2508] );
  assign new_n19145_ = \all_features[2511]  & ((~new_n19146_ & ~\all_features[2509]  & \all_features[2510] ) | (~new_n8454_ & (\all_features[2510]  | (~new_n8450_ & \all_features[2509] ))));
  assign new_n19146_ = (\all_features[2508]  & ~new_n8452_) | (~new_n8457_ & ~\all_features[2508]  & new_n8452_);
  assign new_n19147_ = new_n13408_ & new_n19148_;
  assign new_n19148_ = ~new_n13438_ & ~new_n13441_;
  assign new_n19149_ = new_n10478_ & ~new_n17329_ & ~new_n19150_;
  assign new_n19150_ = ~new_n10456_ & ~new_n10481_;
  assign new_n19151_ = ~new_n19153_ & ~new_n19154_ & (~new_n19152_ | (new_n8741_ & new_n19138_) | (new_n14294_ & ~new_n19138_));
  assign new_n19152_ = ~new_n19137_ & new_n17217_;
  assign new_n19153_ = ~new_n17217_ & new_n19147_ & (new_n9998_ ? ~new_n15477_ : ~new_n19141_);
  assign new_n19154_ = ~new_n17217_ & ~new_n19147_ & ~new_n19149_;
  assign new_n19155_ = ~new_n19161_ & ~new_n19230_ & (new_n19240_ ? (~new_n9869_ | new_n19156_) : ~new_n19239_);
  assign new_n19156_ = new_n19160_ ? new_n18099_ : new_n19157_;
  assign new_n19157_ = new_n19158_ & new_n19159_;
  assign new_n19158_ = new_n16193_ & new_n16224_;
  assign new_n19159_ = new_n16216_ & new_n16222_;
  assign new_n19160_ = ~new_n14042_ & (~new_n14039_ | ~new_n14014_);
  assign new_n19161_ = ~new_n9869_ & ~new_n19162_ & (new_n19197_ ? ~new_n19195_ : ~new_n19196_);
  assign new_n19162_ = ~new_n19191_ & new_n19163_;
  assign new_n19163_ = ~new_n19164_ & ~new_n19190_;
  assign new_n19164_ = new_n19177_ & (~new_n19165_ | (new_n19188_ & new_n19189_ & new_n19185_ & new_n19186_));
  assign new_n19165_ = new_n19166_ & new_n19173_;
  assign new_n19166_ = ~new_n19167_ & ~new_n19169_;
  assign new_n19167_ = ~new_n19168_ & ~\all_features[4439] ;
  assign new_n19168_ = \all_features[4437]  & \all_features[4438]  & (\all_features[4436]  | (\all_features[4434]  & \all_features[4435]  & \all_features[4433] ));
  assign new_n19169_ = ~\all_features[4439]  & (~\all_features[4438]  | ~new_n19170_ | ~new_n19171_ | ~new_n19172_);
  assign new_n19170_ = \all_features[4436]  & \all_features[4437] ;
  assign new_n19171_ = \all_features[4432]  & \all_features[4433] ;
  assign new_n19172_ = \all_features[4434]  & \all_features[4435] ;
  assign new_n19173_ = ~new_n19174_ & ~new_n19175_;
  assign new_n19174_ = ~\all_features[4439]  & (~\all_features[4438]  | (~\all_features[4436]  & ~\all_features[4437]  & ~new_n19172_));
  assign new_n19175_ = ~\all_features[4439]  & (~\all_features[4438]  | (~\all_features[4437]  & (new_n19176_ | ~new_n19172_ | ~\all_features[4436] )));
  assign new_n19176_ = ~\all_features[4432]  & ~\all_features[4433] ;
  assign new_n19177_ = new_n19178_ & new_n19182_;
  assign new_n19178_ = ~new_n19179_ & ~new_n19181_;
  assign new_n19179_ = new_n19180_ & (~\all_features[4437]  | (~\all_features[4436]  & (~\all_features[4435]  | (~\all_features[4434]  & ~\all_features[4433] ))));
  assign new_n19180_ = ~\all_features[4438]  & ~\all_features[4439] ;
  assign new_n19181_ = new_n19180_ & (~\all_features[4435]  | ~new_n19170_ | (~\all_features[4434]  & ~new_n19171_));
  assign new_n19182_ = ~new_n19183_ & ~new_n19184_;
  assign new_n19183_ = ~\all_features[4437]  & new_n19180_ & ((~\all_features[4434]  & new_n19176_) | ~\all_features[4436]  | ~\all_features[4435] );
  assign new_n19184_ = ~\all_features[4439]  & ~\all_features[4438]  & ~\all_features[4437]  & ~\all_features[4435]  & ~\all_features[4436] ;
  assign new_n19185_ = \all_features[4439]  & (\all_features[4438]  | (new_n19170_ & (\all_features[4434]  | \all_features[4435]  | \all_features[4433] )));
  assign new_n19186_ = \all_features[4438]  & \all_features[4439]  & (\all_features[4436]  | \all_features[4437]  | new_n19171_ | ~new_n19187_);
  assign new_n19187_ = ~\all_features[4434]  & ~\all_features[4435] ;
  assign new_n19188_ = \all_features[4439]  & (\all_features[4438]  | (\all_features[4437]  & (\all_features[4436]  | ~new_n19187_ | ~new_n19176_)));
  assign new_n19189_ = \all_features[4439]  & (\all_features[4437]  | \all_features[4438]  | \all_features[4436] );
  assign new_n19190_ = new_n19165_ & new_n19177_;
  assign new_n19191_ = new_n19182_ & (~new_n19178_ | (~new_n19192_ & new_n19173_));
  assign new_n19192_ = new_n19166_ & ((~new_n19193_ & new_n19186_ & new_n19185_) | ~new_n19189_ | ~new_n19188_);
  assign new_n19193_ = \all_features[4439]  & \all_features[4438]  & ~new_n19194_ & \all_features[4437] ;
  assign new_n19194_ = ~\all_features[4435]  & ~\all_features[4436]  & (~\all_features[4434]  | new_n19176_);
  assign new_n19195_ = new_n13284_ & ~new_n13314_ & ~new_n13316_;
  assign new_n19196_ = new_n16607_ & (new_n16603_ | (new_n16596_ & new_n16575_));
  assign new_n19197_ = ~new_n19198_ & new_n19225_;
  assign new_n19198_ = ~new_n19224_ & (~new_n19217_ | (~new_n19222_ & (new_n19215_ | new_n19223_ | ~new_n19199_)));
  assign new_n19199_ = ~new_n19211_ & ~new_n19209_ & ((~new_n19206_ & new_n19200_) | ~new_n19214_ | ~new_n19213_);
  assign new_n19200_ = \all_features[4887]  & \all_features[4886]  & ~new_n19203_ & new_n19201_;
  assign new_n19201_ = \all_features[4887]  & (\all_features[4886]  | (new_n19202_ & (\all_features[4882]  | \all_features[4883]  | \all_features[4881] )));
  assign new_n19202_ = \all_features[4884]  & \all_features[4885] ;
  assign new_n19203_ = new_n19205_ & ~\all_features[4885]  & ~new_n19204_ & ~\all_features[4884] ;
  assign new_n19204_ = \all_features[4880]  & \all_features[4881] ;
  assign new_n19205_ = ~\all_features[4882]  & ~\all_features[4883] ;
  assign new_n19206_ = \all_features[4887]  & \all_features[4886]  & ~new_n19207_ & \all_features[4885] ;
  assign new_n19207_ = ~\all_features[4883]  & ~\all_features[4884]  & (~\all_features[4882]  | new_n19208_);
  assign new_n19208_ = ~\all_features[4880]  & ~\all_features[4881] ;
  assign new_n19209_ = ~new_n19210_ & ~\all_features[4887] ;
  assign new_n19210_ = \all_features[4885]  & \all_features[4886]  & (\all_features[4884]  | (\all_features[4882]  & \all_features[4883]  & \all_features[4881] ));
  assign new_n19211_ = ~\all_features[4887]  & (~\all_features[4886]  | ~new_n19212_ | ~new_n19204_ | ~new_n19202_);
  assign new_n19212_ = \all_features[4882]  & \all_features[4883] ;
  assign new_n19213_ = \all_features[4887]  & (\all_features[4886]  | (\all_features[4885]  & (\all_features[4884]  | ~new_n19205_ | ~new_n19208_)));
  assign new_n19214_ = \all_features[4887]  & (\all_features[4885]  | \all_features[4886]  | \all_features[4884] );
  assign new_n19215_ = ~new_n19209_ & (new_n19211_ | (new_n19214_ & (~new_n19213_ | (~new_n19216_ & new_n19201_))));
  assign new_n19216_ = ~\all_features[4885]  & \all_features[4886]  & \all_features[4887]  & (\all_features[4884]  ? new_n19205_ : (new_n19204_ | ~new_n19205_));
  assign new_n19217_ = ~new_n19221_ & ~new_n19218_ & ~new_n19220_;
  assign new_n19218_ = new_n19219_ & (~\all_features[4885]  | (~\all_features[4884]  & (~\all_features[4883]  | (~\all_features[4882]  & ~\all_features[4881] ))));
  assign new_n19219_ = ~\all_features[4886]  & ~\all_features[4887] ;
  assign new_n19220_ = ~\all_features[4885]  & new_n19219_ & ((~\all_features[4882]  & new_n19208_) | ~\all_features[4884]  | ~\all_features[4883] );
  assign new_n19221_ = new_n19219_ & (~\all_features[4883]  | ~new_n19202_ | (~\all_features[4882]  & ~new_n19204_));
  assign new_n19222_ = ~\all_features[4887]  & (~\all_features[4886]  | (~\all_features[4884]  & ~\all_features[4885]  & ~new_n19212_));
  assign new_n19223_ = ~\all_features[4887]  & (~\all_features[4886]  | (~\all_features[4885]  & (new_n19208_ | ~\all_features[4884]  | ~new_n19212_)));
  assign new_n19224_ = ~\all_features[4887]  & ~\all_features[4886]  & ~\all_features[4885]  & ~\all_features[4883]  & ~\all_features[4884] ;
  assign new_n19225_ = new_n19218_ | ~new_n19228_ | ((new_n19209_ | ~new_n19229_) & (new_n19226_ | new_n19221_));
  assign new_n19226_ = new_n19227_ & (~new_n19200_ | ~new_n19213_ | ~new_n19214_);
  assign new_n19227_ = ~new_n19211_ & ~new_n19209_ & ~new_n19222_ & ~new_n19223_;
  assign new_n19228_ = ~new_n19220_ & ~new_n19224_;
  assign new_n19229_ = ~new_n19221_ & ~new_n19211_ & ~new_n19222_ & ~new_n19223_;
  assign new_n19230_ = ~new_n9869_ & new_n19162_ & new_n19237_ & (~new_n19232_ | ~new_n19231_);
  assign new_n19231_ = new_n8545_ & new_n6955_;
  assign new_n19232_ = new_n8554_ & new_n19233_;
  assign new_n19233_ = ~new_n19234_ & (\all_features[4147]  | \all_features[4148]  | \all_features[4149]  | \all_features[4150]  | \all_features[4151] );
  assign new_n19234_ = ~new_n6971_ & (new_n6966_ | (~new_n6962_ & (new_n6957_ | (~new_n6959_ & ~new_n19235_))));
  assign new_n19235_ = ~new_n6969_ & (new_n6968_ | (new_n8552_ & (~new_n8548_ | (~new_n19236_ & new_n8550_))));
  assign new_n19236_ = ~\all_features[4149]  & \all_features[4150]  & \all_features[4151]  & (\all_features[4148]  ? new_n8549_ : (new_n6964_ | ~new_n8549_));
  assign new_n19237_ = ~new_n6974_ & new_n19238_;
  assign new_n19238_ = ~new_n6998_ & ~new_n7000_;
  assign new_n19239_ = ~new_n8667_ & new_n9869_ & (new_n18568_ | new_n18548_);
  assign new_n19240_ = new_n10271_ & (new_n10249_ | new_n19241_);
  assign new_n19241_ = new_n10273_ & new_n10277_;
  assign new_n19242_ = (~new_n19243_ & ~new_n19314_) | (~new_n19316_ & new_n19314_ & (new_n19318_ | ~new_n19278_));
  assign new_n19243_ = new_n6389_ & ((~new_n19246_ & new_n19273_) ? ~new_n19244_ : ~new_n17804_);
  assign new_n19244_ = new_n19245_ & new_n12980_;
  assign new_n19245_ = new_n12968_ & new_n12978_;
  assign new_n19246_ = ~new_n19272_ & (~new_n19265_ | (~new_n19270_ & (new_n19263_ | new_n19271_ | ~new_n19247_)));
  assign new_n19247_ = ~new_n19259_ & ~new_n19257_ & ((~new_n19254_ & new_n19248_) | ~new_n19262_ | ~new_n19261_);
  assign new_n19248_ = \all_features[1399]  & \all_features[1398]  & ~new_n19251_ & new_n19249_;
  assign new_n19249_ = \all_features[1399]  & (\all_features[1398]  | (new_n19250_ & (\all_features[1394]  | \all_features[1395]  | \all_features[1393] )));
  assign new_n19250_ = \all_features[1396]  & \all_features[1397] ;
  assign new_n19251_ = new_n19253_ & ~\all_features[1397]  & ~new_n19252_ & ~\all_features[1396] ;
  assign new_n19252_ = \all_features[1392]  & \all_features[1393] ;
  assign new_n19253_ = ~\all_features[1394]  & ~\all_features[1395] ;
  assign new_n19254_ = \all_features[1399]  & \all_features[1398]  & ~new_n19255_ & \all_features[1397] ;
  assign new_n19255_ = ~\all_features[1395]  & ~\all_features[1396]  & (~\all_features[1394]  | new_n19256_);
  assign new_n19256_ = ~\all_features[1392]  & ~\all_features[1393] ;
  assign new_n19257_ = ~new_n19258_ & ~\all_features[1399] ;
  assign new_n19258_ = \all_features[1397]  & \all_features[1398]  & (\all_features[1396]  | (\all_features[1394]  & \all_features[1395]  & \all_features[1393] ));
  assign new_n19259_ = ~\all_features[1399]  & (~\all_features[1398]  | ~new_n19260_ | ~new_n19252_ | ~new_n19250_);
  assign new_n19260_ = \all_features[1394]  & \all_features[1395] ;
  assign new_n19261_ = \all_features[1399]  & (\all_features[1398]  | (\all_features[1397]  & (\all_features[1396]  | ~new_n19253_ | ~new_n19256_)));
  assign new_n19262_ = \all_features[1399]  & (\all_features[1397]  | \all_features[1398]  | \all_features[1396] );
  assign new_n19263_ = ~new_n19257_ & (new_n19259_ | (new_n19262_ & (~new_n19261_ | (~new_n19264_ & new_n19249_))));
  assign new_n19264_ = ~\all_features[1397]  & \all_features[1398]  & \all_features[1399]  & (\all_features[1396]  ? new_n19253_ : (new_n19252_ | ~new_n19253_));
  assign new_n19265_ = ~new_n19269_ & ~new_n19266_ & ~new_n19268_;
  assign new_n19266_ = new_n19267_ & (~\all_features[1397]  | (~\all_features[1396]  & (~\all_features[1395]  | (~\all_features[1394]  & ~\all_features[1393] ))));
  assign new_n19267_ = ~\all_features[1398]  & ~\all_features[1399] ;
  assign new_n19268_ = ~\all_features[1397]  & new_n19267_ & ((~\all_features[1394]  & new_n19256_) | ~\all_features[1396]  | ~\all_features[1395] );
  assign new_n19269_ = new_n19267_ & (~\all_features[1395]  | ~new_n19250_ | (~\all_features[1394]  & ~new_n19252_));
  assign new_n19270_ = ~\all_features[1399]  & (~\all_features[1398]  | (~\all_features[1396]  & ~\all_features[1397]  & ~new_n19260_));
  assign new_n19271_ = ~\all_features[1399]  & (~\all_features[1398]  | (~\all_features[1397]  & (new_n19256_ | ~\all_features[1396]  | ~new_n19260_)));
  assign new_n19272_ = ~\all_features[1399]  & ~\all_features[1398]  & ~\all_features[1397]  & ~\all_features[1395]  & ~\all_features[1396] ;
  assign new_n19273_ = new_n19266_ | ~new_n19276_ | ((new_n19257_ | ~new_n19277_) & (new_n19274_ | new_n19269_));
  assign new_n19274_ = new_n19275_ & (~new_n19248_ | ~new_n19261_ | ~new_n19262_);
  assign new_n19275_ = ~new_n19259_ & ~new_n19257_ & ~new_n19270_ & ~new_n19271_;
  assign new_n19276_ = ~new_n19268_ & ~new_n19272_;
  assign new_n19277_ = ~new_n19269_ & ~new_n19259_ & ~new_n19270_ & ~new_n19271_;
  assign new_n19278_ = new_n19279_ & (~new_n17176_ | (~new_n19313_ & ~new_n17154_));
  assign new_n19279_ = ~new_n19309_ & (~new_n19311_ | ~new_n19280_);
  assign new_n19280_ = new_n19281_ & new_n19305_;
  assign new_n19281_ = new_n19297_ & (~new_n19300_ | (~new_n19282_ & ~new_n19303_ & ~new_n19304_));
  assign new_n19282_ = ~new_n19291_ & ~new_n19293_ & (~new_n19296_ | ~new_n19295_ | new_n19283_);
  assign new_n19283_ = new_n19284_ & new_n19286_ & (new_n19289_ | ~\all_features[4869]  | ~\all_features[4870]  | ~\all_features[4871] );
  assign new_n19284_ = \all_features[4871]  & (\all_features[4870]  | (new_n19285_ & (\all_features[4866]  | \all_features[4867]  | \all_features[4865] )));
  assign new_n19285_ = \all_features[4868]  & \all_features[4869] ;
  assign new_n19286_ = \all_features[4870]  & \all_features[4871]  & (\all_features[4868]  | \all_features[4869]  | new_n19287_ | ~new_n19288_);
  assign new_n19287_ = \all_features[4864]  & \all_features[4865] ;
  assign new_n19288_ = ~\all_features[4866]  & ~\all_features[4867] ;
  assign new_n19289_ = ~\all_features[4867]  & ~\all_features[4868]  & (~\all_features[4866]  | new_n19290_);
  assign new_n19290_ = ~\all_features[4864]  & ~\all_features[4865] ;
  assign new_n19291_ = ~new_n19292_ & ~\all_features[4871] ;
  assign new_n19292_ = \all_features[4869]  & \all_features[4870]  & (\all_features[4868]  | (\all_features[4866]  & \all_features[4867]  & \all_features[4865] ));
  assign new_n19293_ = ~\all_features[4871]  & (~\all_features[4870]  | ~new_n19294_ | ~new_n19287_ | ~new_n19285_);
  assign new_n19294_ = \all_features[4866]  & \all_features[4867] ;
  assign new_n19295_ = \all_features[4871]  & (\all_features[4870]  | (\all_features[4869]  & (\all_features[4868]  | ~new_n19288_ | ~new_n19290_)));
  assign new_n19296_ = \all_features[4871]  & (\all_features[4869]  | \all_features[4870]  | \all_features[4868] );
  assign new_n19297_ = ~new_n19298_ & (\all_features[4867]  | \all_features[4868]  | \all_features[4869]  | \all_features[4870]  | \all_features[4871] );
  assign new_n19298_ = ~\all_features[4869]  & new_n19299_ & ((~\all_features[4866]  & new_n19290_) | ~\all_features[4868]  | ~\all_features[4867] );
  assign new_n19299_ = ~\all_features[4870]  & ~\all_features[4871] ;
  assign new_n19300_ = ~new_n19301_ & ~new_n19302_;
  assign new_n19301_ = new_n19299_ & (~\all_features[4869]  | (~\all_features[4868]  & (~\all_features[4867]  | (~\all_features[4866]  & ~\all_features[4865] ))));
  assign new_n19302_ = new_n19299_ & (~\all_features[4867]  | ~new_n19285_ | (~\all_features[4866]  & ~new_n19287_));
  assign new_n19303_ = ~\all_features[4871]  & (~\all_features[4870]  | (~\all_features[4869]  & (new_n19290_ | ~new_n19294_ | ~\all_features[4868] )));
  assign new_n19304_ = ~\all_features[4871]  & (~\all_features[4870]  | (~\all_features[4868]  & ~\all_features[4869]  & ~new_n19294_));
  assign new_n19305_ = ~new_n19306_ & (\all_features[4867]  | \all_features[4868]  | \all_features[4869]  | \all_features[4870]  | \all_features[4871] );
  assign new_n19306_ = ~new_n19298_ & (new_n19301_ | (~new_n19302_ & (new_n19304_ | (~new_n19303_ & ~new_n19307_))));
  assign new_n19307_ = ~new_n19291_ & (new_n19293_ | (new_n19296_ & (~new_n19295_ | (~new_n19308_ & new_n19284_))));
  assign new_n19308_ = ~\all_features[4869]  & \all_features[4870]  & \all_features[4871]  & (\all_features[4868]  ? new_n19288_ : (new_n19287_ | ~new_n19288_));
  assign new_n19309_ = new_n19310_ & new_n19297_ & ~new_n19302_ & ~new_n19303_ & ~new_n19291_ & ~new_n19301_;
  assign new_n19310_ = ~new_n19293_ & ~new_n19304_;
  assign new_n19311_ = new_n19297_ & new_n19300_ & (new_n19312_ | new_n19291_ | new_n19303_ | ~new_n19310_);
  assign new_n19312_ = new_n19296_ & new_n19286_ & new_n19295_ & new_n19284_;
  assign new_n19313_ = new_n17178_ & new_n17182_;
  assign new_n19314_ = new_n11884_ & (new_n11861_ | ~new_n19315_);
  assign new_n19315_ = ~new_n11887_ & ~new_n11891_;
  assign new_n19316_ = new_n19317_ & (new_n7946_ | (new_n7935_ & new_n7943_));
  assign new_n19317_ = ~new_n13503_ & new_n19318_ & (~new_n13506_ | ~new_n13480_);
  assign new_n19318_ = new_n19324_ & new_n19319_ & ~new_n19333_ & ~new_n19332_ & ~new_n19328_ & ~new_n19330_;
  assign new_n19319_ = ~new_n19320_ & ~new_n19322_;
  assign new_n19320_ = new_n19321_ & ~\all_features[4197]  & ~\all_features[4195]  & ~\all_features[4196] ;
  assign new_n19321_ = ~\all_features[4198]  & ~\all_features[4199] ;
  assign new_n19322_ = ~\all_features[4199]  & (~\all_features[4198]  | (~\all_features[4196]  & ~\all_features[4197]  & ~new_n19323_));
  assign new_n19323_ = \all_features[4194]  & \all_features[4195] ;
  assign new_n19324_ = ~new_n19325_ & ~new_n19327_;
  assign new_n19325_ = new_n19321_ & (~new_n19326_ | ~\all_features[4195]  | (~\all_features[4194]  & (~\all_features[4192]  | ~\all_features[4193] )));
  assign new_n19326_ = \all_features[4196]  & \all_features[4197] ;
  assign new_n19327_ = new_n19321_ & (~\all_features[4197]  | (~\all_features[4196]  & (~\all_features[4195]  | (~\all_features[4194]  & ~\all_features[4193] ))));
  assign new_n19328_ = ~new_n19329_ & ~\all_features[4199] ;
  assign new_n19329_ = \all_features[4197]  & \all_features[4198]  & (\all_features[4196]  | (\all_features[4194]  & \all_features[4195]  & \all_features[4193] ));
  assign new_n19330_ = ~\all_features[4197]  & new_n19321_ & ((~\all_features[4194]  & new_n19331_) | ~\all_features[4196]  | ~\all_features[4195] );
  assign new_n19331_ = ~\all_features[4192]  & ~\all_features[4193] ;
  assign new_n19332_ = ~\all_features[4199]  & (~new_n19326_ | ~\all_features[4192]  | ~\all_features[4193]  | ~\all_features[4198]  | ~new_n19323_);
  assign new_n19333_ = ~\all_features[4199]  & (~\all_features[4198]  | (~\all_features[4197]  & (new_n19331_ | ~\all_features[4196]  | ~new_n19323_)));
  assign new_n19334_ = ~new_n19416_ & new_n19335_;
  assign new_n19335_ = ~new_n19336_ & new_n19346_ & (~new_n19378_ | (new_n12849_ & ~new_n19379_) | (new_n19382_ & new_n19379_));
  assign new_n19336_ = new_n19344_ & new_n19337_ & new_n19342_;
  assign new_n19337_ = ~new_n19338_ & ~new_n19339_;
  assign new_n19338_ = ~new_n17327_ & new_n11096_;
  assign new_n19339_ = ~new_n15922_ & new_n19340_;
  assign new_n19340_ = ~new_n15942_ & new_n19341_;
  assign new_n19341_ = ~new_n15951_ & ~new_n15953_;
  assign new_n19342_ = new_n10877_ & new_n19343_;
  assign new_n19343_ = ~new_n10906_ & ~new_n10908_;
  assign new_n19344_ = ~new_n14070_ & new_n19345_;
  assign new_n19345_ = ~new_n14047_ & ~new_n14077_;
  assign new_n19346_ = ~new_n19347_ | (new_n19348_ ? new_n19349_ : ~new_n19350_);
  assign new_n19347_ = ~new_n19344_ & new_n19342_;
  assign new_n19348_ = ~new_n7501_ & new_n7509_;
  assign new_n19349_ = new_n11781_ & (new_n11758_ | ~new_n11783_);
  assign new_n19350_ = ~new_n19370_ & (~new_n19371_ | (~new_n19351_ & ~new_n19375_ & ~new_n19376_ & new_n19377_));
  assign new_n19351_ = ~new_n19368_ & ~new_n19369_ & (~new_n19363_ | (new_n19352_ & (~new_n19358_ | new_n19356_)));
  assign new_n19352_ = \all_features[2215]  & (\all_features[2214]  | (~new_n19353_ & \all_features[2213] ));
  assign new_n19353_ = new_n19354_ & ~\all_features[2212]  & new_n19355_;
  assign new_n19354_ = ~\all_features[2208]  & ~\all_features[2209] ;
  assign new_n19355_ = ~\all_features[2210]  & ~\all_features[2211] ;
  assign new_n19356_ = \all_features[2215]  & \all_features[2214]  & ~new_n19357_ & \all_features[2213] ;
  assign new_n19357_ = ~\all_features[2211]  & ~\all_features[2212]  & (~\all_features[2210]  | new_n19354_);
  assign new_n19358_ = \all_features[2215]  & \all_features[2214]  & ~new_n19361_ & new_n19359_;
  assign new_n19359_ = \all_features[2215]  & (\all_features[2214]  | (new_n19360_ & (\all_features[2210]  | \all_features[2211]  | \all_features[2209] )));
  assign new_n19360_ = \all_features[2212]  & \all_features[2213] ;
  assign new_n19361_ = new_n19355_ & ~\all_features[2213]  & ~new_n19362_ & ~\all_features[2212] ;
  assign new_n19362_ = \all_features[2208]  & \all_features[2209] ;
  assign new_n19363_ = ~new_n19364_ & ~new_n19366_;
  assign new_n19364_ = ~new_n19365_ & ~\all_features[2215] ;
  assign new_n19365_ = \all_features[2213]  & \all_features[2214]  & (\all_features[2212]  | (\all_features[2210]  & \all_features[2211]  & \all_features[2209] ));
  assign new_n19366_ = ~\all_features[2215]  & (~\all_features[2214]  | ~new_n19360_ | ~new_n19362_ | ~new_n19367_);
  assign new_n19367_ = \all_features[2210]  & \all_features[2211] ;
  assign new_n19368_ = ~\all_features[2215]  & (~\all_features[2214]  | (~\all_features[2212]  & ~\all_features[2213]  & ~new_n19367_));
  assign new_n19369_ = ~\all_features[2215]  & (~\all_features[2214]  | (~\all_features[2213]  & (new_n19354_ | ~new_n19367_ | ~\all_features[2212] )));
  assign new_n19370_ = new_n19363_ & new_n19371_ & ~new_n19376_ & ~new_n19375_ & ~new_n19368_ & ~new_n19369_;
  assign new_n19371_ = ~new_n19372_ & ~new_n19374_;
  assign new_n19372_ = ~\all_features[2213]  & new_n19373_ & ((~\all_features[2210]  & new_n19354_) | ~\all_features[2212]  | ~\all_features[2211] );
  assign new_n19373_ = ~\all_features[2214]  & ~\all_features[2215] ;
  assign new_n19374_ = ~\all_features[2215]  & ~\all_features[2214]  & ~\all_features[2213]  & ~\all_features[2211]  & ~\all_features[2212] ;
  assign new_n19375_ = new_n19373_ & (~\all_features[2211]  | ~new_n19360_ | (~new_n19362_ & ~\all_features[2210] ));
  assign new_n19376_ = new_n19373_ & (~\all_features[2213]  | (~\all_features[2212]  & (~\all_features[2211]  | (~\all_features[2210]  & ~\all_features[2209] ))));
  assign new_n19377_ = ~new_n19364_ & ~new_n19366_ & ~new_n19368_ & ~new_n19369_ & (~new_n19358_ | ~new_n19352_);
  assign new_n19378_ = ~new_n19342_ & new_n13522_;
  assign new_n19379_ = new_n19380_ & new_n19381_;
  assign new_n19380_ = ~new_n15172_ & ~new_n15195_;
  assign new_n19381_ = ~new_n15198_ & ~new_n15202_;
  assign new_n19382_ = new_n19414_ & new_n19383_ & new_n19412_;
  assign new_n19383_ = new_n19384_ & new_n19405_;
  assign new_n19384_ = ~new_n19385_ & (\all_features[2851]  | \all_features[2852]  | \all_features[2853]  | \all_features[2854]  | \all_features[2855] );
  assign new_n19385_ = ~new_n19399_ & (new_n19401_ | (~new_n19402_ & (new_n19403_ | (~new_n19386_ & ~new_n19404_))));
  assign new_n19386_ = ~new_n19387_ & (new_n19389_ | (new_n19398_ & (~new_n19393_ | (~new_n19397_ & new_n19396_))));
  assign new_n19387_ = ~new_n19388_ & ~\all_features[2855] ;
  assign new_n19388_ = \all_features[2853]  & \all_features[2854]  & (\all_features[2852]  | (\all_features[2850]  & \all_features[2851]  & \all_features[2849] ));
  assign new_n19389_ = ~\all_features[2855]  & (~\all_features[2854]  | ~new_n19390_ | ~new_n19391_ | ~new_n19392_);
  assign new_n19390_ = \all_features[2848]  & \all_features[2849] ;
  assign new_n19391_ = \all_features[2852]  & \all_features[2853] ;
  assign new_n19392_ = \all_features[2850]  & \all_features[2851] ;
  assign new_n19393_ = \all_features[2855]  & (\all_features[2854]  | (\all_features[2853]  & (\all_features[2852]  | ~new_n19395_ | ~new_n19394_)));
  assign new_n19394_ = ~\all_features[2848]  & ~\all_features[2849] ;
  assign new_n19395_ = ~\all_features[2850]  & ~\all_features[2851] ;
  assign new_n19396_ = \all_features[2855]  & (\all_features[2854]  | (new_n19391_ & (\all_features[2850]  | \all_features[2851]  | \all_features[2849] )));
  assign new_n19397_ = ~\all_features[2853]  & \all_features[2854]  & \all_features[2855]  & (\all_features[2852]  ? new_n19395_ : (new_n19390_ | ~new_n19395_));
  assign new_n19398_ = \all_features[2855]  & (\all_features[2853]  | \all_features[2854]  | \all_features[2852] );
  assign new_n19399_ = ~\all_features[2853]  & new_n19400_ & ((~\all_features[2850]  & new_n19394_) | ~\all_features[2852]  | ~\all_features[2851] );
  assign new_n19400_ = ~\all_features[2854]  & ~\all_features[2855] ;
  assign new_n19401_ = new_n19400_ & (~\all_features[2853]  | (~\all_features[2852]  & (~\all_features[2851]  | (~\all_features[2850]  & ~\all_features[2849] ))));
  assign new_n19402_ = new_n19400_ & (~\all_features[2851]  | ~new_n19391_ | (~\all_features[2850]  & ~new_n19390_));
  assign new_n19403_ = ~\all_features[2855]  & (~\all_features[2854]  | (~\all_features[2852]  & ~\all_features[2853]  & ~new_n19392_));
  assign new_n19404_ = ~\all_features[2855]  & (~\all_features[2854]  | (~\all_features[2853]  & (new_n19394_ | ~new_n19392_ | ~\all_features[2852] )));
  assign new_n19405_ = new_n19410_ & (~new_n19411_ | (~new_n19406_ & ~new_n19403_ & ~new_n19404_));
  assign new_n19406_ = ~new_n19387_ & ~new_n19389_ & (~new_n19398_ | ~new_n19393_ | new_n19407_);
  assign new_n19407_ = new_n19396_ & new_n19408_ & (new_n19409_ | ~\all_features[2853]  | ~\all_features[2854]  | ~\all_features[2855] );
  assign new_n19408_ = \all_features[2854]  & \all_features[2855]  & (\all_features[2852]  | \all_features[2853]  | new_n19390_ | ~new_n19395_);
  assign new_n19409_ = ~\all_features[2851]  & ~\all_features[2852]  & (~\all_features[2850]  | new_n19394_);
  assign new_n19410_ = ~new_n19399_ & (\all_features[2851]  | \all_features[2852]  | \all_features[2853]  | \all_features[2854]  | \all_features[2855] );
  assign new_n19411_ = ~new_n19401_ & ~new_n19402_;
  assign new_n19412_ = new_n19413_ & new_n19410_ & ~new_n19387_ & ~new_n19404_ & ~new_n19401_ & ~new_n19402_;
  assign new_n19413_ = ~new_n19403_ & ~new_n19389_;
  assign new_n19414_ = new_n19410_ & new_n19411_ & (new_n19415_ | new_n19404_ | new_n19387_ | ~new_n19413_);
  assign new_n19415_ = new_n19398_ & new_n19408_ & new_n19393_ & new_n19396_;
  assign new_n19416_ = ~new_n19417_ & ((new_n19342_ & (~new_n19344_ | new_n19337_)) | (new_n19418_ & new_n13522_ & ~new_n19342_));
  assign new_n19417_ = new_n19347_ & ~new_n19348_ & ~new_n19350_;
  assign new_n19418_ = new_n19379_ ? ~new_n19382_ : ~new_n12849_;
  assign new_n19419_ = new_n19420_ & new_n19467_;
  assign new_n19420_ = new_n19421_ & ~new_n19424_ & (~new_n19423_ | ~new_n19425_ | new_n19433_ | new_n11096_);
  assign new_n19421_ = ~new_n19422_ & (~new_n15913_ | ~new_n11096_ | new_n16765_ | new_n8390_);
  assign new_n19422_ = new_n19197_ & new_n17454_ & ~new_n19423_ & ~new_n11096_;
  assign new_n19423_ = ~new_n9168_ & ~new_n7902_;
  assign new_n19424_ = ~new_n16765_ & ~new_n15913_ & new_n11096_ & (new_n11699_ | (~new_n13203_ & new_n11675_));
  assign new_n19425_ = new_n19426_ & new_n19432_;
  assign new_n19426_ = ~new_n19427_ & ~new_n16482_;
  assign new_n19427_ = (new_n19428_ | (new_n16466_ & (~\all_features[1459]  | ~\all_features[1460]  | (~\all_features[1458]  & new_n16465_)))) & (~new_n16466_ | \all_features[1459]  | \all_features[1460] );
  assign new_n19428_ = ~new_n16462_ & (new_n16459_ | (~new_n16473_ & (new_n16476_ | (~new_n19429_ & ~new_n16477_))));
  assign new_n19429_ = ~new_n16475_ & (~\all_features[1463]  | new_n19430_ | (~\all_features[1460]  & ~\all_features[1461]  & ~\all_features[1462] ));
  assign new_n19430_ = \all_features[1463]  & ((~new_n19431_ & ~\all_features[1461]  & \all_features[1462] ) | (~new_n16470_ & (\all_features[1462]  | (~new_n16468_ & \all_features[1461] ))));
  assign new_n19431_ = (\all_features[1460]  & (\all_features[1458]  | \all_features[1459] )) | (~new_n16460_ & ~\all_features[1458]  & ~\all_features[1459]  & ~\all_features[1460] );
  assign new_n19432_ = ~new_n16456_ & ~new_n16479_;
  assign new_n19433_ = new_n19434_ & ~new_n19459_ & ~new_n19463_;
  assign new_n19434_ = ~new_n19435_ & ~new_n19457_;
  assign new_n19435_ = new_n19452_ & ~new_n19456_ & ~new_n19436_ & ~new_n19455_;
  assign new_n19436_ = new_n19437_ & (~new_n19450_ | ~new_n19451_ | ~new_n19447_ | ~new_n19449_);
  assign new_n19437_ = ~new_n19444_ & ~new_n19442_ & ~new_n19438_ & ~new_n19440_;
  assign new_n19438_ = ~\all_features[1223]  & (~\all_features[1222]  | (~\all_features[1220]  & ~\all_features[1221]  & ~new_n19439_));
  assign new_n19439_ = \all_features[1218]  & \all_features[1219] ;
  assign new_n19440_ = ~\all_features[1223]  & (~\all_features[1222]  | (~\all_features[1221]  & (new_n19441_ | ~new_n19439_ | ~\all_features[1220] )));
  assign new_n19441_ = ~\all_features[1216]  & ~\all_features[1217] ;
  assign new_n19442_ = ~new_n19443_ & ~\all_features[1223] ;
  assign new_n19443_ = \all_features[1221]  & \all_features[1222]  & (\all_features[1220]  | (\all_features[1218]  & \all_features[1219]  & \all_features[1217] ));
  assign new_n19444_ = ~\all_features[1223]  & (~\all_features[1222]  | ~new_n19445_ | ~new_n19446_ | ~new_n19439_);
  assign new_n19445_ = \all_features[1216]  & \all_features[1217] ;
  assign new_n19446_ = \all_features[1220]  & \all_features[1221] ;
  assign new_n19447_ = \all_features[1223]  & (\all_features[1222]  | (\all_features[1221]  & (\all_features[1220]  | ~new_n19448_ | ~new_n19441_)));
  assign new_n19448_ = ~\all_features[1218]  & ~\all_features[1219] ;
  assign new_n19449_ = \all_features[1223]  & (\all_features[1222]  | (new_n19446_ & (\all_features[1218]  | \all_features[1219]  | \all_features[1217] )));
  assign new_n19450_ = \all_features[1222]  & \all_features[1223]  & (\all_features[1220]  | \all_features[1221]  | new_n19445_ | ~new_n19448_);
  assign new_n19451_ = \all_features[1223]  & (\all_features[1221]  | \all_features[1222]  | \all_features[1220] );
  assign new_n19452_ = ~new_n19453_ & (\all_features[1219]  | \all_features[1220]  | \all_features[1221]  | \all_features[1222]  | \all_features[1223] );
  assign new_n19453_ = ~\all_features[1221]  & new_n19454_ & ((~\all_features[1218]  & new_n19441_) | ~\all_features[1220]  | ~\all_features[1219] );
  assign new_n19454_ = ~\all_features[1222]  & ~\all_features[1223] ;
  assign new_n19455_ = new_n19454_ & (~\all_features[1221]  | (~\all_features[1220]  & (~\all_features[1219]  | (~\all_features[1218]  & ~\all_features[1217] ))));
  assign new_n19456_ = new_n19454_ & (~\all_features[1219]  | ~new_n19446_ | (~\all_features[1218]  & ~new_n19445_));
  assign new_n19457_ = new_n19458_ & new_n19452_ & ~new_n19455_ & ~new_n19442_;
  assign new_n19458_ = ~new_n19444_ & ~new_n19440_ & ~new_n19456_ & ~new_n19438_;
  assign new_n19459_ = ~new_n19460_ & (\all_features[1219]  | \all_features[1220]  | \all_features[1221]  | \all_features[1222]  | \all_features[1223] );
  assign new_n19460_ = ~new_n19453_ & (new_n19455_ | (~new_n19456_ & (new_n19438_ | (~new_n19461_ & ~new_n19440_))));
  assign new_n19461_ = ~new_n19442_ & (new_n19444_ | (new_n19451_ & (~new_n19447_ | (~new_n19462_ & new_n19449_))));
  assign new_n19462_ = ~\all_features[1221]  & \all_features[1222]  & \all_features[1223]  & (\all_features[1220]  ? new_n19448_ : (new_n19445_ | ~new_n19448_));
  assign new_n19463_ = new_n19452_ & (new_n19456_ | new_n19455_ | (~new_n19464_ & ~new_n19438_ & ~new_n19440_));
  assign new_n19464_ = ~new_n19442_ & ~new_n19444_ & (~new_n19451_ | ~new_n19447_ | new_n19465_);
  assign new_n19465_ = new_n19449_ & new_n19450_ & (new_n19466_ | ~\all_features[1221]  | ~\all_features[1222]  | ~\all_features[1223] );
  assign new_n19466_ = ~\all_features[1219]  & ~\all_features[1220]  & (~\all_features[1218]  | new_n19441_);
  assign new_n19467_ = (new_n19468_ | new_n11096_) & (~new_n16765_ | ~new_n11096_ | (new_n17898_ ? ~new_n19500_ : new_n19499_));
  assign new_n19468_ = (new_n19425_ | ~new_n12266_ | ~new_n19423_) & (new_n19197_ | new_n19469_ | new_n19423_);
  assign new_n19469_ = ~new_n19497_ & ~new_n19470_ & ~new_n19494_;
  assign new_n19470_ = new_n19485_ & (~new_n19490_ | (~new_n19488_ & ~new_n19471_ & ~new_n19493_));
  assign new_n19471_ = ~new_n19482_ & ~new_n19481_ & (~new_n19484_ | ~new_n19480_ | new_n19472_);
  assign new_n19472_ = new_n19473_ & new_n19477_ & (new_n19475_ | ~\all_features[2277]  | ~\all_features[2278]  | ~\all_features[2279] );
  assign new_n19473_ = \all_features[2279]  & (\all_features[2278]  | (new_n19474_ & (\all_features[2274]  | \all_features[2275]  | \all_features[2273] )));
  assign new_n19474_ = \all_features[2276]  & \all_features[2277] ;
  assign new_n19475_ = ~\all_features[2275]  & ~\all_features[2276]  & (~\all_features[2274]  | new_n19476_);
  assign new_n19476_ = ~\all_features[2272]  & ~\all_features[2273] ;
  assign new_n19477_ = \all_features[2278]  & \all_features[2279]  & (\all_features[2276]  | \all_features[2277]  | new_n19479_ | ~new_n19478_);
  assign new_n19478_ = ~\all_features[2274]  & ~\all_features[2275] ;
  assign new_n19479_ = \all_features[2272]  & \all_features[2273] ;
  assign new_n19480_ = \all_features[2279]  & (\all_features[2278]  | (\all_features[2277]  & (\all_features[2276]  | ~new_n19478_ | ~new_n19476_)));
  assign new_n19481_ = ~\all_features[2279]  & (~new_n19479_ | ~\all_features[2274]  | ~\all_features[2275]  | ~\all_features[2278]  | ~new_n19474_);
  assign new_n19482_ = ~new_n19483_ & ~\all_features[2279] ;
  assign new_n19483_ = \all_features[2277]  & \all_features[2278]  & (\all_features[2276]  | (\all_features[2274]  & \all_features[2275]  & \all_features[2273] ));
  assign new_n19484_ = \all_features[2279]  & (\all_features[2277]  | \all_features[2278]  | \all_features[2276] );
  assign new_n19485_ = ~new_n19486_ & (\all_features[2275]  | \all_features[2276]  | \all_features[2277]  | \all_features[2278]  | \all_features[2279] );
  assign new_n19486_ = ~\all_features[2277]  & new_n19487_ & ((~\all_features[2274]  & new_n19476_) | ~\all_features[2276]  | ~\all_features[2275] );
  assign new_n19487_ = ~\all_features[2278]  & ~\all_features[2279] ;
  assign new_n19488_ = ~\all_features[2279]  & (~\all_features[2278]  | new_n19489_);
  assign new_n19489_ = ~\all_features[2277]  & (new_n19476_ | ~\all_features[2275]  | ~\all_features[2276]  | ~\all_features[2274] );
  assign new_n19490_ = ~new_n19491_ & ~new_n19492_;
  assign new_n19491_ = new_n19487_ & (~\all_features[2275]  | ~new_n19474_ | (~new_n19479_ & ~\all_features[2274] ));
  assign new_n19492_ = new_n19487_ & (~\all_features[2277]  | (~\all_features[2276]  & (~\all_features[2275]  | (~\all_features[2274]  & ~\all_features[2273] ))));
  assign new_n19493_ = ~\all_features[2279]  & (~\all_features[2278]  | (~\all_features[2277]  & ~\all_features[2276]  & (~\all_features[2275]  | ~\all_features[2274] )));
  assign new_n19494_ = new_n19490_ & ~new_n19495_ & new_n19485_;
  assign new_n19495_ = ~new_n19493_ & ~new_n19482_ & ~new_n19481_ & ~new_n19488_ & ~new_n19496_;
  assign new_n19496_ = new_n19484_ & new_n19480_ & new_n19473_ & new_n19477_;
  assign new_n19497_ = new_n19485_ & new_n19498_ & ~new_n19482_ & ~new_n19492_;
  assign new_n19498_ = ~new_n19493_ & ~new_n19491_ & ~new_n19488_ & ~new_n19481_;
  assign new_n19499_ = ~new_n14985_ & (~new_n14955_ | new_n17892_);
  assign new_n19500_ = ~new_n17549_ & new_n19501_;
  assign new_n19501_ = ~new_n17553_ & ~new_n17521_ & ~new_n17544_;
  assign new_n19502_ = ~new_n19588_ & new_n19503_;
  assign new_n19503_ = ~new_n19504_ & (new_n12374_ | ~new_n19550_) & (~new_n19587_ | ~new_n19549_);
  assign new_n19504_ = ~new_n19546_ & ((~new_n19505_ & new_n19544_) | (~new_n12117_ & new_n19548_ & ~new_n19544_));
  assign new_n19505_ = new_n19543_ ? new_n19508_ : new_n19506_;
  assign new_n19506_ = new_n9171_ & new_n19507_;
  assign new_n19507_ = ~new_n9204_ & ~new_n9207_;
  assign new_n19508_ = new_n19509_ & ~new_n19538_ & ~new_n19541_;
  assign new_n19509_ = ~new_n19510_ & ~new_n19534_;
  assign new_n19510_ = new_n19525_ & (~new_n19530_ | (~new_n19528_ & ~new_n19511_ & ~new_n19533_));
  assign new_n19511_ = ~new_n19523_ & ~new_n19521_ & (~new_n19524_ | ~new_n19520_ | new_n19512_);
  assign new_n19512_ = new_n19513_ & new_n19515_ & (new_n19518_ | ~\all_features[5301]  | ~\all_features[5302]  | ~\all_features[5303] );
  assign new_n19513_ = \all_features[5303]  & (\all_features[5302]  | (new_n19514_ & (\all_features[5298]  | \all_features[5299]  | \all_features[5297] )));
  assign new_n19514_ = \all_features[5300]  & \all_features[5301] ;
  assign new_n19515_ = \all_features[5302]  & \all_features[5303]  & (\all_features[5300]  | \all_features[5301]  | new_n19517_ | ~new_n19516_);
  assign new_n19516_ = ~\all_features[5298]  & ~\all_features[5299] ;
  assign new_n19517_ = \all_features[5296]  & \all_features[5297] ;
  assign new_n19518_ = ~\all_features[5299]  & ~\all_features[5300]  & (~\all_features[5298]  | new_n19519_);
  assign new_n19519_ = ~\all_features[5296]  & ~\all_features[5297] ;
  assign new_n19520_ = \all_features[5303]  & (\all_features[5302]  | (\all_features[5301]  & (\all_features[5300]  | ~new_n19516_ | ~new_n19519_)));
  assign new_n19521_ = ~new_n19522_ & ~\all_features[5303] ;
  assign new_n19522_ = \all_features[5301]  & \all_features[5302]  & (\all_features[5300]  | (\all_features[5298]  & \all_features[5299]  & \all_features[5297] ));
  assign new_n19523_ = ~\all_features[5303]  & (~new_n19517_ | ~\all_features[5298]  | ~\all_features[5299]  | ~\all_features[5302]  | ~new_n19514_);
  assign new_n19524_ = \all_features[5303]  & (\all_features[5301]  | \all_features[5302]  | \all_features[5300] );
  assign new_n19525_ = ~new_n19526_ & (\all_features[5299]  | \all_features[5300]  | \all_features[5301]  | \all_features[5302]  | \all_features[5303] );
  assign new_n19526_ = ~\all_features[5301]  & new_n19527_ & ((~\all_features[5298]  & new_n19519_) | ~\all_features[5300]  | ~\all_features[5299] );
  assign new_n19527_ = ~\all_features[5302]  & ~\all_features[5303] ;
  assign new_n19528_ = ~\all_features[5303]  & (~\all_features[5302]  | new_n19529_);
  assign new_n19529_ = ~\all_features[5301]  & (new_n19519_ | ~\all_features[5299]  | ~\all_features[5300]  | ~\all_features[5298] );
  assign new_n19530_ = ~new_n19531_ & ~new_n19532_;
  assign new_n19531_ = new_n19527_ & (~\all_features[5299]  | ~new_n19514_ | (~new_n19517_ & ~\all_features[5298] ));
  assign new_n19532_ = new_n19527_ & (~\all_features[5301]  | (~\all_features[5300]  & (~\all_features[5299]  | (~\all_features[5298]  & ~\all_features[5297] ))));
  assign new_n19533_ = ~\all_features[5303]  & (~\all_features[5302]  | (~\all_features[5301]  & ~\all_features[5300]  & (~\all_features[5299]  | ~\all_features[5298] )));
  assign new_n19534_ = ~new_n19535_ & (\all_features[5299]  | \all_features[5300]  | \all_features[5301]  | \all_features[5302]  | \all_features[5303] );
  assign new_n19535_ = ~new_n19526_ & (new_n19532_ | (~new_n19531_ & (new_n19533_ | (~new_n19528_ & ~new_n19536_))));
  assign new_n19536_ = ~new_n19521_ & (new_n19523_ | (new_n19524_ & (~new_n19520_ | (~new_n19537_ & new_n19513_))));
  assign new_n19537_ = ~\all_features[5301]  & \all_features[5302]  & \all_features[5303]  & (\all_features[5300]  ? new_n19516_ : (new_n19517_ | ~new_n19516_));
  assign new_n19538_ = new_n19530_ & ~new_n19539_ & new_n19525_;
  assign new_n19539_ = ~new_n19533_ & ~new_n19523_ & ~new_n19521_ & ~new_n19528_ & ~new_n19540_;
  assign new_n19540_ = new_n19524_ & new_n19520_ & new_n19513_ & new_n19515_;
  assign new_n19541_ = new_n19525_ & new_n19542_ & ~new_n19521_ & ~new_n19532_;
  assign new_n19542_ = ~new_n19533_ & ~new_n19531_ & ~new_n19528_ & ~new_n19523_;
  assign new_n19543_ = new_n18136_ & new_n18132_ & new_n18139_ & ~new_n18143_ & ~new_n18144_;
  assign new_n19544_ = new_n12446_ & new_n19545_;
  assign new_n19545_ = ~new_n8591_ & ~new_n8594_;
  assign new_n19546_ = new_n19547_ & ~new_n19281_ & ~new_n19305_;
  assign new_n19547_ = ~new_n19309_ & ~new_n19311_;
  assign new_n19548_ = new_n17521_ & new_n17553_;
  assign new_n19549_ = ~new_n19548_ & ~new_n19544_ & ~new_n19546_;
  assign new_n19550_ = new_n19546_ & ~new_n19551_ & ~new_n19586_;
  assign new_n19551_ = new_n19552_ & ~new_n19581_ & ~new_n19584_;
  assign new_n19552_ = ~new_n19553_ & ~new_n19577_;
  assign new_n19553_ = new_n19568_ & (~new_n19573_ | (~new_n19571_ & ~new_n19554_ & ~new_n19576_));
  assign new_n19554_ = ~new_n19566_ & ~new_n19564_ & (~new_n19567_ | ~new_n19563_ | new_n19555_);
  assign new_n19555_ = new_n19556_ & new_n19558_ & (new_n19561_ | ~\all_features[4213]  | ~\all_features[4214]  | ~\all_features[4215] );
  assign new_n19556_ = \all_features[4215]  & (\all_features[4214]  | (new_n19557_ & (\all_features[4210]  | \all_features[4211]  | \all_features[4209] )));
  assign new_n19557_ = \all_features[4212]  & \all_features[4213] ;
  assign new_n19558_ = \all_features[4214]  & \all_features[4215]  & (\all_features[4212]  | \all_features[4213]  | new_n19560_ | ~new_n19559_);
  assign new_n19559_ = ~\all_features[4210]  & ~\all_features[4211] ;
  assign new_n19560_ = \all_features[4208]  & \all_features[4209] ;
  assign new_n19561_ = ~\all_features[4211]  & ~\all_features[4212]  & (~\all_features[4210]  | new_n19562_);
  assign new_n19562_ = ~\all_features[4208]  & ~\all_features[4209] ;
  assign new_n19563_ = \all_features[4215]  & (\all_features[4214]  | (\all_features[4213]  & (\all_features[4212]  | ~new_n19559_ | ~new_n19562_)));
  assign new_n19564_ = ~new_n19565_ & ~\all_features[4215] ;
  assign new_n19565_ = \all_features[4213]  & \all_features[4214]  & (\all_features[4212]  | (\all_features[4210]  & \all_features[4211]  & \all_features[4209] ));
  assign new_n19566_ = ~\all_features[4215]  & (~new_n19560_ | ~\all_features[4210]  | ~\all_features[4211]  | ~\all_features[4214]  | ~new_n19557_);
  assign new_n19567_ = \all_features[4215]  & (\all_features[4213]  | \all_features[4214]  | \all_features[4212] );
  assign new_n19568_ = ~new_n19569_ & (\all_features[4211]  | \all_features[4212]  | \all_features[4213]  | \all_features[4214]  | \all_features[4215] );
  assign new_n19569_ = ~\all_features[4213]  & new_n19570_ & ((~\all_features[4210]  & new_n19562_) | ~\all_features[4212]  | ~\all_features[4211] );
  assign new_n19570_ = ~\all_features[4214]  & ~\all_features[4215] ;
  assign new_n19571_ = ~\all_features[4215]  & (~\all_features[4214]  | new_n19572_);
  assign new_n19572_ = ~\all_features[4213]  & (new_n19562_ | ~\all_features[4211]  | ~\all_features[4212]  | ~\all_features[4210] );
  assign new_n19573_ = ~new_n19574_ & ~new_n19575_;
  assign new_n19574_ = new_n19570_ & (~\all_features[4211]  | ~new_n19557_ | (~new_n19560_ & ~\all_features[4210] ));
  assign new_n19575_ = new_n19570_ & (~\all_features[4213]  | (~\all_features[4212]  & (~\all_features[4211]  | (~\all_features[4210]  & ~\all_features[4209] ))));
  assign new_n19576_ = ~\all_features[4215]  & (~\all_features[4214]  | (~\all_features[4213]  & ~\all_features[4212]  & (~\all_features[4211]  | ~\all_features[4210] )));
  assign new_n19577_ = ~new_n19578_ & (\all_features[4211]  | \all_features[4212]  | \all_features[4213]  | \all_features[4214]  | \all_features[4215] );
  assign new_n19578_ = ~new_n19569_ & (new_n19575_ | (~new_n19574_ & (new_n19576_ | (~new_n19571_ & ~new_n19579_))));
  assign new_n19579_ = ~new_n19564_ & (new_n19566_ | (new_n19567_ & (~new_n19563_ | (~new_n19580_ & new_n19556_))));
  assign new_n19580_ = ~\all_features[4213]  & \all_features[4214]  & \all_features[4215]  & (\all_features[4212]  ? new_n19559_ : (new_n19560_ | ~new_n19559_));
  assign new_n19581_ = new_n19573_ & ~new_n19582_ & new_n19568_;
  assign new_n19582_ = ~new_n19576_ & ~new_n19566_ & ~new_n19564_ & ~new_n19571_ & ~new_n19583_;
  assign new_n19583_ = new_n19567_ & new_n19563_ & new_n19556_ & new_n19558_;
  assign new_n19584_ = new_n19568_ & new_n19585_ & ~new_n19564_ & ~new_n19575_;
  assign new_n19585_ = ~new_n19576_ & ~new_n19574_ & ~new_n19571_ & ~new_n19566_;
  assign new_n19586_ = ~new_n11000_ & ~new_n11016_;
  assign new_n19587_ = ~new_n7363_ & (~new_n7341_ | new_n7366_);
  assign new_n19588_ = new_n19589_ & (~new_n12374_ | ~new_n19550_) & (~new_n19549_ | new_n19587_);
  assign new_n19589_ = ~new_n19546_ | ((new_n19590_ | ~new_n19551_) & (new_n17675_ | ~new_n19586_ | new_n19551_));
  assign new_n19590_ = ~new_n14374_ & (new_n18705_ | ~new_n19592_) & (~new_n19591_ | ~new_n14352_);
  assign new_n19591_ = new_n14380_ & new_n14376_;
  assign new_n19592_ = ~new_n18691_ & ~new_n18702_;
  assign new_n19593_ = ~new_n19594_ & new_n19728_;
  assign new_n19594_ = ~new_n19716_ & new_n19595_ & (~new_n19706_ | ~new_n19719_) & (~new_n19705_ | ~new_n19718_);
  assign new_n19595_ = (~new_n19596_ | new_n18121_) & (~new_n19636_ | (~new_n19703_ & ~new_n19648_));
  assign new_n19596_ = new_n19604_ & ~new_n19597_ & new_n19598_;
  assign new_n19597_ = ~new_n12115_ & (~new_n12112_ | new_n12083_);
  assign new_n19598_ = new_n19599_ & ~new_n14008_ & ~new_n19600_;
  assign new_n19599_ = ~new_n13983_ & ~new_n14006_;
  assign new_n19600_ = ~new_n19601_ & (\all_features[4627]  | \all_features[4628]  | \all_features[4629]  | \all_features[4630]  | \all_features[4631] );
  assign new_n19601_ = ~new_n14002_ & (new_n14004_ | (~new_n14005_ & (new_n13995_ | (~new_n13999_ & ~new_n19602_))));
  assign new_n19602_ = ~new_n13993_ & (new_n14000_ | (new_n13991_ & (~new_n13997_ | (~new_n19603_ & new_n13986_))));
  assign new_n19603_ = ~\all_features[4629]  & \all_features[4630]  & \all_features[4631]  & (\all_features[4628]  ? new_n13989_ : (new_n13990_ | ~new_n13989_));
  assign new_n19604_ = ~new_n19632_ & new_n19605_;
  assign new_n19605_ = ~new_n19606_ & ~new_n19630_;
  assign new_n19606_ = new_n19627_ & ~new_n19607_ & new_n19623_;
  assign new_n19607_ = ~new_n19622_ & ~new_n19620_ & ~new_n19619_ & ~new_n19608_ & ~new_n19611_;
  assign new_n19608_ = ~\all_features[5743]  & (~\all_features[5742]  | new_n19609_);
  assign new_n19609_ = ~\all_features[5741]  & (new_n19610_ | ~\all_features[5739]  | ~\all_features[5740]  | ~\all_features[5738] );
  assign new_n19610_ = ~\all_features[5736]  & ~\all_features[5737] ;
  assign new_n19611_ = new_n19618_ & new_n19617_ & new_n19612_ & new_n19614_;
  assign new_n19612_ = \all_features[5743]  & (\all_features[5742]  | (new_n19613_ & (\all_features[5738]  | \all_features[5739]  | \all_features[5737] )));
  assign new_n19613_ = \all_features[5740]  & \all_features[5741] ;
  assign new_n19614_ = \all_features[5742]  & \all_features[5743]  & (\all_features[5740]  | \all_features[5741]  | new_n19616_ | ~new_n19615_);
  assign new_n19615_ = ~\all_features[5738]  & ~\all_features[5739] ;
  assign new_n19616_ = \all_features[5736]  & \all_features[5737] ;
  assign new_n19617_ = \all_features[5743]  & (\all_features[5742]  | (\all_features[5741]  & (\all_features[5740]  | ~new_n19615_ | ~new_n19610_)));
  assign new_n19618_ = \all_features[5743]  & (\all_features[5741]  | \all_features[5742]  | \all_features[5740] );
  assign new_n19619_ = ~\all_features[5743]  & (~new_n19616_ | ~\all_features[5738]  | ~\all_features[5739]  | ~\all_features[5742]  | ~new_n19613_);
  assign new_n19620_ = ~new_n19621_ & ~\all_features[5743] ;
  assign new_n19621_ = \all_features[5741]  & \all_features[5742]  & (\all_features[5740]  | (\all_features[5738]  & \all_features[5739]  & \all_features[5737] ));
  assign new_n19622_ = ~\all_features[5743]  & (~\all_features[5742]  | (~\all_features[5741]  & ~\all_features[5740]  & (~\all_features[5739]  | ~\all_features[5738] )));
  assign new_n19623_ = ~new_n19624_ & ~new_n19626_;
  assign new_n19624_ = ~\all_features[5741]  & new_n19625_ & ((~\all_features[5738]  & new_n19610_) | ~\all_features[5740]  | ~\all_features[5739] );
  assign new_n19625_ = ~\all_features[5742]  & ~\all_features[5743] ;
  assign new_n19626_ = ~\all_features[5743]  & ~\all_features[5742]  & ~\all_features[5741]  & ~\all_features[5739]  & ~\all_features[5740] ;
  assign new_n19627_ = ~new_n19628_ & ~new_n19629_;
  assign new_n19628_ = new_n19625_ & (~\all_features[5739]  | ~new_n19613_ | (~new_n19616_ & ~\all_features[5738] ));
  assign new_n19629_ = new_n19625_ & (~\all_features[5741]  | (~\all_features[5740]  & (~\all_features[5739]  | (~\all_features[5738]  & ~\all_features[5737] ))));
  assign new_n19630_ = new_n19623_ & new_n19631_ & ~new_n19620_ & ~new_n19629_;
  assign new_n19631_ = ~new_n19622_ & ~new_n19628_ & ~new_n19608_ & ~new_n19619_;
  assign new_n19632_ = new_n19623_ & (~new_n19627_ | (~new_n19608_ & ~new_n19633_ & ~new_n19622_));
  assign new_n19633_ = ~new_n19620_ & ~new_n19619_ & (~new_n19618_ | ~new_n19617_ | new_n19634_);
  assign new_n19634_ = new_n19612_ & new_n19614_ & (new_n19635_ | ~\all_features[5741]  | ~\all_features[5742]  | ~\all_features[5743] );
  assign new_n19635_ = ~\all_features[5739]  & ~\all_features[5740]  & (~\all_features[5738]  | new_n19610_);
  assign new_n19636_ = ~new_n19637_ & new_n19597_;
  assign new_n19637_ = ~new_n17414_ & (~new_n17392_ | new_n19638_);
  assign new_n19638_ = ~new_n19639_ & ~new_n19644_;
  assign new_n19639_ = ~new_n17398_ & (new_n17395_ | (~new_n17399_ & (new_n17400_ | (~new_n19640_ & ~new_n17412_))));
  assign new_n19640_ = ~new_n17408_ & (new_n17410_ | (~new_n17413_ & (~new_n19643_ | new_n19641_)));
  assign new_n19641_ = \all_features[3887]  & ((~new_n19642_ & ~\all_features[3885]  & \all_features[3886] ) | (~new_n17405_ & (\all_features[3886]  | (~new_n17403_ & \all_features[3885] ))));
  assign new_n19642_ = (~\all_features[3882]  & ~\all_features[3883]  & ~\all_features[3884]  & (~\all_features[3881]  | ~\all_features[3880] )) | (\all_features[3884]  & (\all_features[3882]  | \all_features[3883] ));
  assign new_n19643_ = \all_features[3887]  & (\all_features[3885]  | \all_features[3886]  | \all_features[3884] );
  assign new_n19644_ = new_n17394_ & (new_n17400_ | new_n17399_ | (~new_n17408_ & ~new_n17412_ & ~new_n19645_));
  assign new_n19645_ = ~new_n17410_ & ~new_n17413_ & (~new_n17402_ | (~new_n19646_ & new_n17404_));
  assign new_n19646_ = \all_features[3887]  & \all_features[3886]  & ~new_n19647_ & \all_features[3885] ;
  assign new_n19647_ = ~\all_features[3883]  & ~\all_features[3884]  & (~\all_features[3882]  | new_n17396_);
  assign new_n19648_ = ~new_n19649_ & new_n19678_;
  assign new_n19649_ = new_n19650_ & new_n19677_;
  assign new_n19650_ = new_n19651_ & new_n19673_;
  assign new_n19651_ = new_n19652_ & (~new_n19661_ | (new_n19671_ & new_n19672_ & new_n19668_ & new_n19670_));
  assign new_n19652_ = new_n19653_ & ~new_n19657_ & ~new_n19658_;
  assign new_n19653_ = ~new_n19654_ & (\all_features[2115]  | \all_features[2116]  | \all_features[2117]  | \all_features[2118]  | \all_features[2119] );
  assign new_n19654_ = ~\all_features[2117]  & new_n19656_ & ((~\all_features[2114]  & new_n19655_) | ~\all_features[2116]  | ~\all_features[2115] );
  assign new_n19655_ = ~\all_features[2112]  & ~\all_features[2113] ;
  assign new_n19656_ = ~\all_features[2118]  & ~\all_features[2119] ;
  assign new_n19657_ = new_n19656_ & (~\all_features[2117]  | (~\all_features[2116]  & (~\all_features[2115]  | (~\all_features[2114]  & ~\all_features[2113] ))));
  assign new_n19658_ = new_n19656_ & (~\all_features[2115]  | ~new_n19659_ | (~\all_features[2114]  & ~new_n19660_));
  assign new_n19659_ = \all_features[2116]  & \all_features[2117] ;
  assign new_n19660_ = \all_features[2112]  & \all_features[2113] ;
  assign new_n19661_ = ~new_n19667_ & ~new_n19666_ & ~new_n19662_ & ~new_n19664_;
  assign new_n19662_ = ~\all_features[2119]  & (~\all_features[2118]  | (~\all_features[2117]  & (new_n19655_ | ~new_n19663_ | ~\all_features[2116] )));
  assign new_n19663_ = \all_features[2114]  & \all_features[2115] ;
  assign new_n19664_ = ~new_n19665_ & ~\all_features[2119] ;
  assign new_n19665_ = \all_features[2117]  & \all_features[2118]  & (\all_features[2116]  | (\all_features[2114]  & \all_features[2115]  & \all_features[2113] ));
  assign new_n19666_ = ~\all_features[2119]  & (~\all_features[2118]  | ~new_n19659_ | ~new_n19660_ | ~new_n19663_);
  assign new_n19667_ = ~\all_features[2119]  & (~\all_features[2118]  | (~\all_features[2116]  & ~\all_features[2117]  & ~new_n19663_));
  assign new_n19668_ = \all_features[2119]  & (\all_features[2118]  | (\all_features[2117]  & (\all_features[2116]  | ~new_n19655_ | ~new_n19669_)));
  assign new_n19669_ = ~\all_features[2114]  & ~\all_features[2115] ;
  assign new_n19670_ = \all_features[2119]  & (\all_features[2118]  | (new_n19659_ & (\all_features[2114]  | \all_features[2115]  | \all_features[2113] )));
  assign new_n19671_ = \all_features[2118]  & \all_features[2119]  & (\all_features[2116]  | \all_features[2117]  | new_n19660_ | ~new_n19669_);
  assign new_n19672_ = \all_features[2119]  & (\all_features[2117]  | \all_features[2118]  | \all_features[2116] );
  assign new_n19673_ = new_n19653_ & (new_n19658_ | new_n19657_ | (~new_n19662_ & ~new_n19667_ & ~new_n19674_));
  assign new_n19674_ = ~new_n19666_ & ~new_n19664_ & (~new_n19672_ | ~new_n19668_ | new_n19675_);
  assign new_n19675_ = new_n19670_ & new_n19671_ & (new_n19676_ | ~\all_features[2117]  | ~\all_features[2118]  | ~\all_features[2119] );
  assign new_n19676_ = ~\all_features[2115]  & ~\all_features[2116]  & (~\all_features[2114]  | new_n19655_);
  assign new_n19677_ = new_n19652_ & new_n19661_;
  assign new_n19678_ = ~new_n19679_ & ~new_n19702_;
  assign new_n19679_ = new_n19680_ & (~new_n19691_ | (new_n19699_ & new_n19701_ & new_n19689_ & new_n19698_));
  assign new_n19680_ = new_n19681_ & ~new_n19686_ & ~new_n19687_;
  assign new_n19681_ = ~new_n19682_ & ~new_n19685_;
  assign new_n19682_ = ~\all_features[2749]  & new_n19684_ & ((~\all_features[2746]  & new_n19683_) | ~\all_features[2748]  | ~\all_features[2747] );
  assign new_n19683_ = ~\all_features[2744]  & ~\all_features[2745] ;
  assign new_n19684_ = ~\all_features[2750]  & ~\all_features[2751] ;
  assign new_n19685_ = ~\all_features[2751]  & ~\all_features[2750]  & ~\all_features[2749]  & ~\all_features[2747]  & ~\all_features[2748] ;
  assign new_n19686_ = new_n19684_ & (~\all_features[2749]  | (~\all_features[2748]  & (~\all_features[2747]  | (~\all_features[2746]  & ~\all_features[2745] ))));
  assign new_n19687_ = new_n19684_ & (~new_n19688_ | ~\all_features[2747]  | (~\all_features[2746]  & (~\all_features[2744]  | ~\all_features[2745] )));
  assign new_n19688_ = \all_features[2748]  & \all_features[2749] ;
  assign new_n19689_ = \all_features[2751]  & (\all_features[2750]  | new_n19690_);
  assign new_n19690_ = \all_features[2749]  & (\all_features[2746]  | \all_features[2747]  | \all_features[2748]  | ~new_n19683_);
  assign new_n19691_ = ~new_n19697_ & ~new_n19696_ & ~new_n19692_ & ~new_n19694_;
  assign new_n19692_ = ~\all_features[2751]  & (~\all_features[2750]  | (~\all_features[2749]  & (new_n19683_ | ~new_n19693_ | ~\all_features[2748] )));
  assign new_n19693_ = \all_features[2746]  & \all_features[2747] ;
  assign new_n19694_ = ~new_n19695_ & ~\all_features[2751] ;
  assign new_n19695_ = \all_features[2749]  & \all_features[2750]  & (\all_features[2748]  | (\all_features[2746]  & \all_features[2747]  & \all_features[2745] ));
  assign new_n19696_ = ~\all_features[2751]  & (~new_n19693_ | ~\all_features[2744]  | ~\all_features[2745]  | ~\all_features[2750]  | ~new_n19688_);
  assign new_n19697_ = ~\all_features[2751]  & (~\all_features[2750]  | (~\all_features[2748]  & ~\all_features[2749]  & ~new_n19693_));
  assign new_n19698_ = \all_features[2751]  & (\all_features[2750]  | (new_n19688_ & (\all_features[2746]  | \all_features[2747]  | \all_features[2745] )));
  assign new_n19699_ = \all_features[2751]  & ~new_n19700_ & \all_features[2750] ;
  assign new_n19700_ = ~\all_features[2746]  & ~\all_features[2747]  & ~\all_features[2748]  & ~\all_features[2749]  & (~\all_features[2745]  | ~\all_features[2744] );
  assign new_n19701_ = \all_features[2751]  & (\all_features[2749]  | \all_features[2750]  | \all_features[2748] );
  assign new_n19702_ = new_n19680_ & new_n19691_;
  assign new_n19703_ = new_n8188_ & ~new_n19678_ & new_n19704_;
  assign new_n19704_ = new_n8166_ & new_n8192_;
  assign new_n19705_ = new_n6847_ ? new_n16957_ : (new_n12490_ | (new_n12487_ & new_n12454_));
  assign new_n19706_ = ~new_n19707_ & ~new_n19597_ & ~new_n19598_;
  assign new_n19707_ = ~new_n18396_ & (~new_n18412_ | (~new_n19712_ & ~new_n19708_));
  assign new_n19708_ = new_n18397_ & (~new_n18419_ | (~new_n19709_ & ~new_n18410_ & ~new_n18406_));
  assign new_n19709_ = ~new_n18407_ & ~new_n18402_ & (~new_n18418_ | ~new_n18414_ | new_n19710_);
  assign new_n19710_ = new_n18416_ & new_n18417_ & (new_n19711_ | ~\all_features[2973]  | ~\all_features[2974]  | ~\all_features[2975] );
  assign new_n19711_ = ~\all_features[2971]  & ~\all_features[2972]  & (~\all_features[2970]  | new_n18400_);
  assign new_n19712_ = ~new_n19713_ & (\all_features[2971]  | \all_features[2972]  | \all_features[2973]  | \all_features[2974]  | \all_features[2975] );
  assign new_n19713_ = ~new_n18398_ & (new_n18409_ | (~new_n18411_ & (new_n18406_ | (~new_n18410_ & ~new_n19714_))));
  assign new_n19714_ = ~new_n18407_ & (new_n18402_ | (new_n18418_ & (~new_n18414_ | (~new_n19715_ & new_n18416_))));
  assign new_n19715_ = ~\all_features[2973]  & \all_features[2974]  & \all_features[2975]  & (\all_features[2972]  ? new_n18415_ : (new_n18404_ | ~new_n18415_));
  assign new_n19716_ = ~new_n19597_ & ((new_n19707_ & ~new_n19598_) | (~new_n19604_ & ~new_n19717_ & new_n19598_));
  assign new_n19717_ = new_n17845_ & new_n18918_;
  assign new_n19718_ = new_n19597_ & new_n19637_;
  assign new_n19719_ = new_n19678_ & new_n19720_;
  assign new_n19720_ = ~new_n19721_ & (new_n19685_ | (~new_n19725_ & ~new_n19682_));
  assign new_n19721_ = new_n19681_ & (new_n19687_ | new_n19686_ | (~new_n19692_ & ~new_n19697_ & ~new_n19722_));
  assign new_n19722_ = ~new_n19696_ & ~new_n19694_ & (~new_n19701_ | new_n19723_ | ~new_n19689_);
  assign new_n19723_ = ~new_n19700_ & new_n19698_ & \all_features[2750]  & \all_features[2751]  & (~\all_features[2749]  | new_n19724_);
  assign new_n19724_ = ~\all_features[2747]  & ~\all_features[2748]  & (~\all_features[2746]  | new_n19683_);
  assign new_n19725_ = ~new_n19686_ & (new_n19687_ | (~new_n19697_ & (new_n19692_ | (~new_n19694_ & ~new_n19726_))));
  assign new_n19726_ = ~new_n19696_ & (~new_n19701_ | (new_n19689_ & (~new_n19698_ | (~new_n19727_ & new_n19699_))));
  assign new_n19727_ = \all_features[2750]  & \all_features[2751]  & (\all_features[2749]  | (\all_features[2748]  & (\all_features[2747]  | \all_features[2746] )));
  assign new_n19728_ = new_n19729_ & (new_n19719_ | ~new_n19706_) & (~new_n19718_ | new_n19705_);
  assign new_n19729_ = (~new_n18121_ | ~new_n19596_) & (new_n19648_ | new_n19703_ | ~new_n19636_);
  assign new_n19730_ = new_n19731_ & (~new_n19775_ | (~new_n19815_ & new_n19814_));
  assign new_n19731_ = new_n19732_ & (~new_n19772_ | (new_n19055_ & new_n6701_) | (new_n19773_ & ~new_n6701_));
  assign new_n19732_ = ~new_n19734_ & (~new_n19769_ | ~new_n19770_ | ~new_n19771_) & (~new_n19733_ | ~new_n19768_);
  assign new_n19733_ = new_n18669_ & new_n18044_;
  assign new_n19734_ = new_n19735_ & (new_n17554_ ? ~new_n12727_ : new_n19767_);
  assign new_n19735_ = ~new_n19736_ & ~new_n19546_;
  assign new_n19736_ = ~new_n19766_ & new_n19737_;
  assign new_n19737_ = ~new_n19738_ & ~new_n19764_;
  assign new_n19738_ = new_n19758_ & (~new_n19754_ | (new_n19750_ & (new_n19739_ | new_n19761_ | new_n19763_)));
  assign new_n19739_ = new_n19740_ & (~new_n19744_ | (~new_n19749_ & \all_features[4357]  & \all_features[4358]  & \all_features[4359] ));
  assign new_n19740_ = \all_features[4359]  & (\all_features[4358]  | (~new_n19741_ & \all_features[4357] ));
  assign new_n19741_ = new_n19742_ & ~\all_features[4356]  & new_n19743_;
  assign new_n19742_ = ~\all_features[4352]  & ~\all_features[4353] ;
  assign new_n19743_ = ~\all_features[4354]  & ~\all_features[4355] ;
  assign new_n19744_ = \all_features[4359]  & \all_features[4358]  & ~new_n19747_ & new_n19745_;
  assign new_n19745_ = \all_features[4359]  & (\all_features[4358]  | (new_n19746_ & (\all_features[4354]  | \all_features[4355]  | \all_features[4353] )));
  assign new_n19746_ = \all_features[4356]  & \all_features[4357] ;
  assign new_n19747_ = new_n19743_ & ~\all_features[4357]  & ~new_n19748_ & ~\all_features[4356] ;
  assign new_n19748_ = \all_features[4352]  & \all_features[4353] ;
  assign new_n19749_ = ~\all_features[4355]  & ~\all_features[4356]  & (~\all_features[4354]  | new_n19742_);
  assign new_n19750_ = ~new_n19751_ & ~new_n19753_;
  assign new_n19751_ = ~\all_features[4359]  & (~\all_features[4358]  | (~\all_features[4356]  & ~\all_features[4357]  & ~new_n19752_));
  assign new_n19752_ = \all_features[4354]  & \all_features[4355] ;
  assign new_n19753_ = ~\all_features[4359]  & (~\all_features[4358]  | (~\all_features[4357]  & (new_n19742_ | ~\all_features[4356]  | ~new_n19752_)));
  assign new_n19754_ = ~new_n19755_ & ~new_n19757_;
  assign new_n19755_ = new_n19756_ & (~\all_features[4355]  | ~new_n19746_ | (~\all_features[4354]  & ~new_n19748_));
  assign new_n19756_ = ~\all_features[4358]  & ~\all_features[4359] ;
  assign new_n19757_ = new_n19756_ & (~\all_features[4357]  | (~\all_features[4356]  & (~\all_features[4355]  | (~\all_features[4354]  & ~\all_features[4353] ))));
  assign new_n19758_ = ~new_n19759_ & ~new_n19760_;
  assign new_n19759_ = ~\all_features[4357]  & new_n19756_ & ((~\all_features[4354]  & new_n19742_) | ~\all_features[4356]  | ~\all_features[4355] );
  assign new_n19760_ = ~\all_features[4359]  & ~\all_features[4358]  & ~\all_features[4357]  & ~\all_features[4355]  & ~\all_features[4356] ;
  assign new_n19761_ = ~new_n19762_ & ~\all_features[4359] ;
  assign new_n19762_ = \all_features[4357]  & \all_features[4358]  & (\all_features[4356]  | (\all_features[4354]  & \all_features[4355]  & \all_features[4353] ));
  assign new_n19763_ = ~\all_features[4359]  & (~\all_features[4358]  | ~new_n19752_ | ~new_n19748_ | ~new_n19746_);
  assign new_n19764_ = new_n19758_ & ~new_n19765_ & new_n19754_;
  assign new_n19765_ = ~new_n19751_ & ~new_n19753_ & ~new_n19761_ & ~new_n19763_ & (~new_n19744_ | ~new_n19740_);
  assign new_n19766_ = new_n19754_ & new_n19750_ & new_n19758_ & ~new_n19761_ & ~new_n19763_;
  assign new_n19767_ = ~new_n13882_ & ~new_n13880_ & ~new_n13851_ & ~new_n13873_;
  assign new_n19768_ = ~new_n19736_ & new_n19546_;
  assign new_n19769_ = new_n18580_ & new_n19736_;
  assign new_n19770_ = ~new_n9058_ & ~new_n9045_ & ~new_n9055_;
  assign new_n19771_ = ~\all_features[3119]  & ~\all_features[3118]  & ~\all_features[3117]  & ~\all_features[3115]  & ~\all_features[3116] ;
  assign new_n19772_ = ~new_n18580_ & new_n19736_;
  assign new_n19773_ = new_n14786_ & new_n19774_;
  assign new_n19774_ = new_n18082_ & new_n18086_;
  assign new_n19775_ = ~new_n19779_ & new_n19776_ & (~new_n19768_ | new_n19780_ | new_n19733_);
  assign new_n19776_ = ~new_n19777_ & (new_n17554_ | new_n19767_ | ~new_n19735_);
  assign new_n19777_ = new_n19769_ & ((~new_n19770_ & new_n19771_) | (~new_n19778_ & ~new_n13196_ & ~new_n19771_));
  assign new_n19778_ = new_n13197_ & new_n13170_;
  assign new_n19779_ = new_n19772_ & (new_n6701_ ? new_n19055_ : new_n19773_);
  assign new_n19780_ = ~new_n18669_ & new_n19781_;
  assign new_n19781_ = new_n19813_ & new_n19811_ & new_n19782_ & new_n19802_;
  assign new_n19782_ = ~new_n19801_ & (new_n19796_ | (~new_n19798_ & (new_n19799_ | (~new_n19783_ & ~new_n19800_))));
  assign new_n19783_ = ~new_n19790_ & (new_n19792_ | (~new_n19794_ & (~new_n19795_ | new_n19784_)));
  assign new_n19784_ = \all_features[4807]  & ((~new_n19789_ & ~\all_features[4805]  & \all_features[4806] ) | (~new_n19787_ & (\all_features[4806]  | (~new_n19785_ & \all_features[4805] ))));
  assign new_n19785_ = new_n19786_ & ~\all_features[4804]  & ~\all_features[4802]  & ~\all_features[4803] ;
  assign new_n19786_ = ~\all_features[4800]  & ~\all_features[4801] ;
  assign new_n19787_ = \all_features[4807]  & (\all_features[4806]  | (new_n19788_ & (\all_features[4802]  | \all_features[4803]  | \all_features[4801] )));
  assign new_n19788_ = \all_features[4804]  & \all_features[4805] ;
  assign new_n19789_ = (~\all_features[4802]  & ~\all_features[4803]  & ~\all_features[4804]  & (~\all_features[4801]  | ~\all_features[4800] )) | (\all_features[4804]  & (\all_features[4802]  | \all_features[4803] ));
  assign new_n19790_ = ~\all_features[4807]  & (~\all_features[4806]  | (~\all_features[4805]  & (new_n19786_ | ~new_n19791_ | ~\all_features[4804] )));
  assign new_n19791_ = \all_features[4802]  & \all_features[4803] ;
  assign new_n19792_ = ~new_n19793_ & ~\all_features[4807] ;
  assign new_n19793_ = \all_features[4805]  & \all_features[4806]  & (\all_features[4804]  | (\all_features[4802]  & \all_features[4803]  & \all_features[4801] ));
  assign new_n19794_ = ~\all_features[4807]  & (~new_n19791_ | ~\all_features[4800]  | ~\all_features[4801]  | ~\all_features[4806]  | ~new_n19788_);
  assign new_n19795_ = \all_features[4807]  & (\all_features[4805]  | \all_features[4806]  | \all_features[4804] );
  assign new_n19796_ = ~\all_features[4805]  & new_n19797_ & ((~\all_features[4802]  & new_n19786_) | ~\all_features[4804]  | ~\all_features[4803] );
  assign new_n19797_ = ~\all_features[4806]  & ~\all_features[4807] ;
  assign new_n19798_ = new_n19797_ & (~\all_features[4805]  | (~\all_features[4804]  & (~\all_features[4803]  | (~\all_features[4802]  & ~\all_features[4801] ))));
  assign new_n19799_ = new_n19797_ & (~new_n19788_ | ~\all_features[4803]  | (~\all_features[4802]  & (~\all_features[4800]  | ~\all_features[4801] )));
  assign new_n19800_ = ~\all_features[4807]  & (~\all_features[4806]  | (~\all_features[4804]  & ~\all_features[4805]  & ~new_n19791_));
  assign new_n19801_ = ~\all_features[4807]  & ~\all_features[4806]  & ~\all_features[4805]  & ~\all_features[4803]  & ~\all_features[4804] ;
  assign new_n19802_ = new_n19808_ & (~new_n19809_ | (new_n19810_ & (new_n19803_ | new_n19792_ | new_n19794_)));
  assign new_n19803_ = new_n19804_ & (~new_n19805_ | (~new_n19807_ & \all_features[4805]  & \all_features[4806]  & \all_features[4807] ));
  assign new_n19804_ = \all_features[4807]  & (\all_features[4806]  | (~new_n19785_ & \all_features[4805] ));
  assign new_n19805_ = \all_features[4807]  & \all_features[4806]  & ~new_n19806_ & new_n19787_;
  assign new_n19806_ = ~\all_features[4802]  & ~\all_features[4803]  & ~\all_features[4804]  & ~\all_features[4805]  & (~\all_features[4801]  | ~\all_features[4800] );
  assign new_n19807_ = ~\all_features[4803]  & ~\all_features[4804]  & (~\all_features[4802]  | new_n19786_);
  assign new_n19808_ = ~new_n19796_ & ~new_n19801_;
  assign new_n19809_ = ~new_n19798_ & ~new_n19799_;
  assign new_n19810_ = ~new_n19800_ & ~new_n19790_;
  assign new_n19811_ = new_n19809_ & ~new_n19812_ & new_n19808_;
  assign new_n19812_ = ~new_n19800_ & ~new_n19790_ & ~new_n19792_ & ~new_n19794_ & (~new_n19805_ | ~new_n19804_);
  assign new_n19813_ = new_n19810_ & new_n19809_ & ~new_n19801_ & ~new_n19794_ & ~new_n19796_ & ~new_n19792_;
  assign new_n19814_ = new_n19780_ & new_n19768_;
  assign new_n19815_ = new_n17554_ & new_n19735_ & new_n12727_;
  assign new_n19816_ = new_n19817_ & (~new_n19847_ | (new_n19877_ & new_n19878_));
  assign new_n19817_ = new_n19818_ & (~new_n19838_ | new_n19846_) & (~new_n19841_ | (~new_n19842_ & ~new_n19845_));
  assign new_n19818_ = (~new_n19837_ | ~new_n19819_) & (new_n19834_ | new_n19830_ | ~new_n19833_);
  assign new_n19819_ = ~new_n19828_ & new_n19820_;
  assign new_n19820_ = ~new_n19821_ & ~new_n19827_;
  assign new_n19821_ = new_n10408_ & new_n19822_;
  assign new_n19822_ = ~new_n10434_ & ~new_n19823_;
  assign new_n19823_ = ~new_n19824_ & (\all_features[2779]  | \all_features[2780]  | \all_features[2781]  | \all_features[2782]  | \all_features[2783] );
  assign new_n19824_ = ~new_n10427_ & (new_n10431_ | (~new_n10430_ & (new_n10425_ | (~new_n10411_ & ~new_n19825_))));
  assign new_n19825_ = ~new_n10423_ & (new_n10422_ | (new_n10421_ & (~new_n10420_ | (~new_n19826_ & new_n10415_))));
  assign new_n19826_ = ~\all_features[2781]  & \all_features[2782]  & \all_features[2783]  & (\all_features[2780]  ? new_n10418_ : (new_n10419_ | ~new_n10418_));
  assign new_n19827_ = ~new_n18256_ & (~new_n18253_ | new_n18224_);
  assign new_n19828_ = new_n19829_ & new_n9271_;
  assign new_n19829_ = new_n9249_ & new_n9275_;
  assign new_n19830_ = new_n19831_ & ~new_n15860_ & new_n19832_;
  assign new_n19831_ = new_n16518_ & (new_n16515_ | ~new_n16486_);
  assign new_n19832_ = ~new_n15853_ & ~new_n15862_;
  assign new_n19833_ = new_n18911_ & new_n19821_;
  assign new_n19834_ = ~new_n19831_ & ~new_n19835_;
  assign new_n19835_ = ~new_n13210_ & new_n19836_;
  assign new_n19836_ = ~new_n13238_ & ~new_n13242_;
  assign new_n19837_ = new_n14394_ & new_n14416_;
  assign new_n19838_ = ~new_n19840_ & new_n19839_;
  assign new_n19839_ = ~new_n18911_ & new_n19821_;
  assign new_n19840_ = ~new_n19721_ & new_n19678_;
  assign new_n19841_ = ~new_n19821_ & new_n19827_;
  assign new_n19842_ = ~new_n8855_ & ~new_n19843_;
  assign new_n19843_ = new_n15957_ & new_n19844_;
  assign new_n19844_ = ~new_n15986_ & ~new_n15990_;
  assign new_n19845_ = new_n8855_ & (~new_n17210_ | ~new_n17206_);
  assign new_n19846_ = ~new_n13160_ & new_n13135_;
  assign new_n19847_ = ~new_n19849_ & new_n19848_ & (~new_n19833_ | ~new_n19834_) & (new_n6497_ | ~new_n19876_);
  assign new_n19848_ = (~new_n19846_ | ~new_n19838_) & (new_n19842_ | new_n19845_ | ~new_n19841_);
  assign new_n19849_ = new_n19820_ & new_n19828_ & ~new_n19874_ & ~new_n19850_ & ~new_n19873_;
  assign new_n19850_ = new_n19865_ & (~new_n19867_ | (~new_n19851_ & new_n19870_));
  assign new_n19851_ = ~new_n19861_ & ~new_n19863_ & (~new_n19852_ | (~new_n19855_ & new_n19857_ & new_n19859_));
  assign new_n19852_ = \all_features[3759]  & (\all_features[3758]  | new_n19853_);
  assign new_n19853_ = \all_features[3757]  & (\all_features[3754]  | \all_features[3755]  | \all_features[3756]  | ~new_n19854_);
  assign new_n19854_ = ~\all_features[3752]  & ~\all_features[3753] ;
  assign new_n19855_ = \all_features[3759]  & \all_features[3758]  & ~new_n19856_ & \all_features[3757] ;
  assign new_n19856_ = ~\all_features[3755]  & ~\all_features[3756]  & (~\all_features[3754]  | new_n19854_);
  assign new_n19857_ = \all_features[3759]  & (\all_features[3758]  | (new_n19858_ & (\all_features[3754]  | \all_features[3755]  | \all_features[3753] )));
  assign new_n19858_ = \all_features[3756]  & \all_features[3757] ;
  assign new_n19859_ = \all_features[3759]  & ~new_n19860_ & \all_features[3758] ;
  assign new_n19860_ = ~\all_features[3754]  & ~\all_features[3755]  & ~\all_features[3756]  & ~\all_features[3757]  & (~\all_features[3753]  | ~\all_features[3752] );
  assign new_n19861_ = ~\all_features[3759]  & (~new_n19862_ | ~\all_features[3752]  | ~\all_features[3753]  | ~\all_features[3758]  | ~new_n19858_);
  assign new_n19862_ = \all_features[3754]  & \all_features[3755] ;
  assign new_n19863_ = ~new_n19864_ & ~\all_features[3759] ;
  assign new_n19864_ = \all_features[3757]  & \all_features[3758]  & (\all_features[3756]  | (\all_features[3754]  & \all_features[3755]  & \all_features[3753] ));
  assign new_n19865_ = \all_features[3757]  | \all_features[3758]  | \all_features[3759]  | (\all_features[3756]  & \all_features[3755]  & ~new_n19866_);
  assign new_n19866_ = ~\all_features[3754]  & new_n19854_;
  assign new_n19867_ = \all_features[3758]  | \all_features[3759]  | (new_n19869_ & new_n19868_);
  assign new_n19868_ = new_n19858_ & \all_features[3755]  & (\all_features[3754]  | (\all_features[3752]  & \all_features[3753] ));
  assign new_n19869_ = \all_features[3757]  & (\all_features[3756]  | (\all_features[3755]  & (\all_features[3754]  | \all_features[3753] )));
  assign new_n19870_ = \all_features[3759]  | (~new_n19872_ & ~new_n19871_ & \all_features[3758] );
  assign new_n19871_ = ~\all_features[3757]  & ~new_n19862_ & ~\all_features[3756] ;
  assign new_n19872_ = ~\all_features[3757]  & (new_n19854_ | ~\all_features[3756]  | ~new_n19862_);
  assign new_n19873_ = new_n19867_ & new_n19865_ & new_n19870_ & ~new_n19861_ & ~new_n19863_;
  assign new_n19874_ = new_n19867_ & new_n19865_ & (~new_n19875_ | (new_n19852_ & new_n19857_ & new_n19859_));
  assign new_n19875_ = ~new_n19861_ & (\all_features[3759]  | (new_n19864_ & \all_features[3758]  & ~new_n19872_ & ~new_n19871_));
  assign new_n19876_ = new_n19839_ & new_n19840_;
  assign new_n19877_ = (new_n19837_ | ~new_n19819_) & (~new_n6497_ | ~new_n19876_);
  assign new_n19878_ = new_n19830_ & new_n19833_;
  assign new_n19879_ = ~new_n19880_ & new_n19896_;
  assign new_n19880_ = ~new_n19835_ & new_n19881_ & ((~new_n17471_ & new_n19883_ & new_n18594_) | (~new_n19890_ & ~new_n18594_));
  assign new_n19881_ = new_n19882_ & (~new_n19835_ | (new_n19884_ & ~new_n16996_) | (new_n19887_ & new_n16996_));
  assign new_n19882_ = new_n19835_ | ~new_n18594_ | (new_n19883_ ? ~new_n17471_ : ~new_n18099_);
  assign new_n19883_ = ~new_n10273_ & new_n10248_;
  assign new_n19884_ = new_n19885_ ? ~new_n19678_ : ~new_n19886_;
  assign new_n19885_ = new_n17625_ & ~new_n12220_ & ~new_n17626_;
  assign new_n19886_ = new_n11094_ & (new_n11092_ | (new_n11083_ & new_n11063_));
  assign new_n19887_ = new_n18223_ ? ~new_n19889_ : new_n19888_;
  assign new_n19888_ = new_n12001_ & (new_n11978_ | ~new_n14085_);
  assign new_n19889_ = new_n17382_ & new_n17388_;
  assign new_n19890_ = new_n17635_ ? new_n19891_ : ~new_n19895_;
  assign new_n19891_ = new_n17250_ & (new_n12677_ | (~new_n19892_ & ~new_n12675_));
  assign new_n19892_ = ~new_n12678_ & (new_n12679_ | (~new_n12670_ & (new_n12672_ | (~new_n12668_ & ~new_n19893_))));
  assign new_n19893_ = ~new_n12673_ & (~new_n12666_ | (new_n12658_ & (~new_n12662_ | (~new_n19894_ & new_n12664_))));
  assign new_n19894_ = \all_features[3782]  & \all_features[3783]  & (\all_features[3781]  | (\all_features[3780]  & (\all_features[3779]  | \all_features[3778] )));
  assign new_n19895_ = ~new_n7935_ & new_n7942_;
  assign new_n19896_ = new_n19897_ & (new_n16996_ | ~new_n19835_ | (new_n19885_ ? new_n19678_ : new_n19886_));
  assign new_n19897_ = ~new_n19899_ & (new_n19835_ | ((new_n19898_ | new_n18594_) & (new_n18099_ | new_n19883_ | ~new_n18594_)));
  assign new_n19898_ = new_n17635_ ? ~new_n19891_ : new_n19895_;
  assign new_n19899_ = new_n16996_ & new_n19835_ & ~new_n19889_ & new_n18223_;
  assign \o[15]  = ~new_n19901_ ^ new_n19902_;
  assign new_n19901_ = (new_n19816_ & new_n19879_) | (~new_n17141_ & (new_n19816_ | new_n19879_));
  assign new_n19902_ = new_n19903_ ? (~new_n19904_ ^ new_n19953_) : (new_n19904_ ^ new_n19953_);
  assign new_n19903_ = (~new_n19031_ & new_n19730_) | (~new_n17142_ & (~new_n19031_ | new_n19730_));
  assign new_n19904_ = new_n19905_ ? (new_n19918_ ^ new_n19919_) : (~new_n19918_ ^ new_n19919_);
  assign new_n19905_ = new_n19906_ ? (~new_n19916_ ^ new_n19917_) : (new_n19916_ ^ new_n19917_);
  assign new_n19906_ = new_n19907_ ? (~new_n19914_ ^ new_n19915_) : (new_n19914_ ^ new_n19915_);
  assign new_n19907_ = new_n19908_ ? (~new_n19912_ ^ new_n19913_) : (new_n19912_ ^ new_n19913_);
  assign new_n19908_ = new_n19909_ ? (new_n19910_ ^ new_n19911_) : (~new_n19910_ ^ new_n19911_);
  assign new_n19909_ = new_n19035_ & new_n19131_;
  assign new_n19910_ = new_n17452_ & new_n17632_;
  assign new_n19911_ = new_n18909_ & new_n18955_;
  assign new_n19912_ = (new_n19155_ & new_n19242_) | (new_n19134_ & (new_n19155_ | new_n19242_));
  assign new_n19913_ = (~new_n17971_ & new_n17890_) | (new_n17810_ & (~new_n17971_ | new_n17890_));
  assign new_n19914_ = (~new_n19133_ & new_n17671_) | (new_n19034_ & (~new_n19133_ | new_n17671_));
  assign new_n19915_ = new_n19135_ & new_n19151_;
  assign new_n19916_ = (new_n18009_ & new_n18106_) | (~new_n17144_ & (new_n18009_ | new_n18106_));
  assign new_n19917_ = (new_n19334_ & new_n19419_) | (~new_n19033_ & (new_n19334_ | new_n19419_));
  assign new_n19918_ = (~new_n18112_ & new_n18957_) | (~new_n17143_ & (~new_n18112_ | new_n18957_));
  assign new_n19919_ = new_n19920_ ? (new_n19933_ ^ new_n19934_) : (~new_n19933_ ^ new_n19934_);
  assign new_n19920_ = new_n19921_ ? (~new_n19931_ ^ new_n19932_) : (new_n19931_ ^ new_n19932_);
  assign new_n19921_ = new_n19922_ ? (new_n19923_ ^ new_n19927_) : (~new_n19923_ ^ new_n19927_);
  assign new_n19922_ = (new_n17290_ & new_n17451_) | (new_n17146_ & (new_n17290_ | new_n17451_));
  assign new_n19923_ = new_n19924_ ? (new_n19925_ ^ new_n19926_) : (~new_n19925_ ^ new_n19926_);
  assign new_n19924_ = new_n18116_ & new_n18179_;
  assign new_n19925_ = new_n18010_ & new_n18103_;
  assign new_n19926_ = new_n19335_ & new_n19416_;
  assign new_n19927_ = new_n19928_ ? (new_n19929_ ^ new_n19930_) : (~new_n19929_ ^ new_n19930_);
  assign new_n19928_ = new_n18183_ & new_n18336_;
  assign new_n19929_ = new_n18666_ & new_n18787_;
  assign new_n19930_ = new_n18958_ & new_n19028_;
  assign new_n19931_ = (~new_n17809_ & new_n17671_) | (~new_n17145_ & (~new_n17809_ | new_n17671_));
  assign new_n19932_ = (new_n18338_ & new_n18339_) | (~new_n18114_ & (new_n18338_ | new_n18339_));
  assign new_n19933_ = (~new_n18372_ & new_n18908_) | (~new_n18113_ & (~new_n18372_ | new_n18908_));
  assign new_n19934_ = new_n19935_ ? (new_n19943_ ^ new_n19944_) : (~new_n19943_ ^ new_n19944_);
  assign new_n19935_ = new_n19936_ ? (~new_n19937_ ^ new_n19942_) : (new_n19937_ ^ new_n19942_);
  assign new_n19936_ = (new_n18182_ & new_n18337_) | (new_n18115_ & (new_n18182_ | new_n18337_));
  assign new_n19937_ = new_n19938_ ? (new_n19940_ ^ new_n19941_) : (~new_n19940_ ^ new_n19941_);
  assign new_n19938_ = new_n19731_ & ~new_n19939_ & new_n19775_;
  assign new_n19939_ = ~new_n19814_ & ~new_n19815_;
  assign new_n19940_ = new_n19503_ & new_n19588_;
  assign new_n19941_ = new_n18791_ & new_n18848_;
  assign new_n19942_ = (new_n18790_ & new_n18852_) | (new_n18665_ & (new_n18790_ | new_n18852_));
  assign new_n19943_ = (~new_n18373_ & ~new_n18664_) | (new_n18338_ & (~new_n18373_ | ~new_n18664_));
  assign new_n19944_ = new_n19945_ ? (~new_n19946_ ^ new_n19949_) : (new_n19946_ ^ new_n19949_);
  assign new_n19945_ = ~new_n18374_ & ~new_n18570_;
  assign new_n19946_ = new_n19947_ ^ new_n19948_;
  assign new_n19947_ = new_n19817_ & new_n19847_;
  assign new_n19948_ = new_n18375_ & new_n18544_;
  assign new_n19949_ = new_n19950_ ? (new_n19951_ ^ new_n19952_) : (~new_n19951_ ^ new_n19952_);
  assign new_n19950_ = new_n18853_ & new_n18904_;
  assign new_n19951_ = new_n19896_ & new_n19881_;
  assign new_n19952_ = new_n18571_ & new_n18591_;
  assign new_n19953_ = (new_n19502_ & new_n19593_) | (~new_n19032_ & (new_n19502_ | new_n19593_));
  assign \o[16]  = ~new_n19955_ ^ new_n19956_;
  assign new_n19955_ = ~new_n19902_ & new_n19901_;
  assign new_n19956_ = new_n19957_ ^ new_n19958_;
  assign new_n19957_ = (~new_n19904_ & new_n19953_) | (new_n19903_ & (~new_n19904_ | new_n19953_));
  assign new_n19958_ = new_n19959_ ? (~new_n19960_ ^ new_n19989_) : (new_n19960_ ^ new_n19989_);
  assign new_n19959_ = (~new_n19919_ & new_n19918_) | (~new_n19905_ & (~new_n19919_ | new_n19918_));
  assign new_n19960_ = new_n19961_ ? (new_n19969_ ^ new_n19970_) : (~new_n19969_ ^ new_n19970_);
  assign new_n19961_ = new_n19962_ ? (~new_n19963_ ^ new_n19968_) : (new_n19963_ ^ new_n19968_);
  assign new_n19962_ = (new_n19914_ & new_n19915_) | (~new_n19907_ & (new_n19914_ | new_n19915_));
  assign new_n19963_ = ~new_n19964_ ^ new_n19965_;
  assign new_n19964_ = (new_n19912_ & new_n19913_) | (~new_n19908_ & (new_n19912_ | new_n19913_));
  assign new_n19965_ = new_n19966_ ^ new_n19967_;
  assign new_n19966_ = (new_n19910_ & new_n19911_) | (new_n19909_ & (new_n19910_ | new_n19911_));
  assign new_n19967_ = (new_n19925_ & new_n19926_) | (new_n19924_ & (new_n19925_ | new_n19926_));
  assign new_n19968_ = (new_n19931_ & new_n19932_) | (~new_n19921_ & (new_n19931_ | new_n19932_));
  assign new_n19969_ = (~new_n19934_ & new_n19933_) | (~new_n19920_ & (~new_n19934_ | new_n19933_));
  assign new_n19970_ = new_n19971_ ? (new_n19975_ ^ new_n19976_) : (~new_n19975_ ^ new_n19976_);
  assign new_n19971_ = new_n19972_ ? (new_n19973_ ^ new_n19974_) : (~new_n19973_ ^ new_n19974_);
  assign new_n19972_ = (~new_n19923_ & ~new_n19927_) | (new_n19922_ & (~new_n19923_ | ~new_n19927_));
  assign new_n19973_ = (~new_n19937_ & new_n19942_) | (new_n19936_ & (~new_n19937_ | new_n19942_));
  assign new_n19974_ = (new_n19929_ & new_n19930_) | (new_n19928_ & (new_n19929_ | new_n19930_));
  assign new_n19975_ = (~new_n19944_ & new_n19943_) | (~new_n19935_ & (~new_n19944_ | new_n19943_));
  assign new_n19976_ = new_n19977_ ? (new_n19978_ ^ new_n19986_) : (~new_n19978_ ^ new_n19986_);
  assign new_n19977_ = (~new_n19946_ & ~new_n19949_) | (~new_n19945_ & (~new_n19946_ | ~new_n19949_));
  assign new_n19978_ = new_n19979_ ? (~new_n19980_ ^ new_n19983_) : (new_n19980_ ^ new_n19983_);
  assign new_n19979_ = ~new_n19947_ & ~new_n19948_;
  assign new_n19980_ = ~new_n19981_ ^ new_n19982_;
  assign new_n19981_ = new_n19939_ & new_n19731_ & new_n19775_;
  assign new_n19982_ = new_n19594_ & new_n19728_;
  assign new_n19983_ = new_n19984_ ^ new_n19985_;
  assign new_n19984_ = new_n19817_ & new_n19877_ & ~new_n19878_ & new_n19847_;
  assign new_n19985_ = new_n18477_ & new_n18544_ & new_n18376_;
  assign new_n19986_ = ~new_n19987_ ^ new_n19988_;
  assign new_n19987_ = (new_n19940_ & new_n19941_) | (new_n19938_ & (new_n19940_ | new_n19941_));
  assign new_n19988_ = (new_n19951_ & new_n19952_) | (new_n19950_ & (new_n19951_ | new_n19952_));
  assign new_n19989_ = (new_n19916_ & new_n19917_) | (~new_n19906_ & (new_n19916_ | new_n19917_));
  assign \o[17]  = ((new_n19991_ | new_n19992_) & (new_n19993_ ^ new_n19994_)) | (~new_n19991_ & ~new_n19992_ & (~new_n19993_ ^ new_n19994_));
  assign new_n19991_ = ~new_n19956_ & new_n19955_;
  assign new_n19992_ = ~new_n19958_ & new_n19957_;
  assign new_n19993_ = (~new_n19960_ & new_n19989_) | (new_n19959_ & (~new_n19960_ | new_n19989_));
  assign new_n19994_ = new_n19995_ ? (~new_n19996_ ^ new_n20009_) : (new_n19996_ ^ new_n20009_);
  assign new_n19995_ = (~new_n19970_ & new_n19969_) | (~new_n19961_ & (~new_n19970_ | new_n19969_));
  assign new_n19996_ = new_n19997_ ? (new_n20001_ ^ new_n20002_) : (~new_n20001_ ^ new_n20002_);
  assign new_n19997_ = new_n19998_ ? (new_n19999_ ^ new_n20000_) : (~new_n19999_ ^ new_n20000_);
  assign new_n19998_ = new_n19964_ & new_n19965_;
  assign new_n19999_ = (new_n19973_ & new_n19974_) | (new_n19972_ & (new_n19973_ | new_n19974_));
  assign new_n20000_ = new_n19966_ & new_n19967_;
  assign new_n20001_ = (~new_n19976_ & new_n19975_) | (~new_n19971_ & (~new_n19976_ | new_n19975_));
  assign new_n20002_ = new_n20003_ ? (~new_n20004_ ^ new_n20008_) : (new_n20004_ ^ new_n20008_);
  assign new_n20003_ = (~new_n19978_ & ~new_n19986_) | (new_n19977_ & (~new_n19978_ | ~new_n19986_));
  assign new_n20004_ = new_n20005_ ? (~new_n20006_ ^ new_n20007_) : (new_n20006_ ^ new_n20007_);
  assign new_n20005_ = (~new_n19980_ & ~new_n19983_) | (~new_n19979_ & (~new_n19980_ | ~new_n19983_));
  assign new_n20006_ = ~new_n19984_ & ~new_n19985_;
  assign new_n20007_ = new_n19981_ & new_n19982_;
  assign new_n20008_ = new_n19987_ & new_n19988_;
  assign new_n20009_ = (~new_n19963_ & new_n19968_) | (new_n19962_ & (~new_n19963_ | new_n19968_));
  assign \o[18]  = ~new_n20011_ ^ new_n20012_;
  assign new_n20011_ = (new_n19993_ | (~new_n19994_ & (new_n19992_ | new_n19991_))) & (new_n19992_ | new_n19991_ | ~new_n19994_);
  assign new_n20012_ = new_n20013_ ^ new_n20014_;
  assign new_n20013_ = (~new_n19996_ & new_n20009_) | (new_n19995_ & (~new_n19996_ | new_n20009_));
  assign new_n20014_ = new_n20015_ ? (~new_n20016_ ^ new_n20019_) : (new_n20016_ ^ new_n20019_);
  assign new_n20015_ = (~new_n20002_ & new_n20001_) | (~new_n19997_ & (~new_n20002_ | new_n20001_));
  assign new_n20016_ = ~new_n20017_ ^ new_n20018_;
  assign new_n20017_ = (~new_n20004_ & new_n20008_) | (new_n20003_ & (~new_n20004_ | new_n20008_));
  assign new_n20018_ = (~new_n20006_ & new_n20007_) | (new_n20005_ & (~new_n20006_ | new_n20007_));
  assign new_n20019_ = (new_n19999_ & new_n20000_) | (new_n19998_ & (new_n19999_ | new_n20000_));
  assign \o[19]  = ((new_n20021_ | new_n20022_) & (~new_n20023_ ^ new_n20024_)) | (~new_n20021_ & ~new_n20022_ & (new_n20023_ ^ new_n20024_));
  assign new_n20021_ = ~new_n20012_ & new_n20011_;
  assign new_n20022_ = ~new_n20014_ & new_n20013_;
  assign new_n20023_ = (~new_n20016_ & new_n20019_) | (new_n20015_ & (~new_n20016_ | new_n20019_));
  assign new_n20024_ = new_n20017_ & new_n20018_;
  assign \o[20]  = (new_n20024_ | new_n20021_ | new_n20022_) & (new_n20023_ | (new_n20024_ & (new_n20021_ | new_n20022_)));
  assign \o[21]  = new_n20027_ ? (new_n21945_ ^ new_n22046_) : (~new_n21945_ ^ new_n22046_);
  assign new_n20027_ = new_n20028_ ? (~new_n21761_ ^ new_n21847_) : (new_n21761_ ^ new_n21847_);
  assign new_n20028_ = new_n20029_ ? (new_n21393_ ^ new_n21698_) : (~new_n21393_ ^ new_n21698_);
  assign new_n20029_ = new_n20030_ ? (new_n20873_ ^ new_n21392_) : (~new_n20873_ ^ new_n21392_);
  assign new_n20030_ = new_n20031_ ? (new_n20451_ ^ new_n20805_) : (~new_n20451_ ^ new_n20805_);
  assign new_n20031_ = new_n20032_ ? (~new_n20236_ ^ new_n20269_) : (new_n20236_ ^ new_n20269_);
  assign new_n20032_ = new_n20033_ ? (new_n20092_ ^ new_n20148_) : (~new_n20092_ ^ new_n20148_);
  assign new_n20033_ = ~new_n20034_ & new_n20089_;
  assign new_n20034_ = new_n20035_ & (~new_n20088_ | ~new_n20082_) & (~new_n20084_ | ~new_n20083_);
  assign new_n20035_ = new_n20036_ & (~new_n20050_ | (new_n8164_ & ~new_n18421_) | (new_n20051_ & new_n18421_));
  assign new_n20036_ = ~new_n20037_ & (~new_n20044_ | (new_n20047_ & new_n20046_) | (new_n20049_ & ~new_n20046_));
  assign new_n20037_ = ~new_n20042_ & ~new_n13038_ & new_n20038_ & (~new_n13015_ | ~new_n17844_);
  assign new_n20038_ = new_n20039_ & new_n20040_;
  assign new_n20039_ = ~new_n19158_ & new_n16215_;
  assign new_n20040_ = new_n10478_ & (new_n10456_ | new_n20041_);
  assign new_n20041_ = new_n10481_ & new_n10485_;
  assign new_n20042_ = ~new_n12115_ & (~new_n12112_ | ~new_n20043_);
  assign new_n20043_ = new_n12084_ & new_n12108_;
  assign new_n20044_ = ~new_n20039_ & new_n20045_;
  assign new_n20045_ = ~new_n12187_ & new_n12729_;
  assign new_n20046_ = new_n8735_ & new_n8725_;
  assign new_n20047_ = ~new_n6702_ & new_n20048_;
  assign new_n20048_ = new_n6732_ & new_n6734_;
  assign new_n20049_ = ~new_n15495_ & new_n8165_;
  assign new_n20050_ = ~new_n20039_ & ~new_n20045_;
  assign new_n20051_ = ~new_n20080_ & (~new_n20077_ | ~new_n20052_);
  assign new_n20052_ = new_n20072_ & (~new_n20068_ | (new_n20064_ & (new_n20053_ | new_n20074_ | new_n20076_)));
  assign new_n20053_ = new_n20062_ & new_n20063_ & (~new_n20059_ | ~new_n20057_ | new_n20054_);
  assign new_n20054_ = \all_features[5431]  & \all_features[5430]  & ~new_n20055_ & \all_features[5429] ;
  assign new_n20055_ = ~\all_features[5427]  & ~\all_features[5428]  & (~\all_features[5426]  | new_n20056_);
  assign new_n20056_ = ~\all_features[5424]  & ~\all_features[5425] ;
  assign new_n20057_ = \all_features[5431]  & (\all_features[5430]  | (new_n20058_ & (\all_features[5426]  | \all_features[5427]  | \all_features[5425] )));
  assign new_n20058_ = \all_features[5428]  & \all_features[5429] ;
  assign new_n20059_ = \all_features[5430]  & \all_features[5431]  & (\all_features[5428]  | \all_features[5429]  | new_n20060_ | ~new_n20061_);
  assign new_n20060_ = \all_features[5424]  & \all_features[5425] ;
  assign new_n20061_ = ~\all_features[5426]  & ~\all_features[5427] ;
  assign new_n20062_ = \all_features[5431]  & (\all_features[5430]  | (\all_features[5429]  & (\all_features[5428]  | ~new_n20061_ | ~new_n20056_)));
  assign new_n20063_ = \all_features[5431]  & (\all_features[5429]  | \all_features[5430]  | \all_features[5428] );
  assign new_n20064_ = ~new_n20065_ & ~new_n20067_;
  assign new_n20065_ = ~\all_features[5431]  & (~\all_features[5430]  | (~\all_features[5428]  & ~\all_features[5429]  & ~new_n20066_));
  assign new_n20066_ = \all_features[5426]  & \all_features[5427] ;
  assign new_n20067_ = ~\all_features[5431]  & (~\all_features[5430]  | (~\all_features[5429]  & (new_n20056_ | ~\all_features[5428]  | ~new_n20066_)));
  assign new_n20068_ = ~new_n20069_ & ~new_n20071_;
  assign new_n20069_ = new_n20070_ & (~\all_features[5429]  | (~\all_features[5428]  & (~\all_features[5427]  | (~\all_features[5426]  & ~\all_features[5425] ))));
  assign new_n20070_ = ~\all_features[5430]  & ~\all_features[5431] ;
  assign new_n20071_ = new_n20070_ & (~\all_features[5427]  | ~new_n20058_ | (~\all_features[5426]  & ~new_n20060_));
  assign new_n20072_ = ~new_n20073_ & (\all_features[5427]  | \all_features[5428]  | \all_features[5429]  | \all_features[5430]  | \all_features[5431] );
  assign new_n20073_ = ~\all_features[5429]  & new_n20070_ & ((~\all_features[5426]  & new_n20056_) | ~\all_features[5428]  | ~\all_features[5427] );
  assign new_n20074_ = ~new_n20075_ & ~\all_features[5431] ;
  assign new_n20075_ = \all_features[5429]  & \all_features[5430]  & (\all_features[5428]  | (\all_features[5426]  & \all_features[5427]  & \all_features[5425] ));
  assign new_n20076_ = ~\all_features[5431]  & (~\all_features[5430]  | ~new_n20066_ | ~new_n20060_ | ~new_n20058_);
  assign new_n20077_ = new_n20072_ & ~new_n20078_ & new_n20068_;
  assign new_n20078_ = new_n20079_ & (~new_n20062_ | ~new_n20063_ | ~new_n20057_ | ~new_n20059_);
  assign new_n20079_ = ~new_n20076_ & ~new_n20074_ & ~new_n20065_ & ~new_n20067_;
  assign new_n20080_ = new_n20068_ & new_n20064_ & new_n20081_ & ~new_n20074_ & ~new_n20073_;
  assign new_n20081_ = ~new_n20076_ & (\all_features[5427]  | \all_features[5428]  | \all_features[5429]  | \all_features[5430]  | \all_features[5431] );
  assign new_n20082_ = new_n20038_ & new_n20042_;
  assign new_n20083_ = ~new_n20040_ & new_n20039_;
  assign new_n20084_ = new_n20085_ ? new_n20087_ : new_n10910_;
  assign new_n20085_ = ~new_n10677_ & (~new_n10679_ | ~new_n20086_);
  assign new_n20086_ = new_n10649_ & new_n10670_;
  assign new_n20087_ = new_n7269_ & ~new_n7295_ & ~new_n7299_;
  assign new_n20088_ = ~new_n10677_ & new_n13942_;
  assign new_n20089_ = new_n20090_ & (new_n20084_ | ~new_n20083_) & (~new_n20082_ | new_n20088_);
  assign new_n20090_ = ~new_n20091_ & (~new_n20044_ | (~new_n20047_ & new_n20046_) | (~new_n20049_ & ~new_n20046_));
  assign new_n20091_ = new_n20050_ & (new_n18421_ ? new_n20051_ : new_n8164_);
  assign new_n20092_ = ~new_n20093_ & ~new_n20147_;
  assign new_n20093_ = new_n20094_ & (new_n20096_ | ((new_n17974_ | ~new_n10205_) & (new_n20102_ | new_n20118_ | new_n10205_)));
  assign new_n20094_ = ~new_n20095_ & ((new_n20111_ & (new_n20112_ | ~new_n20116_)) | ~new_n20096_ | (new_n20117_ & ~new_n20112_ & ~new_n20116_));
  assign new_n20095_ = ~new_n10205_ & ~new_n20096_ & new_n20102_ & (~new_n15247_ | ~new_n20103_);
  assign new_n20096_ = ~new_n20097_ & new_n19238_;
  assign new_n20097_ = new_n6974_ & new_n20098_;
  assign new_n20098_ = ~new_n20099_ & (\all_features[3091]  | \all_features[3092]  | \all_features[3093]  | \all_features[3094]  | \all_features[3095] );
  assign new_n20099_ = ~new_n6991_ & (new_n6994_ | (~new_n6995_ & (new_n6997_ | (~new_n6996_ & ~new_n20100_))));
  assign new_n20100_ = ~new_n6984_ & (new_n6986_ | (new_n6989_ & (~new_n6988_ | (~new_n20101_ & new_n6977_))));
  assign new_n20101_ = ~\all_features[3093]  & \all_features[3094]  & \all_features[3095]  & (\all_features[3092]  ? new_n6981_ : (new_n6980_ | ~new_n6981_));
  assign new_n20102_ = ~new_n17845_ & new_n13837_;
  assign new_n20103_ = ~new_n15260_ & ~new_n15256_ & ~new_n15252_ & ~new_n20104_ & ~new_n15262_;
  assign new_n20104_ = ~new_n15261_ & ~new_n15263_ & ~new_n15257_ & ~new_n15248_ & ~new_n20105_;
  assign new_n20105_ = new_n20110_ & new_n20109_ & new_n20106_ & new_n20108_;
  assign new_n20106_ = \all_features[1231]  & (\all_features[1230]  | (\all_features[1229]  & (\all_features[1228]  | ~new_n20107_ | ~new_n15250_)));
  assign new_n20107_ = ~\all_features[1226]  & ~\all_features[1227] ;
  assign new_n20108_ = \all_features[1231]  & (\all_features[1230]  | (new_n15255_ & (\all_features[1226]  | \all_features[1227]  | \all_features[1225] )));
  assign new_n20109_ = \all_features[1230]  & \all_features[1231]  & (\all_features[1228]  | \all_features[1229]  | new_n15254_ | ~new_n20107_);
  assign new_n20110_ = \all_features[1231]  & (\all_features[1229]  | \all_features[1230]  | \all_features[1228] );
  assign new_n20111_ = new_n16639_ & new_n20112_ & new_n20113_;
  assign new_n20112_ = new_n18158_ & new_n10513_;
  assign new_n20113_ = ~new_n20114_ & new_n20115_;
  assign new_n20114_ = ~new_n14014_ & ~new_n16364_;
  assign new_n20115_ = new_n14039_ & new_n14042_;
  assign new_n20116_ = ~new_n14679_ & (~new_n14656_ | new_n14681_);
  assign new_n20117_ = new_n12301_ & (new_n12298_ | new_n18188_);
  assign new_n20118_ = ~new_n20143_ & new_n20119_;
  assign new_n20119_ = new_n20142_ | ~new_n20140_ | ((new_n20131_ | new_n20129_) & (new_n20137_ | ~new_n20120_));
  assign new_n20120_ = new_n20121_ & ~new_n20127_ & ~new_n20129_;
  assign new_n20121_ = ~new_n20122_ & ~new_n20126_;
  assign new_n20122_ = ~\all_features[4295]  & (~\all_features[4294]  | ~new_n20123_ | ~new_n20124_ | ~new_n20125_);
  assign new_n20123_ = \all_features[4290]  & \all_features[4291] ;
  assign new_n20124_ = \all_features[4288]  & \all_features[4289] ;
  assign new_n20125_ = \all_features[4292]  & \all_features[4293] ;
  assign new_n20126_ = ~\all_features[4295]  & (~\all_features[4294]  | (~\all_features[4292]  & ~\all_features[4293]  & ~new_n20123_));
  assign new_n20127_ = ~\all_features[4295]  & (~\all_features[4294]  | (~\all_features[4293]  & (new_n20128_ | ~new_n20123_ | ~\all_features[4292] )));
  assign new_n20128_ = ~\all_features[4288]  & ~\all_features[4289] ;
  assign new_n20129_ = new_n20130_ & (~\all_features[4291]  | ~new_n20125_ | (~\all_features[4290]  & ~new_n20124_));
  assign new_n20130_ = ~\all_features[4294]  & ~\all_features[4295] ;
  assign new_n20131_ = ~new_n20137_ & ~new_n20127_ & new_n20121_ & (~new_n20139_ | ~new_n20132_);
  assign new_n20132_ = new_n20136_ & new_n20133_ & new_n20134_;
  assign new_n20133_ = \all_features[4295]  & (\all_features[4294]  | (new_n20125_ & (\all_features[4290]  | \all_features[4291]  | \all_features[4289] )));
  assign new_n20134_ = \all_features[4294]  & \all_features[4295]  & (\all_features[4292]  | \all_features[4293]  | new_n20124_ | ~new_n20135_);
  assign new_n20135_ = ~\all_features[4290]  & ~\all_features[4291] ;
  assign new_n20136_ = \all_features[4295]  & (\all_features[4293]  | \all_features[4294]  | \all_features[4292] );
  assign new_n20137_ = ~new_n20138_ & ~\all_features[4295] ;
  assign new_n20138_ = \all_features[4293]  & \all_features[4294]  & (\all_features[4292]  | (\all_features[4290]  & \all_features[4291]  & \all_features[4289] ));
  assign new_n20139_ = \all_features[4295]  & (\all_features[4294]  | (\all_features[4293]  & (\all_features[4292]  | ~new_n20135_ | ~new_n20128_)));
  assign new_n20140_ = ~new_n20141_ & (\all_features[4291]  | \all_features[4292]  | \all_features[4293]  | \all_features[4294]  | \all_features[4295] );
  assign new_n20141_ = ~\all_features[4293]  & new_n20130_ & ((~\all_features[4290]  & new_n20128_) | ~\all_features[4292]  | ~\all_features[4291] );
  assign new_n20142_ = new_n20130_ & (~\all_features[4293]  | (~\all_features[4292]  & (~\all_features[4291]  | (~\all_features[4290]  & ~\all_features[4289] ))));
  assign new_n20143_ = new_n20140_ & (new_n20129_ | new_n20142_ | (~new_n20144_ & ~new_n20127_ & ~new_n20126_));
  assign new_n20144_ = ~new_n20137_ & ~new_n20122_ & (~new_n20136_ | ~new_n20139_ | new_n20145_);
  assign new_n20145_ = new_n20133_ & new_n20134_ & (new_n20146_ | ~\all_features[4293]  | ~\all_features[4294]  | ~\all_features[4295] );
  assign new_n20146_ = ~\all_features[4291]  & ~\all_features[4292]  & (~\all_features[4290]  | new_n20128_);
  assign new_n20147_ = ~new_n20096_ & ((~new_n20102_ & new_n20118_ & ~new_n10205_) | (new_n17974_ & new_n10205_));
  assign new_n20148_ = new_n20170_ & (new_n20149_ | new_n20171_) & (new_n20157_ | new_n15164_ | ~new_n14046_ | ~new_n20171_);
  assign new_n20149_ = new_n20116_ ? (new_n20155_ | (new_n20156_ & new_n17176_)) : ~new_n20150_;
  assign new_n20150_ = new_n16612_ & (~new_n20151_ | ~new_n16640_);
  assign new_n20151_ = ~new_n16633_ & (new_n16632_ | new_n20152_);
  assign new_n20152_ = ~new_n16628_ & (new_n16630_ | (~new_n16623_ & (new_n16624_ | (~new_n16616_ & ~new_n20153_))));
  assign new_n20153_ = ~new_n16618_ & (~new_n16638_ | (new_n16637_ & (~new_n16634_ | (~new_n20154_ & new_n16635_))));
  assign new_n20154_ = \all_features[4430]  & \all_features[4431]  & (\all_features[4429]  | (~new_n16636_ & \all_features[4428] ));
  assign new_n20155_ = new_n15831_ & new_n16106_;
  assign new_n20156_ = new_n17154_ & new_n17178_;
  assign new_n20157_ = (new_n8927_ & (~new_n8893_ | new_n8924_)) ? new_n20168_ : ~new_n20158_;
  assign new_n20158_ = ~new_n20159_ & new_n17816_;
  assign new_n20159_ = ~new_n20160_ & ~new_n20164_;
  assign new_n20160_ = new_n17835_ & (~new_n17841_ | (~new_n20161_ & ~new_n17829_ & ~new_n17833_));
  assign new_n20161_ = ~new_n17834_ & ~new_n17827_ & (~new_n17825_ | ~new_n17831_ | new_n20162_);
  assign new_n20162_ = new_n17820_ & new_n17822_ & (new_n20163_ | ~\all_features[4813]  | ~\all_features[4814]  | ~\all_features[4815] );
  assign new_n20163_ = ~\all_features[4811]  & ~\all_features[4812]  & (~\all_features[4810]  | new_n17832_);
  assign new_n20164_ = ~new_n20165_ & (\all_features[4811]  | \all_features[4812]  | \all_features[4813]  | \all_features[4814]  | \all_features[4815] );
  assign new_n20165_ = ~new_n17836_ & (new_n17838_ | (~new_n17839_ & (new_n17829_ | (~new_n17833_ & ~new_n20166_))));
  assign new_n20166_ = ~new_n17827_ & (new_n17834_ | (new_n17825_ & (~new_n17831_ | (~new_n20167_ & new_n17820_))));
  assign new_n20167_ = ~\all_features[4813]  & \all_features[4814]  & \all_features[4815]  & (\all_features[4812]  ? new_n17823_ : (new_n17824_ | ~new_n17823_));
  assign new_n20168_ = ~new_n20169_ & new_n12721_;
  assign new_n20169_ = ~new_n12709_ & ~new_n12718_;
  assign new_n20170_ = (new_n20150_ | new_n20116_ | ~new_n20235_ | new_n20171_) & (~new_n20233_ | ~new_n20206_ | ~new_n20171_);
  assign new_n20171_ = ~new_n20172_ & new_n20201_;
  assign new_n20172_ = ~new_n20173_ & ~new_n20194_;
  assign new_n20173_ = ~new_n20174_ & (\all_features[1691]  | \all_features[1692]  | \all_features[1693]  | \all_features[1694]  | \all_features[1695] );
  assign new_n20174_ = ~new_n20188_ & (new_n20190_ | (~new_n20191_ & (new_n20192_ | (~new_n20175_ & ~new_n20193_))));
  assign new_n20175_ = ~new_n20176_ & (new_n20185_ | (new_n20187_ & (~new_n20178_ | (~new_n20183_ & new_n20181_))));
  assign new_n20176_ = ~new_n20177_ & ~\all_features[1695] ;
  assign new_n20177_ = \all_features[1693]  & \all_features[1694]  & (\all_features[1692]  | (\all_features[1690]  & \all_features[1691]  & \all_features[1689] ));
  assign new_n20178_ = \all_features[1695]  & (\all_features[1694]  | (\all_features[1693]  & (\all_features[1692]  | ~new_n20180_ | ~new_n20179_)));
  assign new_n20179_ = ~\all_features[1688]  & ~\all_features[1689] ;
  assign new_n20180_ = ~\all_features[1690]  & ~\all_features[1691] ;
  assign new_n20181_ = \all_features[1695]  & (\all_features[1694]  | (new_n20182_ & (\all_features[1690]  | \all_features[1691]  | \all_features[1689] )));
  assign new_n20182_ = \all_features[1692]  & \all_features[1693] ;
  assign new_n20183_ = ~\all_features[1693]  & \all_features[1694]  & \all_features[1695]  & (\all_features[1692]  ? new_n20180_ : (new_n20184_ | ~new_n20180_));
  assign new_n20184_ = \all_features[1688]  & \all_features[1689] ;
  assign new_n20185_ = ~\all_features[1695]  & (~\all_features[1694]  | ~new_n20184_ | ~new_n20182_ | ~new_n20186_);
  assign new_n20186_ = \all_features[1690]  & \all_features[1691] ;
  assign new_n20187_ = \all_features[1695]  & (\all_features[1693]  | \all_features[1694]  | \all_features[1692] );
  assign new_n20188_ = ~\all_features[1693]  & new_n20189_ & ((~\all_features[1690]  & new_n20179_) | ~\all_features[1692]  | ~\all_features[1691] );
  assign new_n20189_ = ~\all_features[1694]  & ~\all_features[1695] ;
  assign new_n20190_ = new_n20189_ & (~\all_features[1693]  | (~\all_features[1692]  & (~\all_features[1691]  | (~\all_features[1690]  & ~\all_features[1689] ))));
  assign new_n20191_ = new_n20189_ & (~\all_features[1691]  | ~new_n20182_ | (~\all_features[1690]  & ~new_n20184_));
  assign new_n20192_ = ~\all_features[1695]  & (~\all_features[1694]  | (~\all_features[1692]  & ~\all_features[1693]  & ~new_n20186_));
  assign new_n20193_ = ~\all_features[1695]  & (~\all_features[1694]  | (~\all_features[1693]  & (new_n20179_ | ~new_n20186_ | ~\all_features[1692] )));
  assign new_n20194_ = new_n20200_ & (~new_n20199_ | (~new_n20195_ & ~new_n20192_ & ~new_n20193_));
  assign new_n20195_ = ~new_n20185_ & ~new_n20176_ & (~new_n20187_ | ~new_n20178_ | new_n20196_);
  assign new_n20196_ = new_n20181_ & new_n20197_ & (new_n20198_ | ~\all_features[1693]  | ~\all_features[1694]  | ~\all_features[1695] );
  assign new_n20197_ = \all_features[1694]  & \all_features[1695]  & (\all_features[1692]  | \all_features[1693]  | new_n20184_ | ~new_n20180_);
  assign new_n20198_ = ~\all_features[1691]  & ~\all_features[1692]  & (~\all_features[1690]  | new_n20179_);
  assign new_n20199_ = ~new_n20190_ & ~new_n20191_;
  assign new_n20200_ = ~new_n20188_ & (\all_features[1691]  | \all_features[1692]  | \all_features[1693]  | \all_features[1694]  | \all_features[1695] );
  assign new_n20201_ = new_n20202_ & new_n20205_;
  assign new_n20202_ = new_n20199_ & new_n20200_ & (new_n20203_ | new_n20193_ | new_n20185_ | ~new_n20204_);
  assign new_n20203_ = new_n20187_ & new_n20197_ & new_n20178_ & new_n20181_;
  assign new_n20204_ = ~new_n20192_ & ~new_n20176_;
  assign new_n20205_ = new_n20200_ & new_n20199_ & new_n20204_ & ~new_n20193_ & ~new_n20185_;
  assign new_n20206_ = (~new_n20207_ | ~new_n20232_) & (new_n15164_ | ~new_n14046_);
  assign new_n20207_ = new_n20218_ & new_n20226_ & (new_n20208_ | new_n20229_ | new_n20231_ | ~new_n20222_);
  assign new_n20208_ = new_n20217_ & new_n20215_ & new_n20209_ & new_n20212_;
  assign new_n20209_ = \all_features[1007]  & (\all_features[1006]  | new_n20210_);
  assign new_n20210_ = \all_features[1005]  & (\all_features[1002]  | \all_features[1003]  | \all_features[1004]  | ~new_n20211_);
  assign new_n20211_ = ~\all_features[1000]  & ~\all_features[1001] ;
  assign new_n20212_ = \all_features[1007]  & ~new_n20213_ & \all_features[1006] ;
  assign new_n20213_ = ~\all_features[1005]  & ~\all_features[1004]  & ~\all_features[1003]  & ~new_n20214_ & ~\all_features[1002] ;
  assign new_n20214_ = \all_features[1000]  & \all_features[1001] ;
  assign new_n20215_ = \all_features[1007]  & (\all_features[1006]  | (new_n20216_ & (\all_features[1002]  | \all_features[1003]  | \all_features[1001] )));
  assign new_n20216_ = \all_features[1004]  & \all_features[1005] ;
  assign new_n20217_ = \all_features[1007]  & (\all_features[1005]  | \all_features[1006]  | \all_features[1004] );
  assign new_n20218_ = ~new_n20219_ & ~new_n20221_;
  assign new_n20219_ = ~\all_features[1005]  & new_n20220_ & ((~\all_features[1002]  & new_n20211_) | ~\all_features[1004]  | ~\all_features[1003] );
  assign new_n20220_ = ~\all_features[1006]  & ~\all_features[1007] ;
  assign new_n20221_ = ~\all_features[1007]  & ~\all_features[1006]  & ~\all_features[1005]  & ~\all_features[1003]  & ~\all_features[1004] ;
  assign new_n20222_ = ~new_n20223_ & ~new_n20225_;
  assign new_n20223_ = ~\all_features[1007]  & (~\all_features[1006]  | ~new_n20224_ | ~new_n20214_ | ~new_n20216_);
  assign new_n20224_ = \all_features[1002]  & \all_features[1003] ;
  assign new_n20225_ = ~\all_features[1007]  & (~\all_features[1006]  | (~\all_features[1004]  & ~\all_features[1005]  & ~new_n20224_));
  assign new_n20226_ = ~new_n20227_ & ~new_n20228_;
  assign new_n20227_ = new_n20220_ & (~\all_features[1005]  | (~\all_features[1004]  & (~\all_features[1003]  | (~\all_features[1002]  & ~\all_features[1001] ))));
  assign new_n20228_ = new_n20220_ & (~\all_features[1003]  | ~new_n20216_ | (~\all_features[1002]  & ~new_n20214_));
  assign new_n20229_ = ~new_n20230_ & ~\all_features[1007] ;
  assign new_n20230_ = \all_features[1005]  & \all_features[1006]  & (\all_features[1004]  | (\all_features[1002]  & \all_features[1003]  & \all_features[1001] ));
  assign new_n20231_ = ~\all_features[1007]  & (~\all_features[1006]  | (~\all_features[1005]  & (new_n20211_ | ~new_n20224_ | ~\all_features[1004] )));
  assign new_n20232_ = new_n20222_ & new_n20218_ & ~new_n20228_ & ~new_n20231_ & ~new_n20229_ & ~new_n20227_;
  assign new_n20233_ = new_n10490_ & new_n20234_;
  assign new_n20234_ = ~new_n10516_ & ~new_n10520_;
  assign new_n20235_ = ~new_n16231_ & ~new_n9018_;
  assign new_n20236_ = new_n20237_ & new_n20266_;
  assign new_n20237_ = new_n20238_ & new_n20249_;
  assign new_n20238_ = (~new_n20239_ | new_n20248_) & (~new_n20244_ | (new_n20245_ ? ~new_n20115_ : new_n20247_));
  assign new_n20239_ = ~new_n18786_ & new_n20240_;
  assign new_n20240_ = ~new_n20241_ & new_n20243_;
  assign new_n20241_ = ~new_n20242_ & new_n6490_;
  assign new_n20242_ = ~new_n6462_ & ~new_n6484_;
  assign new_n20243_ = new_n16943_ & new_n16670_;
  assign new_n20244_ = ~new_n20243_ & new_n14388_;
  assign new_n20245_ = ~new_n20246_ & new_n15493_;
  assign new_n20246_ = ~new_n15445_ & ~new_n15469_;
  assign new_n20247_ = new_n7550_ & new_n7547_ & new_n7518_;
  assign new_n20248_ = new_n17154_ & new_n17176_;
  assign new_n20249_ = (~new_n20251_ | new_n20250_) & (~new_n20261_ | (new_n20262_ ? ~new_n20264_ : new_n15330_));
  assign new_n20250_ = ~new_n16479_ & (~new_n16456_ | new_n19426_);
  assign new_n20251_ = new_n20241_ & new_n20243_ & new_n9893_ & (new_n20257_ | ~new_n20252_);
  assign new_n20252_ = ~new_n9870_ & ~new_n20253_;
  assign new_n20253_ = ~new_n9892_ & ~new_n9891_ & (~new_n9894_ | (~new_n20254_ & ~new_n9872_ & ~new_n9878_));
  assign new_n20254_ = ~new_n9886_ & ~new_n9876_ & (~new_n9885_ | ~new_n9887_ | new_n20255_);
  assign new_n20255_ = new_n9880_ & new_n9882_ & (new_n20256_ | ~\all_features[4181]  | ~\all_features[4182]  | ~\all_features[4183] );
  assign new_n20256_ = ~\all_features[4179]  & ~\all_features[4180]  & (~\all_features[4178]  | new_n9874_);
  assign new_n20257_ = ~new_n20258_ & ~new_n9892_;
  assign new_n20258_ = ~new_n9891_ & (new_n9890_ | (~new_n9888_ & (new_n9878_ | (~new_n9872_ & ~new_n20259_))));
  assign new_n20259_ = ~new_n9876_ & (new_n9886_ | (new_n9885_ & (~new_n9887_ | (~new_n20260_ & new_n9880_))));
  assign new_n20260_ = ~\all_features[4181]  & \all_features[4182]  & \all_features[4183]  & (\all_features[4180]  ? new_n9884_ : (new_n9883_ | ~new_n9884_));
  assign new_n20261_ = ~new_n14388_ & ~new_n20243_;
  assign new_n20262_ = new_n13355_ & new_n20263_;
  assign new_n20263_ = ~new_n7137_ & ~new_n7159_;
  assign new_n20264_ = new_n20265_ & new_n12624_;
  assign new_n20265_ = new_n12601_ & new_n18169_;
  assign new_n20266_ = new_n20268_ & new_n20267_ & (~new_n20261_ | (new_n20264_ & new_n20262_) | (~new_n15330_ & ~new_n20262_));
  assign new_n20267_ = (~new_n20248_ | ~new_n20239_) & (~new_n20244_ | (new_n20245_ ? new_n20115_ : ~new_n20247_));
  assign new_n20268_ = (~new_n20250_ | ~new_n20251_) & (~new_n20240_ | ~new_n18786_);
  assign new_n20269_ = (new_n20306_ & ~new_n20439_ & (new_n20441_ | ~new_n20438_)) | (new_n20270_ & ~new_n20305_ & new_n20439_);
  assign new_n20270_ = (new_n13560_ | ~new_n20272_ | ~new_n20271_) & (new_n12535_ | ~new_n17812_ | new_n20271_);
  assign new_n20271_ = new_n11704_ & ~new_n18469_ & new_n18460_;
  assign new_n20272_ = new_n20303_ & (new_n20301_ | ~new_n20273_);
  assign new_n20273_ = ~new_n20274_ & (new_n20293_ | (~new_n20291_ & (new_n20296_ | new_n20298_)));
  assign new_n20274_ = new_n20290_ & (new_n20297_ | new_n20296_ | (~new_n20294_ & ~new_n20295_ & ~new_n20275_));
  assign new_n20275_ = ~new_n20287_ & ~new_n20285_ & (~new_n20276_ | (~new_n20289_ & new_n20280_));
  assign new_n20276_ = \all_features[1391]  & (\all_features[1390]  | (~new_n20277_ & \all_features[1389] ));
  assign new_n20277_ = new_n20278_ & ~\all_features[1388]  & new_n20279_;
  assign new_n20278_ = ~\all_features[1386]  & ~\all_features[1387] ;
  assign new_n20279_ = ~\all_features[1384]  & ~\all_features[1385] ;
  assign new_n20280_ = new_n20281_ & new_n20283_ & (new_n20284_ | \all_features[1388]  | \all_features[1389]  | ~new_n20278_);
  assign new_n20281_ = \all_features[1391]  & (\all_features[1390]  | (new_n20282_ & (\all_features[1386]  | \all_features[1387]  | \all_features[1385] )));
  assign new_n20282_ = \all_features[1388]  & \all_features[1389] ;
  assign new_n20283_ = \all_features[1390]  & \all_features[1391] ;
  assign new_n20284_ = \all_features[1384]  & \all_features[1385] ;
  assign new_n20285_ = ~new_n20286_ & ~\all_features[1391] ;
  assign new_n20286_ = \all_features[1389]  & \all_features[1390]  & (\all_features[1388]  | (\all_features[1386]  & \all_features[1387]  & \all_features[1385] ));
  assign new_n20287_ = ~\all_features[1391]  & (~\all_features[1390]  | ~new_n20282_ | ~new_n20284_ | ~new_n20288_);
  assign new_n20288_ = \all_features[1386]  & \all_features[1387] ;
  assign new_n20289_ = new_n20283_ & \all_features[1389]  & ((~new_n20279_ & \all_features[1386] ) | \all_features[1388]  | \all_features[1387] );
  assign new_n20290_ = ~new_n20291_ & ~new_n20293_;
  assign new_n20291_ = ~\all_features[1389]  & new_n20292_ & ((~\all_features[1386]  & new_n20279_) | ~\all_features[1388]  | ~\all_features[1387] );
  assign new_n20292_ = ~\all_features[1390]  & ~\all_features[1391] ;
  assign new_n20293_ = ~\all_features[1391]  & ~\all_features[1390]  & ~\all_features[1389]  & ~\all_features[1387]  & ~\all_features[1388] ;
  assign new_n20294_ = ~\all_features[1391]  & (~\all_features[1390]  | (~\all_features[1389]  & (new_n20279_ | ~new_n20288_ | ~\all_features[1388] )));
  assign new_n20295_ = ~\all_features[1391]  & (~\all_features[1390]  | (~\all_features[1388]  & ~\all_features[1389]  & ~new_n20288_));
  assign new_n20296_ = new_n20292_ & (~\all_features[1389]  | (~\all_features[1388]  & (~\all_features[1387]  | (~\all_features[1386]  & ~\all_features[1385] ))));
  assign new_n20297_ = new_n20292_ & (~\all_features[1387]  | ~new_n20282_ | (~\all_features[1386]  & ~new_n20284_));
  assign new_n20298_ = ~new_n20297_ & (new_n20295_ | (~new_n20294_ & (new_n20285_ | (~new_n20287_ & ~new_n20299_))));
  assign new_n20299_ = \all_features[1391]  & ((new_n20300_ & (\all_features[1390]  | \all_features[1389] )) | (~\all_features[1390]  & (\all_features[1389]  ? new_n20277_ : \all_features[1388] )));
  assign new_n20300_ = new_n20281_ & (\all_features[1389]  | ~new_n20283_ | (~new_n20284_ & ~\all_features[1388]  & new_n20278_) | (\all_features[1388]  & ~new_n20278_));
  assign new_n20301_ = new_n20290_ & ~new_n20297_ & ~new_n20302_ & ~new_n20296_;
  assign new_n20302_ = ~new_n20294_ & ~new_n20285_ & ~new_n20287_ & ~new_n20295_ & (~new_n20280_ | ~new_n20276_);
  assign new_n20303_ = new_n20304_ & new_n20290_ & ~new_n20285_ & ~new_n20296_;
  assign new_n20304_ = ~new_n20297_ & ~new_n20295_ & ~new_n20294_ & ~new_n20287_;
  assign new_n20305_ = new_n13560_ & new_n20271_;
  assign new_n20306_ = (new_n20341_ | ~new_n20375_ | new_n20309_) & (~new_n20307_ | ~new_n20309_ | (~new_n20436_ & ~new_n20407_));
  assign new_n20307_ = ~new_n11364_ & new_n20308_;
  assign new_n20308_ = new_n11339_ & new_n11361_;
  assign new_n20309_ = ~new_n20333_ & ~new_n20337_ & (~new_n20310_ | (~new_n20338_ & ~new_n20327_));
  assign new_n20310_ = new_n20311_ & (\all_features[1179]  | \all_features[1180]  | \all_features[1181]  | \all_features[1182]  | \all_features[1183] );
  assign new_n20311_ = new_n20326_ & (new_n20332_ | new_n20331_ | (~new_n20329_ & ~new_n20330_ & ~new_n20312_));
  assign new_n20312_ = ~new_n20323_ & ~new_n20321_ & (~new_n20325_ | new_n20316_ | ~new_n20313_);
  assign new_n20313_ = \all_features[1183]  & (\all_features[1182]  | new_n20314_);
  assign new_n20314_ = \all_features[1181]  & (\all_features[1178]  | \all_features[1179]  | \all_features[1180]  | ~new_n20315_);
  assign new_n20315_ = ~\all_features[1176]  & ~\all_features[1177] ;
  assign new_n20316_ = ~new_n20320_ & new_n20317_ & \all_features[1182]  & \all_features[1183]  & (~\all_features[1181]  | new_n20319_);
  assign new_n20317_ = \all_features[1183]  & (\all_features[1182]  | (new_n20318_ & (\all_features[1178]  | \all_features[1179]  | \all_features[1177] )));
  assign new_n20318_ = \all_features[1180]  & \all_features[1181] ;
  assign new_n20319_ = ~\all_features[1179]  & ~\all_features[1180]  & (~\all_features[1178]  | new_n20315_);
  assign new_n20320_ = ~\all_features[1178]  & ~\all_features[1179]  & ~\all_features[1180]  & ~\all_features[1181]  & (~\all_features[1177]  | ~\all_features[1176] );
  assign new_n20321_ = ~new_n20322_ & ~\all_features[1183] ;
  assign new_n20322_ = \all_features[1181]  & \all_features[1182]  & (\all_features[1180]  | (\all_features[1178]  & \all_features[1179]  & \all_features[1177] ));
  assign new_n20323_ = ~\all_features[1183]  & (~new_n20324_ | ~\all_features[1176]  | ~\all_features[1177]  | ~\all_features[1182]  | ~new_n20318_);
  assign new_n20324_ = \all_features[1178]  & \all_features[1179] ;
  assign new_n20325_ = \all_features[1183]  & (\all_features[1181]  | \all_features[1182]  | \all_features[1180] );
  assign new_n20326_ = ~new_n20327_ & (\all_features[1179]  | \all_features[1180]  | \all_features[1181]  | \all_features[1182]  | \all_features[1183] );
  assign new_n20327_ = ~\all_features[1181]  & new_n20328_ & ((~\all_features[1178]  & new_n20315_) | ~\all_features[1180]  | ~\all_features[1179] );
  assign new_n20328_ = ~\all_features[1182]  & ~\all_features[1183] ;
  assign new_n20329_ = ~\all_features[1183]  & (~\all_features[1182]  | (~\all_features[1181]  & (new_n20315_ | ~new_n20324_ | ~\all_features[1180] )));
  assign new_n20330_ = ~\all_features[1183]  & (~\all_features[1182]  | (~\all_features[1180]  & ~\all_features[1181]  & ~new_n20324_));
  assign new_n20331_ = new_n20328_ & (~\all_features[1181]  | (~\all_features[1180]  & (~\all_features[1179]  | (~\all_features[1178]  & ~\all_features[1177] ))));
  assign new_n20332_ = new_n20328_ & (~new_n20318_ | ~\all_features[1179]  | (~\all_features[1178]  & (~\all_features[1176]  | ~\all_features[1177] )));
  assign new_n20333_ = new_n20334_ & (~new_n20335_ | (new_n20336_ & new_n20325_ & new_n20313_ & new_n20317_));
  assign new_n20334_ = new_n20326_ & ~new_n20331_ & ~new_n20332_;
  assign new_n20335_ = ~new_n20330_ & ~new_n20323_ & ~new_n20329_ & ~new_n20321_;
  assign new_n20336_ = \all_features[1183]  & ~new_n20320_ & \all_features[1182] ;
  assign new_n20337_ = new_n20334_ & new_n20335_;
  assign new_n20338_ = ~new_n20331_ & (new_n20332_ | (~new_n20330_ & (new_n20329_ | (~new_n20321_ & ~new_n20339_))));
  assign new_n20339_ = ~new_n20323_ & (~new_n20325_ | (new_n20313_ & (~new_n20317_ | (~new_n20340_ & new_n20336_))));
  assign new_n20340_ = \all_features[1182]  & \all_features[1183]  & (\all_features[1181]  | (\all_features[1180]  & (\all_features[1179]  | \all_features[1178] )));
  assign new_n20341_ = ~new_n20371_ & new_n20342_;
  assign new_n20342_ = ~new_n20343_ & ~new_n20365_;
  assign new_n20343_ = ~new_n20344_ & ~new_n20364_;
  assign new_n20344_ = ~new_n20361_ & (new_n20359_ | (~new_n20362_ & (new_n20363_ | (~new_n20345_ & ~new_n20348_))));
  assign new_n20345_ = ~\all_features[2079]  & (~\all_features[2078]  | new_n20346_);
  assign new_n20346_ = ~\all_features[2077]  & (new_n20347_ | ~\all_features[2075]  | ~\all_features[2076]  | ~\all_features[2074] );
  assign new_n20347_ = ~\all_features[2072]  & ~\all_features[2073] ;
  assign new_n20348_ = ~new_n20353_ & (new_n20355_ | (new_n20358_ & (~new_n20349_ | (~new_n20357_ & new_n20351_))));
  assign new_n20349_ = \all_features[2079]  & (\all_features[2078]  | (\all_features[2077]  & (\all_features[2076]  | ~new_n20347_ | ~new_n20350_)));
  assign new_n20350_ = ~\all_features[2074]  & ~\all_features[2075] ;
  assign new_n20351_ = \all_features[2079]  & (\all_features[2078]  | (new_n20352_ & (\all_features[2074]  | \all_features[2075]  | \all_features[2073] )));
  assign new_n20352_ = \all_features[2076]  & \all_features[2077] ;
  assign new_n20353_ = ~new_n20354_ & ~\all_features[2079] ;
  assign new_n20354_ = \all_features[2077]  & \all_features[2078]  & (\all_features[2076]  | (\all_features[2074]  & \all_features[2075]  & \all_features[2073] ));
  assign new_n20355_ = ~\all_features[2079]  & (~new_n20356_ | ~\all_features[2074]  | ~\all_features[2075]  | ~\all_features[2078]  | ~new_n20352_);
  assign new_n20356_ = \all_features[2072]  & \all_features[2073] ;
  assign new_n20357_ = ~\all_features[2077]  & \all_features[2078]  & \all_features[2079]  & (\all_features[2076]  ? new_n20350_ : (new_n20356_ | ~new_n20350_));
  assign new_n20358_ = \all_features[2079]  & (\all_features[2077]  | \all_features[2078]  | \all_features[2076] );
  assign new_n20359_ = new_n20360_ & (~\all_features[2077]  | (~\all_features[2076]  & (~\all_features[2075]  | (~\all_features[2074]  & ~\all_features[2073] ))));
  assign new_n20360_ = ~\all_features[2078]  & ~\all_features[2079] ;
  assign new_n20361_ = ~\all_features[2077]  & new_n20360_ & ((~\all_features[2074]  & new_n20347_) | ~\all_features[2076]  | ~\all_features[2075] );
  assign new_n20362_ = new_n20360_ & (~\all_features[2075]  | ~new_n20352_ | (~\all_features[2074]  & ~new_n20356_));
  assign new_n20363_ = ~\all_features[2079]  & (~\all_features[2078]  | (~\all_features[2077]  & ~\all_features[2076]  & (~\all_features[2075]  | ~\all_features[2074] )));
  assign new_n20364_ = ~\all_features[2079]  & ~\all_features[2078]  & ~\all_features[2077]  & ~\all_features[2075]  & ~\all_features[2076] ;
  assign new_n20365_ = ~new_n20361_ & ~new_n20364_ & (~new_n20370_ | (~new_n20345_ & ~new_n20366_ & ~new_n20363_));
  assign new_n20366_ = ~new_n20355_ & ~new_n20353_ & (~new_n20358_ | ~new_n20349_ | new_n20367_);
  assign new_n20367_ = new_n20351_ & new_n20368_ & (new_n20369_ | ~\all_features[2077]  | ~\all_features[2078]  | ~\all_features[2079] );
  assign new_n20368_ = \all_features[2078]  & \all_features[2079]  & (\all_features[2076]  | \all_features[2077]  | new_n20356_ | ~new_n20350_);
  assign new_n20369_ = ~\all_features[2075]  & ~\all_features[2076]  & (~\all_features[2074]  | new_n20347_);
  assign new_n20370_ = ~new_n20359_ & ~new_n20362_;
  assign new_n20371_ = ~new_n20364_ & ~new_n20362_ & ~new_n20361_ & ~new_n20372_ & ~new_n20359_;
  assign new_n20372_ = ~new_n20345_ & ~new_n20355_ & new_n20374_ & (~new_n20349_ | ~new_n20373_);
  assign new_n20373_ = new_n20358_ & new_n20351_ & new_n20368_;
  assign new_n20374_ = ~new_n20353_ & ~new_n20363_;
  assign new_n20375_ = new_n20406_ & ~new_n20376_ & new_n20405_;
  assign new_n20376_ = ~new_n20377_ & ~new_n20402_;
  assign new_n20377_ = new_n20400_ & (~new_n20388_ | (new_n20392_ & (~new_n20396_ | new_n20378_)));
  assign new_n20378_ = new_n20379_ & (~new_n20382_ | (~new_n20387_ & \all_features[1853]  & \all_features[1854]  & \all_features[1855] ));
  assign new_n20379_ = \all_features[1855]  & (\all_features[1854]  | (~new_n20380_ & \all_features[1853] ));
  assign new_n20380_ = new_n20381_ & ~\all_features[1852]  & ~\all_features[1850]  & ~\all_features[1851] ;
  assign new_n20381_ = ~\all_features[1848]  & ~\all_features[1849] ;
  assign new_n20382_ = \all_features[1855]  & \all_features[1854]  & ~new_n20385_ & new_n20383_;
  assign new_n20383_ = \all_features[1855]  & (\all_features[1854]  | (new_n20384_ & (\all_features[1850]  | \all_features[1851]  | \all_features[1849] )));
  assign new_n20384_ = \all_features[1852]  & \all_features[1853] ;
  assign new_n20385_ = ~\all_features[1853]  & ~\all_features[1852]  & ~\all_features[1851]  & ~new_n20386_ & ~\all_features[1850] ;
  assign new_n20386_ = \all_features[1848]  & \all_features[1849] ;
  assign new_n20387_ = ~\all_features[1851]  & ~\all_features[1852]  & (~\all_features[1850]  | new_n20381_);
  assign new_n20388_ = ~new_n20389_ & ~new_n20390_;
  assign new_n20389_ = ~\all_features[1854]  & ~\all_features[1855]  & (~\all_features[1851]  | ~new_n20384_ | (~\all_features[1850]  & ~new_n20386_));
  assign new_n20390_ = ~\all_features[1855]  & ~new_n20391_ & ~\all_features[1854] ;
  assign new_n20391_ = \all_features[1853]  & (\all_features[1852]  | (\all_features[1851]  & (\all_features[1850]  | \all_features[1849] )));
  assign new_n20392_ = ~new_n20393_ & ~new_n20395_;
  assign new_n20393_ = ~\all_features[1855]  & (~\all_features[1854]  | (~\all_features[1852]  & ~\all_features[1853]  & ~new_n20394_));
  assign new_n20394_ = \all_features[1850]  & \all_features[1851] ;
  assign new_n20395_ = ~\all_features[1855]  & (~\all_features[1854]  | (~\all_features[1853]  & (new_n20381_ | ~new_n20394_ | ~\all_features[1852] )));
  assign new_n20396_ = ~new_n20397_ & ~new_n20398_;
  assign new_n20397_ = ~\all_features[1855]  & (~\all_features[1854]  | ~new_n20386_ | ~new_n20384_ | ~new_n20394_);
  assign new_n20398_ = ~new_n20399_ & ~\all_features[1855] ;
  assign new_n20399_ = \all_features[1853]  & \all_features[1854]  & (\all_features[1852]  | (\all_features[1850]  & \all_features[1851]  & \all_features[1849] ));
  assign new_n20400_ = ~new_n20401_ | (\all_features[1851]  & \all_features[1852]  & (\all_features[1850]  | ~new_n20381_));
  assign new_n20401_ = ~\all_features[1855]  & ~\all_features[1853]  & ~\all_features[1854] ;
  assign new_n20402_ = new_n20403_ & (new_n20395_ | new_n20398_ | ~new_n20404_ | (new_n20382_ & new_n20379_));
  assign new_n20403_ = new_n20388_ & new_n20400_;
  assign new_n20404_ = ~new_n20393_ & ~new_n20397_;
  assign new_n20405_ = new_n20396_ & new_n20403_ & new_n20392_;
  assign new_n20406_ = new_n20374_ & new_n20370_ & ~new_n20364_ & ~new_n20361_ & ~new_n20345_ & ~new_n20355_;
  assign new_n20407_ = new_n20408_ & new_n20431_;
  assign new_n20408_ = new_n20429_ & ~new_n20409_ & new_n20425_;
  assign new_n20409_ = new_n20410_ & (~new_n20423_ | ~new_n20424_ | ~new_n20420_ | ~new_n20422_);
  assign new_n20410_ = ~new_n20417_ & ~new_n20415_ & ~new_n20411_ & ~new_n20413_;
  assign new_n20411_ = ~\all_features[3879]  & (~\all_features[3878]  | (~\all_features[3876]  & ~\all_features[3877]  & ~new_n20412_));
  assign new_n20412_ = \all_features[3874]  & \all_features[3875] ;
  assign new_n20413_ = ~\all_features[3879]  & (~\all_features[3878]  | (~\all_features[3877]  & (new_n20414_ | ~\all_features[3876]  | ~new_n20412_)));
  assign new_n20414_ = ~\all_features[3872]  & ~\all_features[3873] ;
  assign new_n20415_ = ~new_n20416_ & ~\all_features[3879] ;
  assign new_n20416_ = \all_features[3877]  & \all_features[3878]  & (\all_features[3876]  | (\all_features[3874]  & \all_features[3875]  & \all_features[3873] ));
  assign new_n20417_ = ~\all_features[3879]  & (~\all_features[3878]  | ~new_n20412_ | ~new_n20418_ | ~new_n20419_);
  assign new_n20418_ = \all_features[3872]  & \all_features[3873] ;
  assign new_n20419_ = \all_features[3876]  & \all_features[3877] ;
  assign new_n20420_ = \all_features[3879]  & (\all_features[3878]  | (\all_features[3877]  & (\all_features[3876]  | ~new_n20421_ | ~new_n20414_)));
  assign new_n20421_ = ~\all_features[3874]  & ~\all_features[3875] ;
  assign new_n20422_ = \all_features[3879]  & (\all_features[3878]  | (new_n20419_ & (\all_features[3874]  | \all_features[3875]  | \all_features[3873] )));
  assign new_n20423_ = \all_features[3878]  & \all_features[3879]  & (\all_features[3876]  | \all_features[3877]  | new_n20418_ | ~new_n20421_);
  assign new_n20424_ = \all_features[3879]  & (\all_features[3877]  | \all_features[3878]  | \all_features[3876] );
  assign new_n20425_ = ~new_n20426_ & ~new_n20428_;
  assign new_n20426_ = new_n20427_ & (~\all_features[3875]  | ~new_n20419_ | (~\all_features[3874]  & ~new_n20418_));
  assign new_n20427_ = ~\all_features[3878]  & ~\all_features[3879] ;
  assign new_n20428_ = new_n20427_ & (~\all_features[3877]  | (~\all_features[3876]  & (~\all_features[3875]  | (~\all_features[3874]  & ~\all_features[3873] ))));
  assign new_n20429_ = ~new_n20430_ & (\all_features[3875]  | \all_features[3876]  | \all_features[3877]  | \all_features[3878]  | \all_features[3879] );
  assign new_n20430_ = ~\all_features[3877]  & new_n20427_ & ((~\all_features[3874]  & new_n20414_) | ~\all_features[3876]  | ~\all_features[3875] );
  assign new_n20431_ = new_n20429_ & (~new_n20425_ | (new_n20435_ & (new_n20432_ | new_n20415_ | new_n20417_)));
  assign new_n20432_ = new_n20420_ & new_n20424_ & (~new_n20423_ | ~new_n20422_ | new_n20433_);
  assign new_n20433_ = \all_features[3879]  & \all_features[3878]  & ~new_n20434_ & \all_features[3877] ;
  assign new_n20434_ = ~\all_features[3875]  & ~\all_features[3876]  & (~\all_features[3874]  | new_n20414_);
  assign new_n20435_ = ~new_n20411_ & ~new_n20413_;
  assign new_n20436_ = new_n20425_ & new_n20435_ & new_n20437_ & ~new_n20415_ & ~new_n20430_;
  assign new_n20437_ = ~new_n20417_ & (\all_features[3875]  | \all_features[3876]  | \all_features[3877]  | \all_features[3878]  | \all_features[3879] );
  assign new_n20438_ = ~new_n20307_ & new_n20309_;
  assign new_n20439_ = new_n8535_ & (new_n8533_ | ~new_n20440_);
  assign new_n20440_ = ~new_n8508_ & ~new_n18329_;
  assign new_n20441_ = ~new_n20442_ & new_n18961_;
  assign new_n20442_ = new_n20443_ & new_n20447_;
  assign new_n20443_ = ~new_n20444_ & (\all_features[2843]  | \all_features[2844]  | \all_features[2845]  | \all_features[2846]  | \all_features[2847] );
  assign new_n20444_ = ~new_n18981_ & (new_n18983_ | (~new_n18984_ & (new_n18974_ | (~new_n18978_ & ~new_n20445_))));
  assign new_n20445_ = ~new_n18972_ & (new_n18979_ | (new_n18970_ & (~new_n18976_ | (~new_n20446_ & new_n18965_))));
  assign new_n20446_ = ~\all_features[2845]  & \all_features[2846]  & \all_features[2847]  & (\all_features[2844]  ? new_n18968_ : (new_n18969_ | ~new_n18968_));
  assign new_n20447_ = new_n18980_ & (~new_n18986_ | (~new_n20448_ & ~new_n18974_ & ~new_n18978_));
  assign new_n20448_ = ~new_n18979_ & ~new_n18972_ & (~new_n18970_ | ~new_n18976_ | new_n20449_);
  assign new_n20449_ = new_n18965_ & new_n18967_ & (new_n20450_ | ~\all_features[2845]  | ~\all_features[2846]  | ~\all_features[2847] );
  assign new_n20450_ = ~\all_features[2843]  & ~\all_features[2844]  & (~\all_features[2842]  | new_n18977_);
  assign new_n20451_ = new_n20452_ ? (new_n20627_ ^ new_n20236_) : (~new_n20627_ ^ new_n20236_);
  assign new_n20452_ = new_n20453_ ? (new_n20490_ ^ new_n20574_) : (~new_n20490_ ^ new_n20574_);
  assign new_n20453_ = ~new_n20454_ & new_n20487_;
  assign new_n20454_ = new_n20455_ & ((~new_n15527_ & new_n20482_ & new_n20462_) | (new_n19499_ & new_n20457_));
  assign new_n20455_ = new_n20456_ & (~new_n20486_ | (new_n20485_ & new_n19821_) | (new_n18324_ & ~new_n19821_));
  assign new_n20456_ = (~new_n20457_ | new_n19499_) & (new_n15527_ | (new_n20482_ ? new_n20462_ : new_n20484_));
  assign new_n20457_ = new_n15527_ & ~new_n20458_ & new_n20460_;
  assign new_n20458_ = new_n20459_ & new_n20273_;
  assign new_n20459_ = ~new_n20301_ & ~new_n20303_;
  assign new_n20460_ = new_n19142_ & new_n20461_;
  assign new_n20461_ = ~new_n8447_ & ~new_n8475_;
  assign new_n20462_ = ~new_n11975_ & ~new_n20463_ & ~new_n11943_;
  assign new_n20463_ = new_n20464_ & new_n20473_;
  assign new_n20464_ = ~new_n20465_ & ~new_n15332_;
  assign new_n20465_ = ~new_n15345_ & ~new_n15341_ & ~new_n15337_ & ~new_n20466_ & ~new_n15347_;
  assign new_n20466_ = ~new_n15346_ & ~new_n15348_ & ~new_n15342_ & ~new_n15333_ & ~new_n20467_;
  assign new_n20467_ = new_n20472_ & new_n20471_ & new_n20468_ & new_n20470_;
  assign new_n20468_ = \all_features[5679]  & (\all_features[5678]  | (\all_features[5677]  & (\all_features[5676]  | ~new_n20469_ | ~new_n15335_)));
  assign new_n20469_ = ~\all_features[5674]  & ~\all_features[5675] ;
  assign new_n20470_ = \all_features[5679]  & (\all_features[5678]  | (new_n15340_ & (\all_features[5674]  | \all_features[5675]  | \all_features[5673] )));
  assign new_n20471_ = \all_features[5678]  & \all_features[5679]  & (\all_features[5676]  | \all_features[5677]  | new_n15339_ | ~new_n20469_);
  assign new_n20472_ = \all_features[5679]  & (\all_features[5677]  | \all_features[5678]  | \all_features[5676] );
  assign new_n20473_ = ~new_n20474_ & ~new_n20478_;
  assign new_n20474_ = ~new_n15345_ & ~new_n15347_ & (~new_n15336_ | (~new_n15333_ & ~new_n20475_ & ~new_n15346_));
  assign new_n20475_ = ~new_n15342_ & ~new_n15348_ & (~new_n20472_ | ~new_n20468_ | new_n20476_);
  assign new_n20476_ = new_n20470_ & new_n20471_ & (new_n20477_ | ~\all_features[5677]  | ~\all_features[5678]  | ~\all_features[5679] );
  assign new_n20477_ = ~\all_features[5675]  & ~\all_features[5676]  & (~\all_features[5674]  | new_n15335_);
  assign new_n20478_ = ~new_n20479_ & ~new_n15345_;
  assign new_n20479_ = ~new_n15347_ & (new_n15341_ | (~new_n15337_ & (new_n15346_ | (~new_n15333_ & ~new_n20480_))));
  assign new_n20480_ = ~new_n15342_ & (new_n15348_ | (new_n20472_ & (~new_n20468_ | (~new_n20481_ & new_n20470_))));
  assign new_n20481_ = ~\all_features[5677]  & \all_features[5678]  & \all_features[5679]  & (\all_features[5676]  ? new_n20469_ : (new_n15339_ | ~new_n20469_));
  assign new_n20482_ = new_n12626_ & new_n20483_;
  assign new_n20483_ = ~new_n12682_ & ~new_n12685_;
  assign new_n20484_ = new_n14528_ & (new_n14531_ | new_n14505_);
  assign new_n20485_ = ~new_n6388_ & (~new_n6385_ | new_n6355_);
  assign new_n20486_ = new_n20458_ & new_n15527_;
  assign new_n20487_ = new_n20488_ & (~new_n20486_ | (~new_n20485_ & new_n19821_) | (~new_n18324_ & ~new_n19821_));
  assign new_n20488_ = (new_n20460_ | new_n20458_ | ~new_n15527_) & (new_n20482_ | new_n20489_ | ~new_n20484_ | new_n15527_);
  assign new_n20489_ = new_n12600_ & ~new_n18165_ & ~new_n18169_;
  assign new_n20490_ = ~new_n20491_ & new_n20571_;
  assign new_n20491_ = ~new_n20534_ & new_n20492_ & (~new_n20569_ | (~new_n16810_ & new_n10248_) | (~new_n20570_ & ~new_n10248_));
  assign new_n20492_ = ~new_n20493_ & (~new_n20496_ | (~new_n20497_ & ~new_n20498_));
  assign new_n20493_ = new_n20495_ & new_n19147_ & ~new_n18119_ & ~new_n20494_;
  assign new_n20494_ = ~new_n20086_ & new_n18395_;
  assign new_n20495_ = new_n18893_ & (~new_n18895_ | ~new_n12784_);
  assign new_n20496_ = ~new_n19147_ & ~new_n20112_;
  assign new_n20497_ = ~new_n19717_ & new_n19843_;
  assign new_n20498_ = new_n19717_ & new_n20499_;
  assign new_n20499_ = new_n20533_ & (new_n20531_ | new_n20500_);
  assign new_n20500_ = ~new_n20530_ & new_n20519_ & (new_n20529_ | (~new_n20527_ & ~new_n20501_));
  assign new_n20501_ = ~new_n20514_ & (new_n20511_ | (~new_n20513_ & (new_n20516_ | (~new_n20502_ & ~new_n20518_))));
  assign new_n20502_ = ~new_n20503_ & \all_features[1831]  & (\all_features[1830]  | \all_features[1829]  | \all_features[1828] );
  assign new_n20503_ = \all_features[1831]  & ((~new_n20509_ & ~\all_features[1829]  & \all_features[1830] ) | (~new_n20507_ & (\all_features[1830]  | (~new_n20504_ & \all_features[1829] ))));
  assign new_n20504_ = new_n20505_ & ~\all_features[1828]  & new_n20506_;
  assign new_n20505_ = ~\all_features[1824]  & ~\all_features[1825] ;
  assign new_n20506_ = ~\all_features[1826]  & ~\all_features[1827] ;
  assign new_n20507_ = \all_features[1831]  & (\all_features[1830]  | (new_n20508_ & (\all_features[1826]  | \all_features[1827]  | \all_features[1825] )));
  assign new_n20508_ = \all_features[1828]  & \all_features[1829] ;
  assign new_n20509_ = (\all_features[1828]  & ~new_n20506_) | (~new_n20510_ & ~\all_features[1828]  & new_n20506_);
  assign new_n20510_ = \all_features[1824]  & \all_features[1825] ;
  assign new_n20511_ = ~\all_features[1831]  & (~\all_features[1830]  | (~\all_features[1828]  & ~\all_features[1829]  & ~new_n20512_));
  assign new_n20512_ = \all_features[1826]  & \all_features[1827] ;
  assign new_n20513_ = ~\all_features[1831]  & (~\all_features[1830]  | (~\all_features[1829]  & (new_n20505_ | ~\all_features[1828]  | ~new_n20512_)));
  assign new_n20514_ = new_n20515_ & (~\all_features[1827]  | ~new_n20508_ | (~\all_features[1826]  & ~new_n20510_));
  assign new_n20515_ = ~\all_features[1830]  & ~\all_features[1831] ;
  assign new_n20516_ = ~new_n20517_ & ~\all_features[1831] ;
  assign new_n20517_ = \all_features[1829]  & \all_features[1830]  & (\all_features[1828]  | (\all_features[1826]  & \all_features[1827]  & \all_features[1825] ));
  assign new_n20518_ = ~\all_features[1831]  & (~\all_features[1830]  | ~new_n20512_ | ~new_n20510_ | ~new_n20508_);
  assign new_n20519_ = new_n20528_ & (~new_n20526_ | (new_n20525_ & (new_n20520_ | new_n20516_ | new_n20518_)));
  assign new_n20520_ = new_n20521_ & (~new_n20522_ | (~new_n20524_ & \all_features[1829]  & \all_features[1830]  & \all_features[1831] ));
  assign new_n20521_ = \all_features[1831]  & (\all_features[1830]  | (~new_n20504_ & \all_features[1829] ));
  assign new_n20522_ = \all_features[1831]  & \all_features[1830]  & ~new_n20523_ & new_n20507_;
  assign new_n20523_ = new_n20506_ & ~\all_features[1829]  & ~new_n20510_ & ~\all_features[1828] ;
  assign new_n20524_ = ~\all_features[1827]  & ~\all_features[1828]  & (~\all_features[1826]  | new_n20505_);
  assign new_n20525_ = ~new_n20511_ & ~new_n20513_;
  assign new_n20526_ = ~new_n20527_ & ~new_n20514_;
  assign new_n20527_ = new_n20515_ & (~\all_features[1829]  | (~\all_features[1828]  & (~\all_features[1827]  | (~\all_features[1826]  & ~\all_features[1825] ))));
  assign new_n20528_ = ~new_n20529_ & ~new_n20530_;
  assign new_n20529_ = ~\all_features[1829]  & new_n20515_ & ((~\all_features[1826]  & new_n20505_) | ~\all_features[1828]  | ~\all_features[1827] );
  assign new_n20530_ = ~\all_features[1831]  & ~\all_features[1830]  & ~\all_features[1829]  & ~\all_features[1827]  & ~\all_features[1828] ;
  assign new_n20531_ = new_n20528_ & ~new_n20532_ & new_n20526_;
  assign new_n20532_ = ~new_n20511_ & ~new_n20513_ & ~new_n20516_ & ~new_n20518_ & (~new_n20522_ | ~new_n20521_);
  assign new_n20533_ = new_n20526_ & new_n20525_ & ~new_n20530_ & ~new_n20518_ & ~new_n20516_ & ~new_n20529_;
  assign new_n20534_ = new_n19147_ & (new_n18119_ ? (new_n20536_ ? ~new_n15282_ : ~new_n20535_) : new_n20494_);
  assign new_n20535_ = new_n10491_ & new_n10513_;
  assign new_n20536_ = ~new_n20537_ & new_n20564_;
  assign new_n20537_ = ~new_n20563_ & (~new_n20556_ | (~new_n20561_ & (new_n20554_ | new_n20562_ | ~new_n20538_)));
  assign new_n20538_ = ~new_n20550_ & ~new_n20548_ & ((~new_n20545_ & new_n20539_) | ~new_n20553_ | ~new_n20552_);
  assign new_n20539_ = \all_features[4743]  & \all_features[4742]  & ~new_n20542_ & new_n20540_;
  assign new_n20540_ = \all_features[4743]  & (\all_features[4742]  | (new_n20541_ & (\all_features[4738]  | \all_features[4739]  | \all_features[4737] )));
  assign new_n20541_ = \all_features[4740]  & \all_features[4741] ;
  assign new_n20542_ = new_n20544_ & ~\all_features[4741]  & ~new_n20543_ & ~\all_features[4740] ;
  assign new_n20543_ = \all_features[4736]  & \all_features[4737] ;
  assign new_n20544_ = ~\all_features[4738]  & ~\all_features[4739] ;
  assign new_n20545_ = \all_features[4743]  & \all_features[4742]  & ~new_n20546_ & \all_features[4741] ;
  assign new_n20546_ = ~\all_features[4739]  & ~\all_features[4740]  & (~\all_features[4738]  | new_n20547_);
  assign new_n20547_ = ~\all_features[4736]  & ~\all_features[4737] ;
  assign new_n20548_ = ~new_n20549_ & ~\all_features[4743] ;
  assign new_n20549_ = \all_features[4741]  & \all_features[4742]  & (\all_features[4740]  | (\all_features[4738]  & \all_features[4739]  & \all_features[4737] ));
  assign new_n20550_ = ~\all_features[4743]  & (~\all_features[4742]  | ~new_n20551_ | ~new_n20543_ | ~new_n20541_);
  assign new_n20551_ = \all_features[4738]  & \all_features[4739] ;
  assign new_n20552_ = \all_features[4743]  & (\all_features[4742]  | (\all_features[4741]  & (\all_features[4740]  | ~new_n20544_ | ~new_n20547_)));
  assign new_n20553_ = \all_features[4743]  & (\all_features[4741]  | \all_features[4742]  | \all_features[4740] );
  assign new_n20554_ = ~new_n20548_ & (new_n20550_ | (new_n20553_ & (~new_n20552_ | (~new_n20555_ & new_n20540_))));
  assign new_n20555_ = ~\all_features[4741]  & \all_features[4742]  & \all_features[4743]  & (\all_features[4740]  ? new_n20544_ : (new_n20543_ | ~new_n20544_));
  assign new_n20556_ = ~new_n20560_ & ~new_n20557_ & ~new_n20559_;
  assign new_n20557_ = new_n20558_ & (~\all_features[4741]  | (~\all_features[4740]  & (~\all_features[4739]  | (~\all_features[4738]  & ~\all_features[4737] ))));
  assign new_n20558_ = ~\all_features[4742]  & ~\all_features[4743] ;
  assign new_n20559_ = ~\all_features[4741]  & new_n20558_ & ((~\all_features[4738]  & new_n20547_) | ~\all_features[4740]  | ~\all_features[4739] );
  assign new_n20560_ = new_n20558_ & (~\all_features[4739]  | ~new_n20541_ | (~\all_features[4738]  & ~new_n20543_));
  assign new_n20561_ = ~\all_features[4743]  & (~\all_features[4742]  | (~\all_features[4740]  & ~\all_features[4741]  & ~new_n20551_));
  assign new_n20562_ = ~\all_features[4743]  & (~\all_features[4742]  | (~\all_features[4741]  & (new_n20547_ | ~\all_features[4740]  | ~new_n20551_)));
  assign new_n20563_ = ~\all_features[4743]  & ~\all_features[4742]  & ~\all_features[4741]  & ~\all_features[4739]  & ~\all_features[4740] ;
  assign new_n20564_ = new_n20557_ | ~new_n20567_ | ((new_n20548_ | ~new_n20568_) & (new_n20565_ | new_n20560_));
  assign new_n20565_ = new_n20566_ & (~new_n20539_ | ~new_n20552_ | ~new_n20553_);
  assign new_n20566_ = ~new_n20550_ & ~new_n20548_ & ~new_n20561_ & ~new_n20562_;
  assign new_n20567_ = ~new_n20559_ & ~new_n20563_;
  assign new_n20568_ = ~new_n20560_ & ~new_n20550_ & ~new_n20561_ & ~new_n20562_;
  assign new_n20569_ = ~new_n19147_ & new_n20112_;
  assign new_n20570_ = new_n8927_ & (new_n8924_ | new_n12733_);
  assign new_n20571_ = ~new_n20572_ & ~new_n20573_ & (new_n20498_ | new_n20497_ | ~new_n20496_);
  assign new_n20572_ = new_n20569_ & (new_n10248_ ? ~new_n16810_ : ~new_n20570_);
  assign new_n20573_ = new_n19147_ & ((new_n15282_ & new_n20536_ & new_n18119_) | (~new_n20494_ & ~new_n20495_ & ~new_n18119_));
  assign new_n20574_ = ~new_n20575_ & new_n20625_;
  assign new_n20575_ = new_n20576_ & (~new_n20585_ | ~new_n20583_ | (new_n20590_ ? new_n19412_ : ~new_n20589_));
  assign new_n20576_ = (new_n20585_ | ~new_n20586_ | ~new_n20583_) & (new_n20583_ | (new_n20588_ ? new_n20581_ : new_n20577_));
  assign new_n20577_ = ~new_n20578_ & new_n20579_;
  assign new_n20578_ = ~new_n16263_ & (~new_n16261_ | new_n18386_);
  assign new_n20579_ = ~new_n7475_ & (~new_n7477_ | new_n20580_);
  assign new_n20580_ = ~new_n7447_ & ~new_n7471_;
  assign new_n20581_ = ~new_n20582_ & ~new_n15034_;
  assign new_n20582_ = ~new_n13977_ & new_n17933_;
  assign new_n20583_ = ~new_n20584_ & new_n18396_;
  assign new_n20584_ = ~new_n19708_ & ~new_n18412_;
  assign new_n20585_ = ~new_n8471_ & new_n20461_;
  assign new_n20586_ = ~new_n20587_ & new_n20337_;
  assign new_n20587_ = ~new_n20333_ & ~new_n20311_;
  assign new_n20588_ = new_n16639_ & (new_n16613_ | new_n16640_ | new_n20151_);
  assign new_n20589_ = ~new_n14042_ & (~new_n14039_ | ~new_n16363_);
  assign new_n20590_ = ~new_n20623_ & ~new_n20612_ & ~new_n20620_ & (new_n20618_ | (~new_n20617_ & ~new_n20591_));
  assign new_n20591_ = ~new_n20605_ & (new_n20607_ | (~new_n20608_ & (new_n20609_ | (~new_n20592_ & ~new_n20610_))));
  assign new_n20592_ = ~new_n20599_ & (~new_n20603_ | (new_n20593_ & (~new_n20602_ | (~new_n20604_ & new_n20596_))));
  assign new_n20593_ = \all_features[1839]  & (\all_features[1838]  | new_n20594_);
  assign new_n20594_ = \all_features[1837]  & (\all_features[1834]  | \all_features[1835]  | \all_features[1836]  | ~new_n20595_);
  assign new_n20595_ = ~\all_features[1832]  & ~\all_features[1833] ;
  assign new_n20596_ = \all_features[1839]  & ~new_n20597_ & \all_features[1838] ;
  assign new_n20597_ = ~\all_features[1837]  & ~\all_features[1836]  & ~\all_features[1835]  & ~new_n20598_ & ~\all_features[1834] ;
  assign new_n20598_ = \all_features[1832]  & \all_features[1833] ;
  assign new_n20599_ = ~\all_features[1839]  & (~\all_features[1838]  | ~new_n20598_ | ~new_n20600_ | ~new_n20601_);
  assign new_n20600_ = \all_features[1836]  & \all_features[1837] ;
  assign new_n20601_ = \all_features[1834]  & \all_features[1835] ;
  assign new_n20602_ = \all_features[1839]  & (\all_features[1838]  | (new_n20600_ & (\all_features[1834]  | \all_features[1835]  | \all_features[1833] )));
  assign new_n20603_ = \all_features[1839]  & (\all_features[1837]  | \all_features[1838]  | \all_features[1836] );
  assign new_n20604_ = \all_features[1838]  & \all_features[1839]  & (\all_features[1837]  | (\all_features[1836]  & (\all_features[1835]  | \all_features[1834] )));
  assign new_n20605_ = new_n20606_ & (~\all_features[1837]  | (~\all_features[1836]  & (~\all_features[1835]  | (~\all_features[1834]  & ~\all_features[1833] ))));
  assign new_n20606_ = ~\all_features[1838]  & ~\all_features[1839] ;
  assign new_n20607_ = new_n20606_ & (~\all_features[1835]  | ~new_n20600_ | (~\all_features[1834]  & ~new_n20598_));
  assign new_n20608_ = ~\all_features[1839]  & (~\all_features[1838]  | (~\all_features[1836]  & ~\all_features[1837]  & ~new_n20601_));
  assign new_n20609_ = ~\all_features[1839]  & (~\all_features[1838]  | (~\all_features[1837]  & (new_n20595_ | ~new_n20601_ | ~\all_features[1836] )));
  assign new_n20610_ = ~new_n20611_ & ~\all_features[1839] ;
  assign new_n20611_ = \all_features[1837]  & \all_features[1838]  & (\all_features[1836]  | (\all_features[1834]  & \all_features[1835]  & \all_features[1833] ));
  assign new_n20612_ = new_n20616_ & (~new_n20619_ | (~new_n20613_ & ~new_n20608_ & ~new_n20609_));
  assign new_n20613_ = ~new_n20599_ & ~new_n20610_ & (~new_n20603_ | new_n20614_ | ~new_n20593_);
  assign new_n20614_ = ~new_n20597_ & new_n20602_ & \all_features[1838]  & \all_features[1839]  & (~\all_features[1837]  | new_n20615_);
  assign new_n20615_ = ~\all_features[1835]  & ~\all_features[1836]  & (~\all_features[1834]  | new_n20595_);
  assign new_n20616_ = ~new_n20617_ & ~new_n20618_;
  assign new_n20617_ = ~\all_features[1837]  & new_n20606_ & ((~\all_features[1834]  & new_n20595_) | ~\all_features[1836]  | ~\all_features[1835] );
  assign new_n20618_ = ~\all_features[1839]  & ~\all_features[1838]  & ~\all_features[1837]  & ~\all_features[1835]  & ~\all_features[1836] ;
  assign new_n20619_ = ~new_n20605_ & ~new_n20607_;
  assign new_n20620_ = new_n20619_ & ~new_n20621_ & new_n20616_;
  assign new_n20621_ = new_n20622_ & (~new_n20602_ | ~new_n20603_ | ~new_n20596_ | ~new_n20593_);
  assign new_n20622_ = ~new_n20599_ & ~new_n20610_ & ~new_n20608_ & ~new_n20609_;
  assign new_n20623_ = new_n20624_ & new_n20616_ & ~new_n20605_ & ~new_n20610_;
  assign new_n20624_ = ~new_n20599_ & ~new_n20609_ & ~new_n20607_ & ~new_n20608_;
  assign new_n20625_ = (new_n20626_ | ~new_n20583_) & (new_n20578_ | new_n20588_ | ~new_n20579_ | new_n20583_);
  assign new_n20626_ = (new_n20586_ | new_n20585_) & (~new_n20590_ | ~new_n19412_ | ~new_n20585_);
  assign new_n20627_ = new_n20628_ ^ new_n20779_;
  assign new_n20628_ = ~new_n20629_ & new_n20772_;
  assign new_n20629_ = new_n20630_ & (new_n20737_ | ~new_n20736_) & (~new_n20728_ | new_n20729_);
  assign new_n20630_ = (~new_n20661_ | ~new_n20631_) & (~new_n20634_ | (new_n19781_ ? ~new_n18099_ : new_n20695_));
  assign new_n20631_ = ~new_n20633_ & new_n20632_;
  assign new_n20632_ = ~new_n7601_ & ~new_n19598_;
  assign new_n20633_ = ~new_n10271_ & (~new_n10249_ | ~new_n19241_);
  assign new_n20634_ = new_n7601_ & new_n20635_;
  assign new_n20635_ = new_n20660_ | ~new_n20657_ | ((new_n20651_ | ~new_n20654_) & (new_n20636_ | new_n20655_));
  assign new_n20636_ = ~new_n20651_ & ~new_n20653_ & new_n20644_ & (~new_n20648_ | ~new_n20637_);
  assign new_n20637_ = new_n20643_ & new_n20638_ & new_n20641_;
  assign new_n20638_ = \all_features[5703]  & ~new_n20639_ & \all_features[5702] ;
  assign new_n20639_ = ~\all_features[5701]  & ~\all_features[5700]  & ~\all_features[5699]  & ~new_n20640_ & ~\all_features[5698] ;
  assign new_n20640_ = \all_features[5696]  & \all_features[5697] ;
  assign new_n20641_ = \all_features[5703]  & (\all_features[5702]  | (new_n20642_ & (\all_features[5698]  | \all_features[5699]  | \all_features[5697] )));
  assign new_n20642_ = \all_features[5700]  & \all_features[5701] ;
  assign new_n20643_ = \all_features[5703]  & (\all_features[5701]  | \all_features[5702]  | \all_features[5700] );
  assign new_n20644_ = ~new_n20645_ & ~new_n20647_;
  assign new_n20645_ = ~\all_features[5703]  & (~\all_features[5702]  | ~new_n20646_ | ~new_n20640_ | ~new_n20642_);
  assign new_n20646_ = \all_features[5698]  & \all_features[5699] ;
  assign new_n20647_ = ~\all_features[5703]  & (~\all_features[5702]  | (~\all_features[5700]  & ~\all_features[5701]  & ~new_n20646_));
  assign new_n20648_ = \all_features[5703]  & (\all_features[5702]  | new_n20649_);
  assign new_n20649_ = \all_features[5701]  & (\all_features[5698]  | \all_features[5699]  | \all_features[5700]  | ~new_n20650_);
  assign new_n20650_ = ~\all_features[5696]  & ~\all_features[5697] ;
  assign new_n20651_ = ~new_n20652_ & ~\all_features[5703] ;
  assign new_n20652_ = \all_features[5701]  & \all_features[5702]  & (\all_features[5700]  | (\all_features[5698]  & \all_features[5699]  & \all_features[5697] ));
  assign new_n20653_ = ~\all_features[5703]  & (~\all_features[5702]  | (~\all_features[5701]  & (new_n20650_ | ~new_n20646_ | ~\all_features[5700] )));
  assign new_n20654_ = new_n20644_ & ~new_n20653_ & ~new_n20655_;
  assign new_n20655_ = new_n20656_ & (~\all_features[5699]  | ~new_n20642_ | (~\all_features[5698]  & ~new_n20640_));
  assign new_n20656_ = ~\all_features[5702]  & ~\all_features[5703] ;
  assign new_n20657_ = ~new_n20658_ & ~new_n20659_;
  assign new_n20658_ = ~\all_features[5701]  & new_n20656_ & ((~\all_features[5698]  & new_n20650_) | ~\all_features[5700]  | ~\all_features[5699] );
  assign new_n20659_ = ~\all_features[5703]  & ~\all_features[5702]  & ~\all_features[5701]  & ~\all_features[5699]  & ~\all_features[5700] ;
  assign new_n20660_ = new_n20656_ & (~\all_features[5701]  | (~\all_features[5700]  & (~\all_features[5699]  | (~\all_features[5698]  & ~\all_features[5697] ))));
  assign new_n20661_ = ~new_n20693_ & (~new_n20662_ | (~new_n20684_ & ~new_n20689_));
  assign new_n20662_ = ~new_n20683_ & ~new_n20682_ & ~new_n20681_ & ~new_n20663_ & ~new_n20679_;
  assign new_n20663_ = ~new_n20678_ & ~new_n20677_ & ~new_n20675_ & ~new_n20664_ & ~new_n20667_;
  assign new_n20664_ = ~\all_features[2095]  & (~\all_features[2094]  | new_n20665_);
  assign new_n20665_ = ~\all_features[2093]  & (new_n20666_ | ~\all_features[2091]  | ~\all_features[2092]  | ~\all_features[2090] );
  assign new_n20666_ = ~\all_features[2088]  & ~\all_features[2089] ;
  assign new_n20667_ = new_n20674_ & new_n20672_ & new_n20668_ & new_n20670_;
  assign new_n20668_ = \all_features[2095]  & (\all_features[2094]  | (\all_features[2093]  & (\all_features[2092]  | ~new_n20669_ | ~new_n20666_)));
  assign new_n20669_ = ~\all_features[2090]  & ~\all_features[2091] ;
  assign new_n20670_ = \all_features[2095]  & (\all_features[2094]  | (new_n20671_ & (\all_features[2090]  | \all_features[2091]  | \all_features[2089] )));
  assign new_n20671_ = \all_features[2092]  & \all_features[2093] ;
  assign new_n20672_ = \all_features[2094]  & \all_features[2095]  & (\all_features[2092]  | \all_features[2093]  | new_n20673_ | ~new_n20669_);
  assign new_n20673_ = \all_features[2088]  & \all_features[2089] ;
  assign new_n20674_ = \all_features[2095]  & (\all_features[2093]  | \all_features[2094]  | \all_features[2092] );
  assign new_n20675_ = ~new_n20676_ & ~\all_features[2095] ;
  assign new_n20676_ = \all_features[2093]  & \all_features[2094]  & (\all_features[2092]  | (\all_features[2090]  & \all_features[2091]  & \all_features[2089] ));
  assign new_n20677_ = ~\all_features[2095]  & (~new_n20671_ | ~\all_features[2090]  | ~\all_features[2091]  | ~\all_features[2094]  | ~new_n20673_);
  assign new_n20678_ = ~\all_features[2095]  & (~\all_features[2094]  | (~\all_features[2093]  & ~\all_features[2092]  & (~\all_features[2091]  | ~\all_features[2090] )));
  assign new_n20679_ = ~\all_features[2093]  & new_n20680_ & ((~\all_features[2090]  & new_n20666_) | ~\all_features[2092]  | ~\all_features[2091] );
  assign new_n20680_ = ~\all_features[2094]  & ~\all_features[2095] ;
  assign new_n20681_ = new_n20680_ & (~\all_features[2091]  | ~new_n20671_ | (~\all_features[2090]  & ~new_n20673_));
  assign new_n20682_ = new_n20680_ & (~\all_features[2093]  | (~\all_features[2092]  & (~\all_features[2091]  | (~\all_features[2090]  & ~\all_features[2089] ))));
  assign new_n20683_ = ~\all_features[2095]  & ~\all_features[2094]  & ~\all_features[2093]  & ~\all_features[2091]  & ~\all_features[2092] ;
  assign new_n20684_ = ~new_n20683_ & ~new_n20679_ & (~new_n20688_ | (~new_n20685_ & ~new_n20664_ & ~new_n20678_));
  assign new_n20685_ = ~new_n20675_ & ~new_n20677_ & (~new_n20674_ | ~new_n20668_ | new_n20686_);
  assign new_n20686_ = new_n20670_ & new_n20672_ & (new_n20687_ | ~\all_features[2093]  | ~\all_features[2094]  | ~\all_features[2095] );
  assign new_n20687_ = ~\all_features[2091]  & ~\all_features[2092]  & (~\all_features[2090]  | new_n20666_);
  assign new_n20688_ = ~new_n20681_ & ~new_n20682_;
  assign new_n20689_ = ~new_n20690_ & ~new_n20683_;
  assign new_n20690_ = ~new_n20679_ & (new_n20682_ | (~new_n20681_ & (new_n20678_ | (~new_n20664_ & ~new_n20691_))));
  assign new_n20691_ = ~new_n20675_ & (new_n20677_ | (new_n20674_ & (~new_n20668_ | (~new_n20692_ & new_n20670_))));
  assign new_n20692_ = ~\all_features[2093]  & \all_features[2094]  & \all_features[2095]  & (\all_features[2092]  ? new_n20669_ : (new_n20673_ | ~new_n20669_));
  assign new_n20693_ = new_n20688_ & new_n20694_ & ~new_n20678_ & ~new_n20679_ & ~new_n20664_ & ~new_n20675_;
  assign new_n20694_ = ~new_n20677_ & ~new_n20683_;
  assign new_n20695_ = ~new_n20696_ & new_n20723_;
  assign new_n20696_ = ~new_n20722_ & (~new_n20715_ | (~new_n20720_ & (new_n20713_ | new_n20721_ | ~new_n20697_)));
  assign new_n20697_ = ~new_n20709_ & ~new_n20707_ & ((~new_n20704_ & new_n20698_) | ~new_n20712_ | ~new_n20711_);
  assign new_n20698_ = \all_features[1615]  & \all_features[1614]  & ~new_n20701_ & new_n20699_;
  assign new_n20699_ = \all_features[1615]  & (\all_features[1614]  | (new_n20700_ & (\all_features[1610]  | \all_features[1611]  | \all_features[1609] )));
  assign new_n20700_ = \all_features[1612]  & \all_features[1613] ;
  assign new_n20701_ = new_n20703_ & ~\all_features[1613]  & ~new_n20702_ & ~\all_features[1612] ;
  assign new_n20702_ = \all_features[1608]  & \all_features[1609] ;
  assign new_n20703_ = ~\all_features[1610]  & ~\all_features[1611] ;
  assign new_n20704_ = \all_features[1615]  & \all_features[1614]  & ~new_n20705_ & \all_features[1613] ;
  assign new_n20705_ = ~\all_features[1611]  & ~\all_features[1612]  & (~\all_features[1610]  | new_n20706_);
  assign new_n20706_ = ~\all_features[1608]  & ~\all_features[1609] ;
  assign new_n20707_ = ~new_n20708_ & ~\all_features[1615] ;
  assign new_n20708_ = \all_features[1613]  & \all_features[1614]  & (\all_features[1612]  | (\all_features[1610]  & \all_features[1611]  & \all_features[1609] ));
  assign new_n20709_ = ~\all_features[1615]  & (~\all_features[1614]  | ~new_n20710_ | ~new_n20702_ | ~new_n20700_);
  assign new_n20710_ = \all_features[1610]  & \all_features[1611] ;
  assign new_n20711_ = \all_features[1615]  & (\all_features[1614]  | (\all_features[1613]  & (\all_features[1612]  | ~new_n20703_ | ~new_n20706_)));
  assign new_n20712_ = \all_features[1615]  & (\all_features[1613]  | \all_features[1614]  | \all_features[1612] );
  assign new_n20713_ = ~new_n20707_ & (new_n20709_ | (new_n20712_ & (~new_n20711_ | (~new_n20714_ & new_n20699_))));
  assign new_n20714_ = ~\all_features[1613]  & \all_features[1614]  & \all_features[1615]  & (\all_features[1612]  ? new_n20703_ : (new_n20702_ | ~new_n20703_));
  assign new_n20715_ = ~new_n20719_ & ~new_n20716_ & ~new_n20718_;
  assign new_n20716_ = new_n20717_ & (~\all_features[1613]  | (~\all_features[1612]  & (~\all_features[1611]  | (~\all_features[1610]  & ~\all_features[1609] ))));
  assign new_n20717_ = ~\all_features[1614]  & ~\all_features[1615] ;
  assign new_n20718_ = ~\all_features[1613]  & new_n20717_ & ((~\all_features[1610]  & new_n20706_) | ~\all_features[1612]  | ~\all_features[1611] );
  assign new_n20719_ = new_n20717_ & (~\all_features[1611]  | ~new_n20700_ | (~\all_features[1610]  & ~new_n20702_));
  assign new_n20720_ = ~\all_features[1615]  & (~\all_features[1614]  | (~\all_features[1612]  & ~\all_features[1613]  & ~new_n20710_));
  assign new_n20721_ = ~\all_features[1615]  & (~\all_features[1614]  | (~\all_features[1613]  & (new_n20706_ | ~\all_features[1612]  | ~new_n20710_)));
  assign new_n20722_ = ~\all_features[1615]  & ~\all_features[1614]  & ~\all_features[1613]  & ~\all_features[1611]  & ~\all_features[1612] ;
  assign new_n20723_ = new_n20716_ | ~new_n20726_ | ((new_n20707_ | ~new_n20727_) & (new_n20724_ | new_n20719_));
  assign new_n20724_ = new_n20725_ & (~new_n20698_ | ~new_n20711_ | ~new_n20712_);
  assign new_n20725_ = ~new_n20709_ & ~new_n20707_ & ~new_n20720_ & ~new_n20721_;
  assign new_n20726_ = ~new_n20718_ & ~new_n20722_;
  assign new_n20727_ = ~new_n20719_ & ~new_n20709_ & ~new_n20720_ & ~new_n20721_;
  assign new_n20728_ = new_n20632_ & new_n20633_;
  assign new_n20729_ = ~new_n14947_ & (~new_n14924_ | ~new_n20730_);
  assign new_n20730_ = new_n20731_ & new_n14950_;
  assign new_n20731_ = (new_n20732_ | (new_n14934_ & (~\all_features[2331]  | ~\all_features[2332]  | (~\all_features[2330]  & new_n14933_)))) & (~new_n14934_ | \all_features[2331]  | \all_features[2332] );
  assign new_n20732_ = ~new_n14930_ & (new_n14927_ | (~new_n14941_ & (new_n14944_ | (~new_n20733_ & ~new_n14945_))));
  assign new_n20733_ = ~new_n14943_ & (~\all_features[2335]  | new_n20734_ | (~\all_features[2332]  & ~\all_features[2333]  & ~\all_features[2334] ));
  assign new_n20734_ = \all_features[2335]  & ((~new_n20735_ & ~\all_features[2333]  & \all_features[2334] ) | (~new_n14938_ & (\all_features[2334]  | (~new_n14936_ & \all_features[2333] ))));
  assign new_n20735_ = (\all_features[2332]  & (\all_features[2330]  | \all_features[2331] )) | (~new_n14928_ & ~\all_features[2330]  & ~\all_features[2331]  & ~\all_features[2332] );
  assign new_n20736_ = ~new_n7601_ & new_n19598_;
  assign new_n20737_ = (~new_n19433_ | (~new_n20768_ & new_n20738_)) & (new_n16712_ | new_n16744_ | ~new_n18042_ | new_n19433_);
  assign new_n20738_ = ~new_n20767_ & ~new_n20739_ & ~new_n20761_;
  assign new_n20739_ = new_n20756_ & ~new_n20760_ & ~new_n20740_ & ~new_n20759_;
  assign new_n20740_ = new_n20741_ & ~new_n20749_ & (~new_n20754_ | ~new_n20755_ | ~new_n20751_ | ~new_n20753_);
  assign new_n20741_ = ~new_n20746_ & ~new_n20742_ & ~new_n20744_;
  assign new_n20742_ = ~\all_features[5199]  & (~\all_features[5198]  | (~\all_features[5196]  & ~\all_features[5197]  & ~new_n20743_));
  assign new_n20743_ = \all_features[5194]  & \all_features[5195] ;
  assign new_n20744_ = ~new_n20745_ & ~\all_features[5199] ;
  assign new_n20745_ = \all_features[5197]  & \all_features[5198]  & (\all_features[5196]  | (\all_features[5194]  & \all_features[5195]  & \all_features[5193] ));
  assign new_n20746_ = ~\all_features[5199]  & (~\all_features[5198]  | ~new_n20747_ | ~new_n20748_ | ~new_n20743_);
  assign new_n20747_ = \all_features[5192]  & \all_features[5193] ;
  assign new_n20748_ = \all_features[5196]  & \all_features[5197] ;
  assign new_n20749_ = ~\all_features[5199]  & (~\all_features[5198]  | (~\all_features[5197]  & (new_n20750_ | ~new_n20743_ | ~\all_features[5196] )));
  assign new_n20750_ = ~\all_features[5192]  & ~\all_features[5193] ;
  assign new_n20751_ = \all_features[5199]  & (\all_features[5198]  | (\all_features[5197]  & (\all_features[5196]  | ~new_n20752_ | ~new_n20750_)));
  assign new_n20752_ = ~\all_features[5194]  & ~\all_features[5195] ;
  assign new_n20753_ = \all_features[5199]  & (\all_features[5198]  | (new_n20748_ & (\all_features[5194]  | \all_features[5195]  | \all_features[5193] )));
  assign new_n20754_ = \all_features[5198]  & \all_features[5199]  & (\all_features[5196]  | \all_features[5197]  | new_n20747_ | ~new_n20752_);
  assign new_n20755_ = \all_features[5199]  & (\all_features[5197]  | \all_features[5198]  | \all_features[5196] );
  assign new_n20756_ = ~new_n20757_ & (\all_features[5195]  | \all_features[5196]  | \all_features[5197]  | \all_features[5198]  | \all_features[5199] );
  assign new_n20757_ = new_n20758_ & (~\all_features[5195]  | ~new_n20748_ | (~\all_features[5194]  & ~new_n20747_));
  assign new_n20758_ = ~\all_features[5198]  & ~\all_features[5199] ;
  assign new_n20759_ = ~\all_features[5197]  & new_n20758_ & ((~\all_features[5194]  & new_n20750_) | ~\all_features[5196]  | ~\all_features[5195] );
  assign new_n20760_ = new_n20758_ & (~\all_features[5197]  | (~\all_features[5196]  & (~\all_features[5195]  | (~\all_features[5194]  & ~\all_features[5193] ))));
  assign new_n20761_ = new_n20765_ & (~new_n20766_ | (~new_n20762_ & ~new_n20742_ & ~new_n20749_));
  assign new_n20762_ = ~new_n20744_ & ~new_n20746_ & (~new_n20755_ | ~new_n20751_ | new_n20763_);
  assign new_n20763_ = new_n20753_ & new_n20754_ & (new_n20764_ | ~\all_features[5197]  | ~\all_features[5198]  | ~\all_features[5199] );
  assign new_n20764_ = ~\all_features[5195]  & ~\all_features[5196]  & (~\all_features[5194]  | new_n20750_);
  assign new_n20765_ = ~new_n20759_ & (\all_features[5195]  | \all_features[5196]  | \all_features[5197]  | \all_features[5198]  | \all_features[5199] );
  assign new_n20766_ = ~new_n20760_ & ~new_n20757_;
  assign new_n20767_ = new_n20741_ & new_n20766_ & ~new_n20749_ & new_n20765_;
  assign new_n20768_ = ~new_n20769_ & (\all_features[5195]  | \all_features[5196]  | \all_features[5197]  | \all_features[5198]  | \all_features[5199] );
  assign new_n20769_ = ~new_n20759_ & (new_n20760_ | (~new_n20757_ & (new_n20742_ | (~new_n20770_ & ~new_n20749_))));
  assign new_n20770_ = ~new_n20744_ & (new_n20746_ | (new_n20755_ & (~new_n20751_ | (~new_n20771_ & new_n20753_))));
  assign new_n20771_ = ~\all_features[5197]  & \all_features[5198]  & \all_features[5199]  & (\all_features[5196]  ? new_n20752_ : (new_n20747_ | ~new_n20752_));
  assign new_n20772_ = new_n20773_ & (new_n20661_ | ~new_n20631_) & (new_n20775_ | new_n20777_ | ~new_n20774_);
  assign new_n20773_ = (~new_n20737_ | ~new_n20736_) & (~new_n20634_ | (new_n19781_ ? new_n18099_ : ~new_n20695_));
  assign new_n20774_ = ~new_n20635_ & new_n7601_;
  assign new_n20775_ = new_n9893_ & new_n20776_ & new_n9870_;
  assign new_n20776_ = new_n20257_ & new_n20253_;
  assign new_n20777_ = ~new_n20778_ & new_n16777_;
  assign new_n20778_ = new_n16806_ & new_n16802_;
  assign new_n20779_ = new_n20780_ & (new_n20796_ | (~new_n20795_ & (~new_n20804_ | ~new_n20802_)));
  assign new_n20780_ = new_n20782_ & (new_n20789_ | new_n20794_ | ~new_n20781_);
  assign new_n20781_ = ~new_n7556_ & new_n6532_;
  assign new_n20782_ = new_n6532_ | (new_n20788_ ? (new_n16957_ ? new_n20786_ : ~new_n20787_) : new_n20783_);
  assign new_n20783_ = new_n7443_ & new_n20784_;
  assign new_n20784_ = new_n19457_ & (new_n19435_ | new_n20785_);
  assign new_n20785_ = new_n19459_ & new_n19463_;
  assign new_n20786_ = new_n13209_ & new_n19836_;
  assign new_n20787_ = ~new_n20274_ & new_n20459_;
  assign new_n20788_ = new_n8202_ & new_n8225_;
  assign new_n20789_ = ~new_n12082_ & (~new_n20119_ | (new_n20790_ & new_n20143_));
  assign new_n20790_ = ~new_n20791_ & (\all_features[4291]  | \all_features[4292]  | \all_features[4293]  | \all_features[4294]  | \all_features[4295] );
  assign new_n20791_ = ~new_n20141_ & (new_n20142_ | (~new_n20129_ & (new_n20126_ | (~new_n20127_ & ~new_n20792_))));
  assign new_n20792_ = ~new_n20137_ & (new_n20122_ | (new_n20136_ & (~new_n20139_ | (~new_n20793_ & new_n20133_))));
  assign new_n20793_ = ~\all_features[4293]  & \all_features[4294]  & \all_features[4295]  & (\all_features[4292]  ? new_n20135_ : (new_n20124_ | ~new_n20135_));
  assign new_n20794_ = new_n12082_ & new_n16282_;
  assign new_n20795_ = new_n20781_ & new_n20789_;
  assign new_n20796_ = new_n7556_ & new_n6532_ & (new_n20797_ ? ~new_n20800_ : ~new_n20799_);
  assign new_n20797_ = ~new_n20798_ & new_n17676_;
  assign new_n20798_ = new_n17701_ & new_n17705_;
  assign new_n20799_ = new_n16958_ & (~new_n16959_ | ~new_n16054_);
  assign new_n20800_ = ~new_n20801_ & new_n13169_;
  assign new_n20801_ = new_n13197_ & new_n13978_;
  assign new_n20802_ = ~new_n20803_ & (~new_n6532_ | ((new_n20797_ | ~new_n20799_ | ~new_n7556_) & (~new_n20794_ | new_n7556_)));
  assign new_n20803_ = new_n16957_ & new_n20788_ & ~new_n6532_ & new_n20786_;
  assign new_n20804_ = ~new_n6532_ & ((new_n7443_ & new_n20784_ & ~new_n20788_) | (~new_n16957_ & ~new_n20787_ & new_n20788_));
  assign new_n20805_ = new_n20806_ & new_n20867_;
  assign new_n20806_ = ~new_n20809_ & (~new_n20844_ | (new_n20807_ & new_n20851_) | (~new_n20845_ & ~new_n20852_ & ~new_n20851_));
  assign new_n20807_ = ~new_n18385_ & new_n20808_;
  assign new_n20808_ = ~new_n8739_ & (~new_n8736_ | ~new_n8704_);
  assign new_n20809_ = ~new_n14293_ & ~new_n20844_ & (new_n16777_ ? new_n20843_ : new_n20810_);
  assign new_n20810_ = new_n20811_ & new_n20842_;
  assign new_n20811_ = new_n20812_ & new_n20838_;
  assign new_n20812_ = ~new_n20813_ & (\all_features[5219]  | \all_features[5220]  | \all_features[5221]  | \all_features[5222]  | \all_features[5223] );
  assign new_n20813_ = new_n20831_ & (new_n20837_ | (~new_n20836_ & new_n20814_ & (new_n20823_ | new_n20829_)));
  assign new_n20814_ = ~new_n20823_ & ~new_n20825_ & (~new_n20828_ | ~new_n20827_ | new_n20815_);
  assign new_n20815_ = new_n20816_ & ~new_n20821_ & new_n20818_;
  assign new_n20816_ = \all_features[5223]  & (\all_features[5222]  | (new_n20817_ & (\all_features[5218]  | \all_features[5219]  | \all_features[5217] )));
  assign new_n20817_ = \all_features[5220]  & \all_features[5221] ;
  assign new_n20818_ = new_n20820_ & (\all_features[5220]  | \all_features[5221]  | ~new_n20819_ | (\all_features[5217]  & \all_features[5216] ));
  assign new_n20819_ = ~\all_features[5218]  & ~\all_features[5219] ;
  assign new_n20820_ = \all_features[5222]  & \all_features[5223] ;
  assign new_n20821_ = new_n20820_ & \all_features[5221]  & ((~new_n20822_ & \all_features[5218] ) | \all_features[5220]  | \all_features[5219] );
  assign new_n20822_ = ~\all_features[5216]  & ~\all_features[5217] ;
  assign new_n20823_ = ~new_n20824_ & ~\all_features[5223] ;
  assign new_n20824_ = \all_features[5221]  & \all_features[5222]  & (\all_features[5220]  | (\all_features[5218]  & \all_features[5219]  & \all_features[5217] ));
  assign new_n20825_ = ~\all_features[5223]  & (~new_n20817_ | ~\all_features[5216]  | ~\all_features[5217]  | ~\all_features[5222]  | ~new_n20826_);
  assign new_n20826_ = \all_features[5218]  & \all_features[5219] ;
  assign new_n20827_ = \all_features[5223]  & (\all_features[5222]  | (\all_features[5221]  & (\all_features[5220]  | ~new_n20819_ | ~new_n20822_)));
  assign new_n20828_ = \all_features[5223]  & (\all_features[5221]  | \all_features[5222]  | \all_features[5220] );
  assign new_n20829_ = ~new_n20825_ & (~new_n20828_ | (new_n20827_ & (~new_n20816_ | (~new_n20830_ & new_n20818_))));
  assign new_n20830_ = new_n20820_ & (\all_features[5221]  | (~new_n20819_ & \all_features[5220] ));
  assign new_n20831_ = ~new_n20835_ & ~new_n20832_ & ~new_n20834_;
  assign new_n20832_ = new_n20833_ & (~\all_features[5221]  | (~\all_features[5220]  & (~\all_features[5219]  | (~\all_features[5218]  & ~\all_features[5217] ))));
  assign new_n20833_ = ~\all_features[5222]  & ~\all_features[5223] ;
  assign new_n20834_ = new_n20833_ & (~new_n20817_ | ~\all_features[5219]  | (~\all_features[5218]  & (~\all_features[5216]  | ~\all_features[5217] )));
  assign new_n20835_ = ~\all_features[5221]  & new_n20833_ & ((~\all_features[5218]  & new_n20822_) | ~\all_features[5220]  | ~\all_features[5219] );
  assign new_n20836_ = ~\all_features[5223]  & (~\all_features[5222]  | (~\all_features[5221]  & (new_n20822_ | ~\all_features[5220]  | ~new_n20826_)));
  assign new_n20837_ = ~\all_features[5223]  & (~\all_features[5222]  | (~\all_features[5220]  & ~\all_features[5221]  & ~new_n20826_));
  assign new_n20838_ = new_n20839_ & (~new_n20841_ | (new_n20818_ & new_n20828_ & new_n20827_ & new_n20816_));
  assign new_n20839_ = new_n20840_ & ~new_n20832_ & ~new_n20834_;
  assign new_n20840_ = ~new_n20835_ & (\all_features[5219]  | \all_features[5220]  | \all_features[5221]  | \all_features[5222]  | \all_features[5223] );
  assign new_n20841_ = ~new_n20837_ & ~new_n20825_ & ~new_n20836_ & ~new_n20823_;
  assign new_n20842_ = new_n20839_ & new_n20841_;
  assign new_n20843_ = ~new_n19650_ & ~new_n19677_;
  assign new_n20844_ = ~new_n11201_ & (~new_n11199_ | ~new_n11173_);
  assign new_n20845_ = ~new_n19766_ & (~new_n19764_ | new_n20846_);
  assign new_n20846_ = ~new_n19738_ & (new_n19760_ | (~new_n19759_ & (new_n19757_ | new_n20847_)));
  assign new_n20847_ = ~new_n19755_ & (new_n19751_ | (~new_n19753_ & (new_n19761_ | (~new_n20848_ & ~new_n19763_))));
  assign new_n20848_ = ~new_n20849_ & \all_features[4359]  & (\all_features[4358]  | \all_features[4357]  | \all_features[4356] );
  assign new_n20849_ = \all_features[4359]  & ((~new_n20850_ & ~\all_features[4357]  & \all_features[4358] ) | (~new_n19745_ & (\all_features[4358]  | (~new_n19741_ & \all_features[4357] ))));
  assign new_n20850_ = (\all_features[4356]  & ~new_n19743_) | (~new_n19748_ & ~\all_features[4356]  & new_n19743_);
  assign new_n20851_ = new_n11361_ & (new_n11365_ | new_n11339_);
  assign new_n20852_ = new_n20853_ & ~new_n20866_ & ~new_n20865_ & ~new_n20862_ & ~new_n20864_;
  assign new_n20853_ = ~new_n20861_ & ~new_n20860_ & ~new_n20854_ & ~new_n20857_;
  assign new_n20854_ = ~\all_features[3527]  & (~\all_features[3526]  | (~\all_features[3525]  & (new_n20856_ | ~\all_features[3524]  | ~new_n20855_)));
  assign new_n20855_ = \all_features[3522]  & \all_features[3523] ;
  assign new_n20856_ = ~\all_features[3520]  & ~\all_features[3521] ;
  assign new_n20857_ = new_n20858_ & (~new_n20859_ | ~\all_features[3523]  | (~\all_features[3522]  & (~\all_features[3520]  | ~\all_features[3521] )));
  assign new_n20858_ = ~\all_features[3526]  & ~\all_features[3527] ;
  assign new_n20859_ = \all_features[3524]  & \all_features[3525] ;
  assign new_n20860_ = ~\all_features[3525]  & new_n20858_ & ((~\all_features[3522]  & new_n20856_) | ~\all_features[3524]  | ~\all_features[3523] );
  assign new_n20861_ = ~\all_features[3527]  & (~\all_features[3526]  | (~\all_features[3524]  & ~\all_features[3525]  & ~new_n20855_));
  assign new_n20862_ = ~new_n20863_ & ~\all_features[3527] ;
  assign new_n20863_ = \all_features[3525]  & \all_features[3526]  & (\all_features[3524]  | (\all_features[3522]  & \all_features[3523]  & \all_features[3521] ));
  assign new_n20864_ = new_n20858_ & (~\all_features[3525]  | (~\all_features[3524]  & (~\all_features[3523]  | (~\all_features[3522]  & ~\all_features[3521] ))));
  assign new_n20865_ = ~\all_features[3527]  & (~new_n20859_ | ~\all_features[3520]  | ~\all_features[3521]  | ~\all_features[3526]  | ~new_n20855_);
  assign new_n20866_ = ~\all_features[3527]  & ~\all_features[3526]  & ~\all_features[3525]  & ~\all_features[3523]  & ~\all_features[3524] ;
  assign new_n20867_ = new_n20844_ ? new_n20868_ : (new_n14293_ ? new_n20869_ : ~new_n20872_);
  assign new_n20868_ = (new_n18385_ | ~new_n20808_ | ~new_n20851_) & (new_n20845_ | new_n20852_ | new_n20851_);
  assign new_n20869_ = new_n9787_ & new_n9763_ & ~new_n9789_ & new_n20870_;
  assign new_n20870_ = new_n7700_ & new_n20871_;
  assign new_n20871_ = ~new_n7733_ & ~new_n7736_;
  assign new_n20872_ = new_n16777_ ? ~new_n20843_ : ~new_n20810_;
  assign new_n20873_ = new_n20874_ ? (~new_n20805_ ^ new_n21348_) : (new_n20805_ ^ new_n21348_);
  assign new_n20874_ = new_n20875_ ? (~new_n21184_ ^ new_n21347_) : (new_n21184_ ^ new_n21347_);
  assign new_n20875_ = new_n20876_ ? (~new_n20961_ ^ new_n21052_) : (new_n20961_ ^ new_n21052_);
  assign new_n20876_ = new_n20877_ & new_n20889_;
  assign new_n20877_ = (~new_n20878_ | new_n20887_) & (~new_n20885_ | (new_n11614_ ? new_n14618_ : new_n20888_));
  assign new_n20878_ = ~new_n20884_ & new_n20879_;
  assign new_n20879_ = ~new_n20880_ & new_n20882_;
  assign new_n20880_ = ~new_n8631_ & new_n20881_;
  assign new_n20881_ = ~new_n8663_ & ~new_n8666_;
  assign new_n20882_ = new_n18008_ & new_n20883_;
  assign new_n20883_ = ~new_n13480_ & ~new_n13503_;
  assign new_n20884_ = ~new_n16639_ & (~new_n16613_ | ~new_n16640_);
  assign new_n20885_ = ~new_n20886_ & new_n20880_;
  assign new_n20886_ = new_n12115_ & (new_n12112_ | new_n12084_);
  assign new_n20887_ = ~new_n19315_ & new_n11860_;
  assign new_n20888_ = new_n16613_ & new_n16639_;
  assign new_n20889_ = (new_n20958_ | ~new_n20890_) & (new_n20894_ | ~new_n20893_) & (~new_n20892_ | ~new_n20960_);
  assign new_n20890_ = new_n20891_ & new_n19340_;
  assign new_n20891_ = new_n20880_ & new_n20886_;
  assign new_n20892_ = new_n20879_ & new_n20884_;
  assign new_n20893_ = ~new_n20880_ & ~new_n20882_;
  assign new_n20894_ = (new_n20895_ & ~new_n20923_) | (~new_n10877_ & new_n20957_ & new_n20923_);
  assign new_n20895_ = new_n20896_ & new_n20921_;
  assign new_n20896_ = new_n20915_ & ~new_n20920_ & ~new_n20897_ & ~new_n20919_;
  assign new_n20897_ = ~new_n20913_ & ~new_n20914_ & new_n20908_ & (~new_n20905_ | ~new_n20898_);
  assign new_n20898_ = new_n20904_ & new_n20899_ & new_n20902_;
  assign new_n20899_ = \all_features[783]  & ~new_n20900_ & \all_features[782] ;
  assign new_n20900_ = ~\all_features[781]  & ~\all_features[780]  & ~\all_features[779]  & ~new_n20901_ & ~\all_features[778] ;
  assign new_n20901_ = \all_features[776]  & \all_features[777] ;
  assign new_n20902_ = \all_features[783]  & (\all_features[782]  | (new_n20903_ & (\all_features[778]  | \all_features[779]  | \all_features[777] )));
  assign new_n20903_ = \all_features[780]  & \all_features[781] ;
  assign new_n20904_ = \all_features[783]  & (\all_features[781]  | \all_features[782]  | \all_features[780] );
  assign new_n20905_ = \all_features[783]  & (\all_features[782]  | new_n20906_);
  assign new_n20906_ = \all_features[781]  & (\all_features[778]  | \all_features[779]  | \all_features[780]  | ~new_n20907_);
  assign new_n20907_ = ~\all_features[776]  & ~\all_features[777] ;
  assign new_n20908_ = ~new_n20909_ & ~new_n20911_;
  assign new_n20909_ = ~new_n20910_ & ~\all_features[783] ;
  assign new_n20910_ = \all_features[781]  & \all_features[782]  & (\all_features[780]  | (\all_features[778]  & \all_features[779]  & \all_features[777] ));
  assign new_n20911_ = ~\all_features[783]  & (~\all_features[782]  | (~\all_features[780]  & ~\all_features[781]  & ~new_n20912_));
  assign new_n20912_ = \all_features[778]  & \all_features[779] ;
  assign new_n20913_ = ~\all_features[783]  & (~\all_features[782]  | (~\all_features[781]  & (new_n20907_ | ~new_n20912_ | ~\all_features[780] )));
  assign new_n20914_ = ~\all_features[783]  & (~\all_features[782]  | ~new_n20903_ | ~new_n20901_ | ~new_n20912_);
  assign new_n20915_ = ~new_n20916_ & ~new_n20918_;
  assign new_n20916_ = ~\all_features[781]  & new_n20917_ & ((~\all_features[778]  & new_n20907_) | ~\all_features[780]  | ~\all_features[779] );
  assign new_n20917_ = ~\all_features[782]  & ~\all_features[783] ;
  assign new_n20918_ = ~\all_features[783]  & ~\all_features[782]  & ~\all_features[781]  & ~\all_features[779]  & ~\all_features[780] ;
  assign new_n20919_ = new_n20917_ & (~\all_features[781]  | (~\all_features[780]  & (~\all_features[779]  | (~\all_features[778]  & ~\all_features[777] ))));
  assign new_n20920_ = new_n20917_ & (~\all_features[779]  | ~new_n20903_ | (~\all_features[778]  & ~new_n20901_));
  assign new_n20921_ = new_n20915_ & new_n20908_ & new_n20922_ & ~new_n20913_ & ~new_n20914_;
  assign new_n20922_ = ~new_n20919_ & ~new_n20920_;
  assign new_n20923_ = new_n20956_ & new_n20924_ & new_n20954_;
  assign new_n20924_ = new_n20925_ & new_n20945_;
  assign new_n20925_ = ~new_n20944_ & (new_n20939_ | (~new_n20941_ & (new_n20942_ | (~new_n20926_ & ~new_n20943_))));
  assign new_n20926_ = ~new_n20933_ & (new_n20935_ | (~new_n20937_ & (~new_n20938_ | new_n20927_)));
  assign new_n20927_ = \all_features[2823]  & ((~new_n20932_ & ~\all_features[2821]  & \all_features[2822] ) | (~new_n20930_ & (\all_features[2822]  | (~new_n20928_ & \all_features[2821] ))));
  assign new_n20928_ = new_n20929_ & ~\all_features[2820]  & ~\all_features[2818]  & ~\all_features[2819] ;
  assign new_n20929_ = ~\all_features[2816]  & ~\all_features[2817] ;
  assign new_n20930_ = \all_features[2823]  & (\all_features[2822]  | (new_n20931_ & (\all_features[2818]  | \all_features[2819]  | \all_features[2817] )));
  assign new_n20931_ = \all_features[2820]  & \all_features[2821] ;
  assign new_n20932_ = (~\all_features[2818]  & ~\all_features[2819]  & ~\all_features[2820]  & (~\all_features[2817]  | ~\all_features[2816] )) | (\all_features[2820]  & (\all_features[2818]  | \all_features[2819] ));
  assign new_n20933_ = ~\all_features[2823]  & (~\all_features[2822]  | (~\all_features[2821]  & (new_n20929_ | ~new_n20934_ | ~\all_features[2820] )));
  assign new_n20934_ = \all_features[2818]  & \all_features[2819] ;
  assign new_n20935_ = ~new_n20936_ & ~\all_features[2823] ;
  assign new_n20936_ = \all_features[2821]  & \all_features[2822]  & (\all_features[2820]  | (\all_features[2818]  & \all_features[2819]  & \all_features[2817] ));
  assign new_n20937_ = ~\all_features[2823]  & (~new_n20934_ | ~\all_features[2816]  | ~\all_features[2817]  | ~\all_features[2822]  | ~new_n20931_);
  assign new_n20938_ = \all_features[2823]  & (\all_features[2821]  | \all_features[2822]  | \all_features[2820] );
  assign new_n20939_ = ~\all_features[2821]  & new_n20940_ & ((~\all_features[2818]  & new_n20929_) | ~\all_features[2820]  | ~\all_features[2819] );
  assign new_n20940_ = ~\all_features[2822]  & ~\all_features[2823] ;
  assign new_n20941_ = new_n20940_ & (~\all_features[2821]  | (~\all_features[2820]  & (~\all_features[2819]  | (~\all_features[2818]  & ~\all_features[2817] ))));
  assign new_n20942_ = new_n20940_ & (~new_n20931_ | ~\all_features[2819]  | (~\all_features[2818]  & (~\all_features[2816]  | ~\all_features[2817] )));
  assign new_n20943_ = ~\all_features[2823]  & (~\all_features[2822]  | (~\all_features[2820]  & ~\all_features[2821]  & ~new_n20934_));
  assign new_n20944_ = ~\all_features[2823]  & ~\all_features[2822]  & ~\all_features[2821]  & ~\all_features[2819]  & ~\all_features[2820] ;
  assign new_n20945_ = new_n20951_ & (~new_n20952_ | (new_n20953_ & (new_n20946_ | new_n20935_ | new_n20937_)));
  assign new_n20946_ = new_n20947_ & (~new_n20948_ | (~new_n20950_ & \all_features[2821]  & \all_features[2822]  & \all_features[2823] ));
  assign new_n20947_ = \all_features[2823]  & (\all_features[2822]  | (~new_n20928_ & \all_features[2821] ));
  assign new_n20948_ = \all_features[2823]  & \all_features[2822]  & ~new_n20949_ & new_n20930_;
  assign new_n20949_ = ~\all_features[2818]  & ~\all_features[2819]  & ~\all_features[2820]  & ~\all_features[2821]  & (~\all_features[2817]  | ~\all_features[2816] );
  assign new_n20950_ = ~\all_features[2819]  & ~\all_features[2820]  & (~\all_features[2818]  | new_n20929_);
  assign new_n20951_ = ~new_n20939_ & ~new_n20944_;
  assign new_n20952_ = ~new_n20941_ & ~new_n20942_;
  assign new_n20953_ = ~new_n20943_ & ~new_n20933_;
  assign new_n20954_ = new_n20952_ & ~new_n20955_ & new_n20951_;
  assign new_n20955_ = ~new_n20943_ & ~new_n20933_ & ~new_n20935_ & ~new_n20937_ & (~new_n20948_ | ~new_n20947_);
  assign new_n20956_ = new_n20952_ & new_n20951_ & new_n20953_ & ~new_n20935_ & ~new_n20937_;
  assign new_n20957_ = new_n10906_ & new_n10908_;
  assign new_n20958_ = ~new_n17849_ & new_n20959_;
  assign new_n20959_ = new_n15676_ & new_n15702_;
  assign new_n20960_ = ~new_n19125_ & (~new_n19127_ | ~new_n19096_);
  assign new_n20961_ = ~new_n21051_ & (~new_n20962_ | (~new_n21050_ & new_n21013_ & (~new_n20968_ | ~new_n20964_)));
  assign new_n20962_ = new_n20963_ & (~new_n20975_ | (~new_n20976_ & new_n21012_) | (new_n21011_ & ~new_n21012_));
  assign new_n20963_ = (new_n20968_ | ~new_n20964_) & (new_n12686_ | ~new_n20972_) & (~new_n20970_ | ~new_n20973_);
  assign new_n20964_ = new_n20965_ & ~new_n8927_ & new_n20967_;
  assign new_n20965_ = new_n10871_ & (new_n10868_ | new_n20966_);
  assign new_n20966_ = new_n10840_ & new_n10861_;
  assign new_n20967_ = new_n12933_ & new_n12910_ & new_n12936_;
  assign new_n20968_ = new_n14947_ & ~new_n20969_ & new_n14924_;
  assign new_n20969_ = ~new_n20731_ & ~new_n14950_;
  assign new_n20970_ = new_n20971_ & ~new_n20967_ & ~new_n13437_;
  assign new_n20971_ = new_n16454_ & new_n20242_;
  assign new_n20972_ = new_n8927_ & ~new_n12758_ & new_n20967_;
  assign new_n20973_ = ~new_n20974_ & new_n10738_;
  assign new_n20974_ = new_n10763_ & new_n10767_;
  assign new_n20975_ = ~new_n20967_ & new_n13437_;
  assign new_n20976_ = new_n20977_ & ~new_n21003_ & ~new_n21007_;
  assign new_n20977_ = ~new_n20978_ & ~new_n21001_;
  assign new_n20978_ = new_n20996_ & ~new_n21000_ & ~new_n20979_ & ~new_n20999_;
  assign new_n20979_ = ~new_n20992_ & ~new_n20994_ & new_n20987_ & (~new_n20995_ | ~new_n20980_);
  assign new_n20980_ = new_n20986_ & new_n20981_ & new_n20983_;
  assign new_n20981_ = \all_features[4303]  & (\all_features[4302]  | (new_n20982_ & (\all_features[4298]  | \all_features[4299]  | \all_features[4297] )));
  assign new_n20982_ = \all_features[4300]  & \all_features[4301] ;
  assign new_n20983_ = \all_features[4302]  & \all_features[4303]  & (\all_features[4300]  | \all_features[4301]  | new_n20984_ | ~new_n20985_);
  assign new_n20984_ = \all_features[4296]  & \all_features[4297] ;
  assign new_n20985_ = ~\all_features[4298]  & ~\all_features[4299] ;
  assign new_n20986_ = \all_features[4303]  & (\all_features[4301]  | \all_features[4302]  | \all_features[4300] );
  assign new_n20987_ = ~new_n20988_ & ~new_n20990_;
  assign new_n20988_ = ~\all_features[4303]  & (~\all_features[4302]  | (~\all_features[4300]  & ~\all_features[4301]  & ~new_n20989_));
  assign new_n20989_ = \all_features[4298]  & \all_features[4299] ;
  assign new_n20990_ = ~new_n20991_ & ~\all_features[4303] ;
  assign new_n20991_ = \all_features[4301]  & \all_features[4302]  & (\all_features[4300]  | (\all_features[4298]  & \all_features[4299]  & \all_features[4297] ));
  assign new_n20992_ = ~\all_features[4303]  & (~\all_features[4302]  | (~\all_features[4301]  & (new_n20993_ | ~new_n20989_ | ~\all_features[4300] )));
  assign new_n20993_ = ~\all_features[4296]  & ~\all_features[4297] ;
  assign new_n20994_ = ~\all_features[4303]  & (~\all_features[4302]  | ~new_n20984_ | ~new_n20982_ | ~new_n20989_);
  assign new_n20995_ = \all_features[4303]  & (\all_features[4302]  | (\all_features[4301]  & (\all_features[4300]  | ~new_n20985_ | ~new_n20993_)));
  assign new_n20996_ = ~new_n20997_ & (\all_features[4299]  | \all_features[4300]  | \all_features[4301]  | \all_features[4302]  | \all_features[4303] );
  assign new_n20997_ = ~\all_features[4301]  & new_n20998_ & ((~\all_features[4298]  & new_n20993_) | ~\all_features[4300]  | ~\all_features[4299] );
  assign new_n20998_ = ~\all_features[4302]  & ~\all_features[4303] ;
  assign new_n20999_ = new_n20998_ & (~\all_features[4301]  | (~\all_features[4300]  & (~\all_features[4299]  | (~\all_features[4298]  & ~\all_features[4297] ))));
  assign new_n21000_ = new_n20998_ & (~\all_features[4299]  | ~new_n20982_ | (~\all_features[4298]  & ~new_n20984_));
  assign new_n21001_ = new_n20996_ & new_n20987_ & new_n21002_ & ~new_n20992_ & ~new_n20994_;
  assign new_n21002_ = ~new_n20999_ & ~new_n21000_;
  assign new_n21003_ = ~new_n21004_ & (\all_features[4299]  | \all_features[4300]  | \all_features[4301]  | \all_features[4302]  | \all_features[4303] );
  assign new_n21004_ = ~new_n20997_ & (new_n20999_ | (~new_n21000_ & (new_n20988_ | (~new_n21005_ & ~new_n20992_))));
  assign new_n21005_ = ~new_n20990_ & (new_n20994_ | (new_n20986_ & (~new_n20995_ | (~new_n21006_ & new_n20981_))));
  assign new_n21006_ = ~\all_features[4301]  & \all_features[4302]  & \all_features[4303]  & (\all_features[4300]  ? new_n20985_ : (new_n20984_ | ~new_n20985_));
  assign new_n21007_ = new_n20996_ & (~new_n21002_ | (~new_n21008_ & ~new_n20988_ & ~new_n20992_));
  assign new_n21008_ = ~new_n20990_ & ~new_n20994_ & (~new_n20986_ | ~new_n20995_ | new_n21009_);
  assign new_n21009_ = new_n20981_ & new_n20983_ & (new_n21010_ | ~\all_features[4301]  | ~\all_features[4302]  | ~\all_features[4303] );
  assign new_n21010_ = ~\all_features[4299]  & ~\all_features[4300]  & (~\all_features[4298]  | new_n20993_);
  assign new_n21011_ = ~new_n18985_ & (~new_n18962_ | ~new_n20442_);
  assign new_n21012_ = new_n9122_ & new_n16648_;
  assign new_n21013_ = new_n21014_ & (~new_n12686_ | ~new_n20972_) & (~new_n20970_ | new_n20973_);
  assign new_n21014_ = ~new_n20967_ | ((new_n20965_ | new_n8927_) & (~new_n12758_ | ~new_n21015_ | ~new_n8927_));
  assign new_n21015_ = new_n21016_ & ~new_n21045_ & ~new_n21048_;
  assign new_n21016_ = ~new_n21017_ & ~new_n21041_;
  assign new_n21017_ = new_n21032_ & (~new_n21037_ | (~new_n21035_ & ~new_n21018_ & ~new_n21040_));
  assign new_n21018_ = ~new_n21030_ & ~new_n21028_ & (~new_n21031_ | ~new_n21027_ | new_n21019_);
  assign new_n21019_ = new_n21020_ & new_n21022_ & (new_n21025_ | ~\all_features[1629]  | ~\all_features[1630]  | ~\all_features[1631] );
  assign new_n21020_ = \all_features[1631]  & (\all_features[1630]  | (new_n21021_ & (\all_features[1626]  | \all_features[1627]  | \all_features[1625] )));
  assign new_n21021_ = \all_features[1628]  & \all_features[1629] ;
  assign new_n21022_ = \all_features[1630]  & \all_features[1631]  & (\all_features[1628]  | \all_features[1629]  | new_n21024_ | ~new_n21023_);
  assign new_n21023_ = ~\all_features[1626]  & ~\all_features[1627] ;
  assign new_n21024_ = \all_features[1624]  & \all_features[1625] ;
  assign new_n21025_ = ~\all_features[1627]  & ~\all_features[1628]  & (~\all_features[1626]  | new_n21026_);
  assign new_n21026_ = ~\all_features[1624]  & ~\all_features[1625] ;
  assign new_n21027_ = \all_features[1631]  & (\all_features[1630]  | (\all_features[1629]  & (\all_features[1628]  | ~new_n21023_ | ~new_n21026_)));
  assign new_n21028_ = ~new_n21029_ & ~\all_features[1631] ;
  assign new_n21029_ = \all_features[1629]  & \all_features[1630]  & (\all_features[1628]  | (\all_features[1626]  & \all_features[1627]  & \all_features[1625] ));
  assign new_n21030_ = ~\all_features[1631]  & (~new_n21024_ | ~\all_features[1626]  | ~\all_features[1627]  | ~\all_features[1630]  | ~new_n21021_);
  assign new_n21031_ = \all_features[1631]  & (\all_features[1629]  | \all_features[1630]  | \all_features[1628] );
  assign new_n21032_ = ~new_n21033_ & (\all_features[1627]  | \all_features[1628]  | \all_features[1629]  | \all_features[1630]  | \all_features[1631] );
  assign new_n21033_ = ~\all_features[1629]  & new_n21034_ & ((~\all_features[1626]  & new_n21026_) | ~\all_features[1628]  | ~\all_features[1627] );
  assign new_n21034_ = ~\all_features[1630]  & ~\all_features[1631] ;
  assign new_n21035_ = ~\all_features[1631]  & (~\all_features[1630]  | new_n21036_);
  assign new_n21036_ = ~\all_features[1629]  & (new_n21026_ | ~\all_features[1627]  | ~\all_features[1628]  | ~\all_features[1626] );
  assign new_n21037_ = ~new_n21038_ & ~new_n21039_;
  assign new_n21038_ = new_n21034_ & (~\all_features[1627]  | ~new_n21021_ | (~new_n21024_ & ~\all_features[1626] ));
  assign new_n21039_ = new_n21034_ & (~\all_features[1629]  | (~\all_features[1628]  & (~\all_features[1627]  | (~\all_features[1626]  & ~\all_features[1625] ))));
  assign new_n21040_ = ~\all_features[1631]  & (~\all_features[1630]  | (~\all_features[1629]  & ~\all_features[1628]  & (~\all_features[1627]  | ~\all_features[1626] )));
  assign new_n21041_ = ~new_n21042_ & (\all_features[1627]  | \all_features[1628]  | \all_features[1629]  | \all_features[1630]  | \all_features[1631] );
  assign new_n21042_ = ~new_n21033_ & (new_n21039_ | (~new_n21038_ & (new_n21040_ | (~new_n21035_ & ~new_n21043_))));
  assign new_n21043_ = ~new_n21028_ & (new_n21030_ | (new_n21031_ & (~new_n21027_ | (~new_n21044_ & new_n21020_))));
  assign new_n21044_ = ~\all_features[1629]  & \all_features[1630]  & \all_features[1631]  & (\all_features[1628]  ? new_n21023_ : (new_n21024_ | ~new_n21023_));
  assign new_n21045_ = new_n21037_ & ~new_n21046_ & new_n21032_;
  assign new_n21046_ = ~new_n21040_ & ~new_n21030_ & ~new_n21028_ & ~new_n21035_ & ~new_n21047_;
  assign new_n21047_ = new_n21031_ & new_n21027_ & new_n21020_ & new_n21022_;
  assign new_n21048_ = new_n21032_ & new_n21049_ & ~new_n21028_ & ~new_n21039_;
  assign new_n21049_ = ~new_n21040_ & ~new_n21038_ & ~new_n21035_ & ~new_n21030_;
  assign new_n21050_ = ~new_n20967_ & ((~new_n21012_ & new_n21011_ & new_n13437_) | (~new_n20971_ & ~new_n13437_));
  assign new_n21051_ = new_n21012_ & ~new_n20976_ & new_n20975_;
  assign new_n21052_ = ~new_n21053_ & new_n21182_;
  assign new_n21053_ = new_n21054_ & (~new_n21056_ | (~new_n21133_ & ~new_n21134_));
  assign new_n21054_ = new_n21057_ & (~new_n21055_ | (~new_n19835_ & new_n21111_) | (~new_n21076_ & ~new_n21111_));
  assign new_n21055_ = ~new_n21056_ & new_n15751_;
  assign new_n21056_ = new_n9452_ & new_n9455_;
  assign new_n21057_ = new_n21056_ | new_n15751_ | (new_n21058_ ? ~new_n21059_ : new_n12187_);
  assign new_n21058_ = ~new_n7696_ & (~new_n7905_ | ~new_n7909_ | ~new_n7673_);
  assign new_n21059_ = ~new_n21071_ & new_n21072_;
  assign new_n21071_ = ~\all_features[5191]  & ~\all_features[5190]  & ~\all_features[5189]  & ~\all_features[5187]  & ~\all_features[5188] ;
  assign new_n21072_ = \all_features[5190]  | \all_features[5191]  | (~new_n21073_ & \all_features[5189]  & new_n21075_);
  assign new_n21073_ = ~\all_features[5188]  & (~\all_features[5187]  | (~\all_features[5186]  & ~\all_features[5185] ));
  assign new_n21075_ = \all_features[5187]  & \all_features[5188]  & \all_features[5189]  & (\all_features[5186]  | (\all_features[5185]  & \all_features[5184] ));
  assign new_n21076_ = ~new_n21106_ & (~new_n21108_ | new_n21077_);
  assign new_n21077_ = ~new_n21078_ & ~new_n21102_;
  assign new_n21078_ = new_n21094_ & (~new_n21097_ | (~new_n21079_ & ~new_n21100_ & ~new_n21101_));
  assign new_n21079_ = ~new_n21088_ & ~new_n21090_ & (~new_n21093_ | ~new_n21092_ | new_n21080_);
  assign new_n21080_ = new_n21081_ & new_n21083_ & (new_n21086_ | ~\all_features[1061]  | ~\all_features[1062]  | ~\all_features[1063] );
  assign new_n21081_ = \all_features[1063]  & (\all_features[1062]  | (new_n21082_ & (\all_features[1058]  | \all_features[1059]  | \all_features[1057] )));
  assign new_n21082_ = \all_features[1060]  & \all_features[1061] ;
  assign new_n21083_ = \all_features[1062]  & \all_features[1063]  & (\all_features[1060]  | \all_features[1061]  | new_n21084_ | ~new_n21085_);
  assign new_n21084_ = \all_features[1056]  & \all_features[1057] ;
  assign new_n21085_ = ~\all_features[1058]  & ~\all_features[1059] ;
  assign new_n21086_ = ~\all_features[1059]  & ~\all_features[1060]  & (~\all_features[1058]  | new_n21087_);
  assign new_n21087_ = ~\all_features[1056]  & ~\all_features[1057] ;
  assign new_n21088_ = ~new_n21089_ & ~\all_features[1063] ;
  assign new_n21089_ = \all_features[1061]  & \all_features[1062]  & (\all_features[1060]  | (\all_features[1058]  & \all_features[1059]  & \all_features[1057] ));
  assign new_n21090_ = ~\all_features[1063]  & (~\all_features[1062]  | ~new_n21091_ | ~new_n21084_ | ~new_n21082_);
  assign new_n21091_ = \all_features[1058]  & \all_features[1059] ;
  assign new_n21092_ = \all_features[1063]  & (\all_features[1062]  | (\all_features[1061]  & (\all_features[1060]  | ~new_n21085_ | ~new_n21087_)));
  assign new_n21093_ = \all_features[1063]  & (\all_features[1061]  | \all_features[1062]  | \all_features[1060] );
  assign new_n21094_ = ~new_n21095_ & (\all_features[1059]  | \all_features[1060]  | \all_features[1061]  | \all_features[1062]  | \all_features[1063] );
  assign new_n21095_ = ~\all_features[1061]  & new_n21096_ & ((~\all_features[1058]  & new_n21087_) | ~\all_features[1060]  | ~\all_features[1059] );
  assign new_n21096_ = ~\all_features[1062]  & ~\all_features[1063] ;
  assign new_n21097_ = ~new_n21098_ & ~new_n21099_;
  assign new_n21098_ = new_n21096_ & (~\all_features[1061]  | (~\all_features[1060]  & (~\all_features[1059]  | (~\all_features[1058]  & ~\all_features[1057] ))));
  assign new_n21099_ = new_n21096_ & (~\all_features[1059]  | ~new_n21082_ | (~\all_features[1058]  & ~new_n21084_));
  assign new_n21100_ = ~\all_features[1063]  & (~\all_features[1062]  | (~\all_features[1061]  & (new_n21087_ | ~new_n21091_ | ~\all_features[1060] )));
  assign new_n21101_ = ~\all_features[1063]  & (~\all_features[1062]  | (~\all_features[1060]  & ~\all_features[1061]  & ~new_n21091_));
  assign new_n21102_ = ~new_n21103_ & (\all_features[1059]  | \all_features[1060]  | \all_features[1061]  | \all_features[1062]  | \all_features[1063] );
  assign new_n21103_ = ~new_n21095_ & (new_n21098_ | (~new_n21099_ & (new_n21101_ | (~new_n21100_ & ~new_n21104_))));
  assign new_n21104_ = ~new_n21088_ & (new_n21090_ | (new_n21093_ & (~new_n21092_ | (~new_n21105_ & new_n21081_))));
  assign new_n21105_ = ~\all_features[1061]  & \all_features[1062]  & \all_features[1063]  & (\all_features[1060]  ? new_n21085_ : (new_n21084_ | ~new_n21085_));
  assign new_n21106_ = new_n21107_ & new_n21094_ & ~new_n21099_ & ~new_n21100_ & ~new_n21088_ & ~new_n21098_;
  assign new_n21107_ = ~new_n21090_ & ~new_n21101_;
  assign new_n21108_ = new_n21094_ & new_n21097_ & (new_n21109_ | new_n21088_ | new_n21100_ | ~new_n21107_);
  assign new_n21109_ = new_n21093_ & new_n21083_ & new_n21092_ & new_n21081_;
  assign new_n21111_ = new_n21112_ & ~new_n21116_ & ~new_n21117_;
  assign new_n21112_ = ~new_n21113_ & (\all_features[5667]  | \all_features[5668]  | \all_features[5669]  | \all_features[5670]  | \all_features[5671] );
  assign new_n21113_ = ~\all_features[5669]  & new_n21115_ & ((~\all_features[5666]  & new_n21114_) | ~\all_features[5668]  | ~\all_features[5667] );
  assign new_n21114_ = ~\all_features[5664]  & ~\all_features[5665] ;
  assign new_n21115_ = ~\all_features[5670]  & ~\all_features[5671] ;
  assign new_n21116_ = new_n21115_ & (~\all_features[5669]  | (~\all_features[5668]  & (~\all_features[5667]  | (~\all_features[5666]  & ~\all_features[5665] ))));
  assign new_n21117_ = new_n21115_ & (~\all_features[5667]  | ~new_n21118_ | (~\all_features[5666]  & ~new_n21119_));
  assign new_n21118_ = \all_features[5668]  & \all_features[5669] ;
  assign new_n21119_ = \all_features[5664]  & \all_features[5665] ;
  assign new_n21120_ = new_n21124_ & new_n21121_ & new_n21122_;
  assign new_n21121_ = \all_features[5671]  & (\all_features[5670]  | (new_n21118_ & (\all_features[5666]  | \all_features[5667]  | \all_features[5665] )));
  assign new_n21122_ = \all_features[5670]  & \all_features[5671]  & (\all_features[5668]  | \all_features[5669]  | new_n21119_ | ~new_n21123_);
  assign new_n21123_ = ~\all_features[5666]  & ~\all_features[5667] ;
  assign new_n21124_ = \all_features[5671]  & (\all_features[5669]  | \all_features[5670]  | \all_features[5668] );
  assign new_n21125_ = ~new_n21131_ & ~new_n21130_ & ~new_n21126_ & ~new_n21128_;
  assign new_n21126_ = ~\all_features[5671]  & (~\all_features[5670]  | (~\all_features[5669]  & (new_n21114_ | ~new_n21127_ | ~\all_features[5668] )));
  assign new_n21127_ = \all_features[5666]  & \all_features[5667] ;
  assign new_n21128_ = ~new_n21129_ & ~\all_features[5671] ;
  assign new_n21129_ = \all_features[5669]  & \all_features[5670]  & (\all_features[5668]  | (\all_features[5666]  & \all_features[5667]  & \all_features[5665] ));
  assign new_n21130_ = ~\all_features[5671]  & (~\all_features[5670]  | ~new_n21118_ | ~new_n21119_ | ~new_n21127_);
  assign new_n21131_ = ~\all_features[5671]  & (~\all_features[5670]  | (~\all_features[5668]  & ~\all_features[5669]  & ~new_n21127_));
  assign new_n21132_ = \all_features[5671]  & (\all_features[5670]  | (\all_features[5669]  & (\all_features[5668]  | ~new_n21114_ | ~new_n21123_)));
  assign new_n21133_ = new_n12655_ & new_n17251_;
  assign new_n21134_ = (new_n18597_ | ~new_n21163_ | (~new_n21135_ & ~new_n21164_)) & (new_n21166_ | new_n21135_ | new_n21164_);
  assign new_n21135_ = new_n21152_ & (new_n21161_ | (~new_n21160_ & ~new_n21136_));
  assign new_n21136_ = ~new_n21149_ & (new_n21151_ | (~new_n21148_ & (new_n21144_ | (~new_n21146_ & ~new_n21137_))));
  assign new_n21137_ = ~new_n21138_ & \all_features[4751]  & (\all_features[4750]  | \all_features[4749]  | \all_features[4748] );
  assign new_n21138_ = \all_features[4751]  & ((~new_n21143_ & ~\all_features[4749]  & \all_features[4750] ) | (~new_n21141_ & (\all_features[4750]  | (~new_n21139_ & \all_features[4749] ))));
  assign new_n21139_ = new_n21140_ & ~\all_features[4748]  & ~\all_features[4746]  & ~\all_features[4747] ;
  assign new_n21140_ = ~\all_features[4744]  & ~\all_features[4745] ;
  assign new_n21141_ = \all_features[4751]  & (\all_features[4750]  | (new_n21142_ & (\all_features[4746]  | \all_features[4747]  | \all_features[4745] )));
  assign new_n21142_ = \all_features[4748]  & \all_features[4749] ;
  assign new_n21143_ = (~\all_features[4746]  & ~\all_features[4747]  & ~\all_features[4748]  & (~\all_features[4745]  | ~\all_features[4744] )) | (\all_features[4748]  & (\all_features[4746]  | \all_features[4747] ));
  assign new_n21144_ = ~new_n21145_ & ~\all_features[4751] ;
  assign new_n21145_ = \all_features[4749]  & \all_features[4750]  & (\all_features[4748]  | (\all_features[4746]  & \all_features[4747]  & \all_features[4745] ));
  assign new_n21146_ = ~\all_features[4751]  & (~new_n21142_ | ~\all_features[4744]  | ~\all_features[4745]  | ~\all_features[4750]  | ~new_n21147_);
  assign new_n21147_ = \all_features[4746]  & \all_features[4747] ;
  assign new_n21148_ = ~\all_features[4751]  & (~\all_features[4750]  | (~\all_features[4749]  & (new_n21140_ | ~\all_features[4748]  | ~new_n21147_)));
  assign new_n21149_ = new_n21150_ & (~new_n21142_ | ~\all_features[4747]  | (~\all_features[4746]  & (~\all_features[4744]  | ~\all_features[4745] )));
  assign new_n21150_ = ~\all_features[4750]  & ~\all_features[4751] ;
  assign new_n21151_ = ~\all_features[4751]  & (~\all_features[4750]  | (~\all_features[4748]  & ~\all_features[4749]  & ~new_n21147_));
  assign new_n21152_ = ~new_n21158_ & new_n21159_ & (new_n21146_ | new_n21144_ | new_n21153_);
  assign new_n21153_ = new_n21154_ & (~new_n21155_ | (~new_n21157_ & \all_features[4749]  & \all_features[4750]  & \all_features[4751] ));
  assign new_n21154_ = \all_features[4751]  & (\all_features[4750]  | (~new_n21139_ & \all_features[4749] ));
  assign new_n21155_ = \all_features[4751]  & \all_features[4750]  & ~new_n21156_ & new_n21141_;
  assign new_n21156_ = ~\all_features[4746]  & ~\all_features[4747]  & ~\all_features[4748]  & ~\all_features[4749]  & (~\all_features[4745]  | ~\all_features[4744] );
  assign new_n21157_ = ~\all_features[4747]  & ~\all_features[4748]  & (~\all_features[4746]  | new_n21140_);
  assign new_n21158_ = ~new_n21144_ & ~new_n21146_ & ~new_n21148_ & ~new_n21151_ & (~new_n21155_ | ~new_n21154_);
  assign new_n21159_ = ~new_n21162_ & ~new_n21151_ & ~new_n21161_ & ~new_n21149_ & ~new_n21160_ & ~new_n21148_;
  assign new_n21160_ = new_n21150_ & (~\all_features[4749]  | (~\all_features[4748]  & (~\all_features[4747]  | (~\all_features[4746]  & ~\all_features[4745] ))));
  assign new_n21161_ = ~\all_features[4749]  & new_n21150_ & ((~\all_features[4746]  & new_n21140_) | ~\all_features[4748]  | ~\all_features[4747] );
  assign new_n21162_ = ~\all_features[4751]  & ~\all_features[4750]  & ~\all_features[4749]  & ~\all_features[4747]  & ~\all_features[4748] ;
  assign new_n21163_ = new_n18627_ & new_n18631_;
  assign new_n21164_ = new_n21165_ & ~new_n21162_ & ~new_n21146_ & ~new_n21144_ & ~new_n21160_;
  assign new_n21165_ = ~new_n21151_ & ~new_n21161_ & ~new_n21148_ & ~new_n21149_;
  assign new_n21166_ = new_n21172_ & new_n21167_ & ~new_n21181_ & ~new_n21180_ & ~new_n21176_ & ~new_n21178_;
  assign new_n21167_ = ~new_n21168_ & (\all_features[5747]  | \all_features[5748]  | \all_features[5749]  | \all_features[5750]  | \all_features[5751] );
  assign new_n21168_ = ~\all_features[5751]  & (~\all_features[5750]  | ~new_n21169_ | ~new_n21170_ | ~new_n21171_);
  assign new_n21169_ = \all_features[5744]  & \all_features[5745] ;
  assign new_n21170_ = \all_features[5746]  & \all_features[5747] ;
  assign new_n21171_ = \all_features[5748]  & \all_features[5749] ;
  assign new_n21172_ = ~new_n21173_ & ~new_n21175_;
  assign new_n21173_ = new_n21174_ & (~\all_features[5749]  | (~\all_features[5748]  & (~\all_features[5747]  | (~\all_features[5746]  & ~\all_features[5745] ))));
  assign new_n21174_ = ~\all_features[5750]  & ~\all_features[5751] ;
  assign new_n21175_ = new_n21174_ & (~\all_features[5747]  | ~new_n21171_ | (~\all_features[5746]  & ~new_n21169_));
  assign new_n21176_ = ~new_n21177_ & ~\all_features[5751] ;
  assign new_n21177_ = \all_features[5749]  & \all_features[5750]  & (\all_features[5748]  | (\all_features[5746]  & \all_features[5747]  & \all_features[5745] ));
  assign new_n21178_ = ~\all_features[5749]  & new_n21174_ & ((~\all_features[5746]  & new_n21179_) | ~\all_features[5748]  | ~\all_features[5747] );
  assign new_n21179_ = ~\all_features[5744]  & ~\all_features[5745] ;
  assign new_n21180_ = ~\all_features[5751]  & (~\all_features[5750]  | (~\all_features[5748]  & ~\all_features[5749]  & ~new_n21170_));
  assign new_n21181_ = ~\all_features[5751]  & (~\all_features[5750]  | (~\all_features[5749]  & (new_n21179_ | ~\all_features[5748]  | ~new_n21170_)));
  assign new_n21182_ = new_n21183_ & (~new_n21055_ | (new_n19835_ & new_n21111_) | (new_n21076_ & ~new_n21111_));
  assign new_n21183_ = (new_n21134_ | new_n21133_ | ~new_n21056_) & (new_n15751_ | new_n21059_ | ~new_n21058_ | new_n21056_);
  assign new_n21184_ = new_n20237_ ? (~new_n21185_ ^ new_n21247_) : (new_n21185_ ^ new_n21247_);
  assign new_n21185_ = ~new_n21186_ & new_n21246_;
  assign new_n21186_ = ~new_n21187_ & (new_n21188_ | (new_n21206_ & new_n21209_) | (new_n21210_ & ~new_n21209_));
  assign new_n21187_ = new_n9098_ & new_n21198_ & ~new_n21200_ & new_n21188_;
  assign new_n21188_ = new_n17734_ & new_n21189_ & new_n21194_;
  assign new_n21189_ = new_n17711_ & new_n21190_;
  assign new_n21190_ = new_n17729_ & (~new_n17735_ | (~new_n21191_ & ~new_n17723_ & ~new_n17727_));
  assign new_n21191_ = ~new_n17728_ & ~new_n17721_ & (~new_n17719_ | ~new_n17725_ | new_n21192_);
  assign new_n21192_ = new_n17714_ & new_n17716_ & (new_n21193_ | ~\all_features[5437]  | ~\all_features[5438]  | ~\all_features[5439] );
  assign new_n21193_ = ~\all_features[5435]  & ~\all_features[5436]  & (~\all_features[5434]  | new_n17726_);
  assign new_n21194_ = ~new_n21195_ & (\all_features[5435]  | \all_features[5436]  | \all_features[5437]  | \all_features[5438]  | \all_features[5439] );
  assign new_n21195_ = ~new_n17730_ & (new_n17732_ | (~new_n17733_ & (new_n17723_ | (~new_n17727_ & ~new_n21196_))));
  assign new_n21196_ = ~new_n17721_ & (new_n17728_ | (new_n17719_ & (~new_n17725_ | (~new_n21197_ & new_n17714_))));
  assign new_n21197_ = ~\all_features[5437]  & \all_features[5438]  & \all_features[5439]  & (\all_features[5436]  ? new_n17717_ : (new_n17718_ | ~new_n17717_));
  assign new_n21198_ = ~new_n21199_ & new_n10911_;
  assign new_n21199_ = new_n10939_ & new_n10943_;
  assign new_n21200_ = new_n10099_ & (new_n10097_ | (new_n10072_ & new_n21201_));
  assign new_n21201_ = ~new_n10074_ & (new_n10077_ | (~new_n10089_ & (new_n10088_ | (~new_n21202_ & ~new_n10091_))));
  assign new_n21202_ = ~new_n10093_ & (new_n10095_ | (~new_n10094_ & (~new_n21205_ | new_n21203_)));
  assign new_n21203_ = \all_features[4543]  & ((~new_n21204_ & ~\all_features[4541]  & \all_features[4542] ) | (~new_n10083_ & (\all_features[4542]  | (~new_n10081_ & \all_features[4541] ))));
  assign new_n21204_ = (~\all_features[4538]  & ~\all_features[4539]  & ~\all_features[4540]  & (~\all_features[4537]  | ~\all_features[4536] )) | (\all_features[4540]  & (\all_features[4538]  | \all_features[4539] ));
  assign new_n21205_ = \all_features[4543]  & (\all_features[4541]  | \all_features[4542]  | \all_features[4540] );
  assign new_n21206_ = new_n19843_ ? ~new_n21208_ : new_n21207_;
  assign new_n21207_ = ~new_n14954_ & new_n14985_;
  assign new_n21208_ = ~new_n9995_ & (~new_n9993_ | ~new_n9968_);
  assign new_n21209_ = new_n10271_ & (new_n10249_ | ~new_n10272_);
  assign new_n21210_ = new_n16800_ & (~new_n21211_ | ~new_n21241_) & (new_n20778_ | new_n16778_);
  assign new_n21211_ = ~new_n21212_ & ~new_n21233_;
  assign new_n21212_ = ~new_n21213_ & (\all_features[1643]  | \all_features[1644]  | \all_features[1645]  | \all_features[1646]  | \all_features[1647] );
  assign new_n21213_ = ~new_n21227_ & (new_n21232_ | (~new_n21229_ & (new_n21230_ | (~new_n21231_ & ~new_n21214_))));
  assign new_n21214_ = ~new_n21215_ & (new_n21224_ | (new_n21226_ & (~new_n21217_ | (~new_n21222_ & new_n21220_))));
  assign new_n21215_ = ~new_n21216_ & ~\all_features[1647] ;
  assign new_n21216_ = \all_features[1645]  & \all_features[1646]  & (\all_features[1644]  | (\all_features[1642]  & \all_features[1643]  & \all_features[1641] ));
  assign new_n21217_ = \all_features[1647]  & (\all_features[1646]  | (\all_features[1645]  & (\all_features[1644]  | ~new_n21219_ | ~new_n21218_)));
  assign new_n21218_ = ~\all_features[1640]  & ~\all_features[1641] ;
  assign new_n21219_ = ~\all_features[1642]  & ~\all_features[1643] ;
  assign new_n21220_ = \all_features[1647]  & (\all_features[1646]  | (new_n21221_ & (\all_features[1642]  | \all_features[1643]  | \all_features[1641] )));
  assign new_n21221_ = \all_features[1644]  & \all_features[1645] ;
  assign new_n21222_ = ~\all_features[1645]  & \all_features[1646]  & \all_features[1647]  & (\all_features[1644]  ? new_n21219_ : (new_n21223_ | ~new_n21219_));
  assign new_n21223_ = \all_features[1640]  & \all_features[1641] ;
  assign new_n21224_ = ~\all_features[1647]  & (~\all_features[1646]  | ~new_n21223_ | ~new_n21221_ | ~new_n21225_);
  assign new_n21225_ = \all_features[1642]  & \all_features[1643] ;
  assign new_n21226_ = \all_features[1647]  & (\all_features[1645]  | \all_features[1646]  | \all_features[1644] );
  assign new_n21227_ = ~\all_features[1645]  & new_n21228_ & ((~\all_features[1642]  & new_n21218_) | ~\all_features[1644]  | ~\all_features[1643] );
  assign new_n21228_ = ~\all_features[1646]  & ~\all_features[1647] ;
  assign new_n21229_ = new_n21228_ & (~\all_features[1643]  | ~new_n21221_ | (~\all_features[1642]  & ~new_n21223_));
  assign new_n21230_ = ~\all_features[1647]  & (~\all_features[1646]  | (~\all_features[1644]  & ~\all_features[1645]  & ~new_n21225_));
  assign new_n21231_ = ~\all_features[1647]  & (~\all_features[1646]  | (~\all_features[1645]  & (new_n21218_ | ~new_n21225_ | ~\all_features[1644] )));
  assign new_n21232_ = new_n21228_ & (~\all_features[1645]  | (~\all_features[1644]  & (~\all_features[1643]  | (~\all_features[1642]  & ~\all_features[1641] ))));
  assign new_n21233_ = new_n21239_ & (~new_n21240_ | (~new_n21234_ & ~new_n21230_ & ~new_n21231_));
  assign new_n21234_ = new_n21237_ & ((~new_n21235_ & new_n21220_ & new_n21238_) | ~new_n21226_ | ~new_n21217_);
  assign new_n21235_ = \all_features[1647]  & \all_features[1646]  & ~new_n21236_ & \all_features[1645] ;
  assign new_n21236_ = ~\all_features[1643]  & ~\all_features[1644]  & (~\all_features[1642]  | new_n21218_);
  assign new_n21237_ = ~new_n21215_ & ~new_n21224_;
  assign new_n21238_ = \all_features[1646]  & \all_features[1647]  & (\all_features[1644]  | \all_features[1645]  | new_n21223_ | ~new_n21219_);
  assign new_n21239_ = ~new_n21227_ & (\all_features[1643]  | \all_features[1644]  | \all_features[1645]  | \all_features[1646]  | \all_features[1647] );
  assign new_n21240_ = ~new_n21229_ & ~new_n21232_;
  assign new_n21241_ = ~new_n21242_ & ~new_n21245_;
  assign new_n21242_ = new_n21240_ & ~new_n21243_ & new_n21239_;
  assign new_n21243_ = new_n21244_ & (~new_n21238_ | ~new_n21226_ | ~new_n21217_ | ~new_n21220_);
  assign new_n21244_ = ~new_n21224_ & ~new_n21215_ & ~new_n21230_ & ~new_n21231_;
  assign new_n21245_ = new_n21237_ & new_n21239_ & ~new_n21232_ & ~new_n21231_ & ~new_n21229_ & ~new_n21230_;
  assign new_n21246_ = (~new_n21200_ & new_n21198_ & new_n21188_) | (~new_n21188_ & (new_n21209_ ? ~new_n21206_ : ~new_n21210_));
  assign new_n21247_ = ~new_n21248_ & (~new_n21343_ | (~new_n21312_ & ~new_n21334_ & ~new_n21345_));
  assign new_n21248_ = (~new_n21249_ | new_n21280_) & (new_n20489_ | ~new_n13773_ | ~new_n11297_ | ~new_n21280_);
  assign new_n21249_ = ~new_n21250_ & (~new_n21278_ | (~new_n21252_ & ~new_n21274_));
  assign new_n21250_ = new_n13518_ & new_n21251_ & new_n13090_;
  assign new_n21251_ = new_n13067_ & new_n13095_;
  assign new_n21252_ = new_n21271_ & ~new_n21253_ & new_n21267_;
  assign new_n21253_ = ~new_n21261_ & ~new_n21263_ & ~new_n21265_ & ~new_n21266_ & (~new_n21257_ | ~new_n21254_);
  assign new_n21254_ = \all_features[1287]  & (\all_features[1286]  | (~new_n21255_ & \all_features[1285] ));
  assign new_n21255_ = new_n21256_ & ~\all_features[1284]  & ~\all_features[1282]  & ~\all_features[1283] ;
  assign new_n21256_ = ~\all_features[1280]  & ~\all_features[1281] ;
  assign new_n21257_ = \all_features[1287]  & \all_features[1286]  & ~new_n21260_ & new_n21258_;
  assign new_n21258_ = \all_features[1287]  & (\all_features[1286]  | (new_n21259_ & (\all_features[1282]  | \all_features[1283]  | \all_features[1281] )));
  assign new_n21259_ = \all_features[1284]  & \all_features[1285] ;
  assign new_n21260_ = ~\all_features[1282]  & ~\all_features[1283]  & ~\all_features[1284]  & ~\all_features[1285]  & (~\all_features[1281]  | ~\all_features[1280] );
  assign new_n21261_ = ~new_n21262_ & ~\all_features[1287] ;
  assign new_n21262_ = \all_features[1285]  & \all_features[1286]  & (\all_features[1284]  | (\all_features[1282]  & \all_features[1283]  & \all_features[1281] ));
  assign new_n21263_ = ~\all_features[1287]  & (~\all_features[1286]  | (~\all_features[1284]  & ~\all_features[1285]  & ~new_n21264_));
  assign new_n21264_ = \all_features[1282]  & \all_features[1283] ;
  assign new_n21265_ = ~\all_features[1287]  & (~new_n21259_ | ~\all_features[1280]  | ~\all_features[1281]  | ~\all_features[1286]  | ~new_n21264_);
  assign new_n21266_ = ~\all_features[1287]  & (~\all_features[1286]  | (~\all_features[1285]  & (new_n21256_ | ~\all_features[1284]  | ~new_n21264_)));
  assign new_n21267_ = ~new_n21268_ & ~new_n21270_;
  assign new_n21268_ = new_n21269_ & (~new_n21259_ | ~\all_features[1283]  | (~\all_features[1282]  & (~\all_features[1280]  | ~\all_features[1281] )));
  assign new_n21269_ = ~\all_features[1286]  & ~\all_features[1287] ;
  assign new_n21270_ = new_n21269_ & (~\all_features[1285]  | (~\all_features[1284]  & (~\all_features[1283]  | (~\all_features[1282]  & ~\all_features[1281] ))));
  assign new_n21271_ = ~new_n21272_ & ~new_n21273_;
  assign new_n21272_ = new_n21269_ & ~\all_features[1285]  & ~\all_features[1283]  & ~\all_features[1284] ;
  assign new_n21273_ = ~\all_features[1285]  & new_n21269_ & ((~\all_features[1282]  & new_n21256_) | ~\all_features[1284]  | ~\all_features[1283] );
  assign new_n21274_ = new_n21271_ & (~new_n21267_ | (~new_n21275_ & ~new_n21263_ & ~new_n21266_));
  assign new_n21275_ = ~new_n21261_ & ~new_n21265_ & (~new_n21254_ | (~new_n21276_ & new_n21257_));
  assign new_n21276_ = \all_features[1287]  & \all_features[1286]  & ~new_n21277_ & \all_features[1285] ;
  assign new_n21277_ = ~\all_features[1283]  & ~\all_features[1284]  & (~\all_features[1282]  | new_n21256_);
  assign new_n21278_ = new_n21267_ & new_n21279_ & ~new_n21266_ & ~new_n21273_ & ~new_n21261_ & ~new_n21265_;
  assign new_n21279_ = ~new_n21272_ & ~new_n21263_;
  assign new_n21280_ = ~new_n21281_ & (new_n21296_ | new_n21298_ | new_n21290_ | new_n21307_ | ~new_n21311_);
  assign new_n21281_ = new_n21303_ & (new_n21282_ | new_n21306_) & (new_n21296_ | new_n21290_ | new_n21308_);
  assign new_n21282_ = ~new_n21298_ & (new_n21301_ | (~new_n21302_ & (new_n21300_ | (~new_n21296_ & ~new_n21283_))));
  assign new_n21283_ = ~new_n21290_ & (~new_n21294_ | (new_n21284_ & (~new_n21293_ | (~new_n21295_ & new_n21287_))));
  assign new_n21284_ = \all_features[3183]  & (\all_features[3182]  | new_n21285_);
  assign new_n21285_ = \all_features[3181]  & (\all_features[3178]  | \all_features[3179]  | \all_features[3180]  | ~new_n21286_);
  assign new_n21286_ = ~\all_features[3176]  & ~\all_features[3177] ;
  assign new_n21287_ = \all_features[3183]  & ~new_n21288_ & \all_features[3182] ;
  assign new_n21288_ = ~\all_features[3181]  & ~\all_features[3180]  & ~\all_features[3179]  & ~new_n21289_ & ~\all_features[3178] ;
  assign new_n21289_ = \all_features[3176]  & \all_features[3177] ;
  assign new_n21290_ = ~\all_features[3183]  & (~\all_features[3182]  | ~new_n21289_ | ~new_n21291_ | ~new_n21292_);
  assign new_n21291_ = \all_features[3178]  & \all_features[3179] ;
  assign new_n21292_ = \all_features[3180]  & \all_features[3181] ;
  assign new_n21293_ = \all_features[3183]  & (\all_features[3182]  | (new_n21292_ & (\all_features[3178]  | \all_features[3179]  | \all_features[3177] )));
  assign new_n21294_ = \all_features[3183]  & (\all_features[3181]  | \all_features[3182]  | \all_features[3180] );
  assign new_n21295_ = \all_features[3182]  & \all_features[3183]  & (\all_features[3181]  | (\all_features[3180]  & (\all_features[3179]  | \all_features[3178] )));
  assign new_n21296_ = ~new_n21297_ & ~\all_features[3183] ;
  assign new_n21297_ = \all_features[3181]  & \all_features[3182]  & (\all_features[3180]  | (\all_features[3178]  & \all_features[3179]  & \all_features[3177] ));
  assign new_n21298_ = new_n21299_ & (~\all_features[3181]  | (~\all_features[3180]  & (~\all_features[3179]  | (~\all_features[3178]  & ~\all_features[3177] ))));
  assign new_n21299_ = ~\all_features[3182]  & ~\all_features[3183] ;
  assign new_n21300_ = ~\all_features[3183]  & (~\all_features[3182]  | (~\all_features[3181]  & (new_n21286_ | ~\all_features[3180]  | ~new_n21291_)));
  assign new_n21301_ = new_n21299_ & (~\all_features[3179]  | ~new_n21292_ | (~\all_features[3178]  & ~new_n21289_));
  assign new_n21302_ = ~\all_features[3183]  & (~\all_features[3182]  | (~\all_features[3180]  & ~\all_features[3181]  & ~new_n21291_));
  assign new_n21303_ = new_n21305_ & ~new_n21300_ & (new_n21296_ | new_n21290_ | new_n21304_ | new_n21302_);
  assign new_n21304_ = new_n21294_ & new_n21293_ & new_n21284_ & new_n21287_;
  assign new_n21305_ = ~new_n21307_ & ~new_n21302_ & ~new_n21306_ & ~new_n21298_ & ~new_n21301_;
  assign new_n21306_ = ~\all_features[3181]  & new_n21299_ & ((~\all_features[3178]  & new_n21286_) | ~\all_features[3180]  | ~\all_features[3179] );
  assign new_n21307_ = ~\all_features[3183]  & ~\all_features[3182]  & ~\all_features[3181]  & ~\all_features[3179]  & ~\all_features[3180] ;
  assign new_n21308_ = new_n21294_ & ~new_n21309_ & new_n21284_;
  assign new_n21309_ = ~new_n21288_ & new_n21293_ & \all_features[3182]  & \all_features[3183]  & (~\all_features[3181]  | new_n21310_);
  assign new_n21310_ = ~\all_features[3179]  & ~\all_features[3180]  & (~\all_features[3178]  | new_n21286_);
  assign new_n21311_ = ~new_n21302_ & ~new_n21306_ & ~new_n21300_ & ~new_n21301_;
  assign new_n21312_ = ~new_n21313_ & (\all_features[3835]  | \all_features[3836]  | \all_features[3837]  | \all_features[3838]  | \all_features[3839] );
  assign new_n21313_ = ~new_n21329_ & (new_n21333_ | (~new_n21332_ & (new_n21328_ | (~new_n21331_ & ~new_n21314_))));
  assign new_n21314_ = ~new_n21318_ & (new_n21320_ | (new_n21327_ & (~new_n21315_ | (~new_n21325_ & new_n21324_))));
  assign new_n21315_ = \all_features[3839]  & (\all_features[3838]  | new_n21316_);
  assign new_n21316_ = \all_features[3837]  & (\all_features[3834]  | \all_features[3835]  | \all_features[3836]  | ~new_n21317_);
  assign new_n21317_ = ~\all_features[3832]  & ~\all_features[3833] ;
  assign new_n21318_ = ~new_n21319_ & ~\all_features[3839] ;
  assign new_n21319_ = \all_features[3837]  & \all_features[3838]  & (\all_features[3836]  | (\all_features[3834]  & \all_features[3835]  & \all_features[3833] ));
  assign new_n21320_ = ~\all_features[3839]  & (~\all_features[3838]  | ~new_n21321_ | ~new_n21322_ | ~new_n21323_);
  assign new_n21321_ = \all_features[3832]  & \all_features[3833] ;
  assign new_n21322_ = \all_features[3834]  & \all_features[3835] ;
  assign new_n21323_ = \all_features[3836]  & \all_features[3837] ;
  assign new_n21324_ = \all_features[3839]  & (\all_features[3838]  | (new_n21323_ & (\all_features[3834]  | \all_features[3835]  | \all_features[3833] )));
  assign new_n21325_ = ~\all_features[3837]  & new_n21326_ & ((~\all_features[3836]  & (new_n21321_ | \all_features[3834]  | \all_features[3835] )) | (~\all_features[3834]  & ~\all_features[3835]  & \all_features[3836] ));
  assign new_n21326_ = \all_features[3838]  & \all_features[3839] ;
  assign new_n21327_ = \all_features[3839]  & (\all_features[3837]  | \all_features[3838]  | \all_features[3836] );
  assign new_n21328_ = ~\all_features[3839]  & (~\all_features[3838]  | (~\all_features[3836]  & ~\all_features[3837]  & ~new_n21322_));
  assign new_n21329_ = ~\all_features[3837]  & new_n21330_ & ((~\all_features[3834]  & new_n21317_) | ~\all_features[3836]  | ~\all_features[3835] );
  assign new_n21330_ = ~\all_features[3838]  & ~\all_features[3839] ;
  assign new_n21331_ = ~\all_features[3839]  & (~\all_features[3838]  | (~\all_features[3837]  & (new_n21317_ | ~\all_features[3836]  | ~new_n21322_)));
  assign new_n21332_ = new_n21330_ & (~\all_features[3835]  | ~new_n21323_ | (~\all_features[3834]  & ~new_n21321_));
  assign new_n21333_ = new_n21330_ & (~\all_features[3837]  | (~\all_features[3836]  & (~\all_features[3835]  | (~\all_features[3834]  & ~\all_features[3833] ))));
  assign new_n21334_ = new_n21342_ & (~new_n21339_ | (new_n21341_ & (~new_n21340_ | new_n21335_)));
  assign new_n21335_ = new_n21327_ & ~new_n21336_ & new_n21315_;
  assign new_n21336_ = new_n21337_ & new_n21324_ & (~\all_features[3837]  | ~new_n21326_ | new_n21338_);
  assign new_n21337_ = new_n21326_ & (new_n21321_ | \all_features[3834]  | \all_features[3835]  | \all_features[3836]  | \all_features[3837] );
  assign new_n21338_ = ~\all_features[3835]  & ~\all_features[3836]  & (~\all_features[3834]  | new_n21317_);
  assign new_n21339_ = ~new_n21332_ & ~new_n21333_;
  assign new_n21340_ = ~new_n21318_ & ~new_n21320_;
  assign new_n21341_ = ~new_n21328_ & ~new_n21331_;
  assign new_n21342_ = ~new_n21329_ & (\all_features[3835]  | \all_features[3836]  | \all_features[3837]  | \all_features[3838]  | \all_features[3839] );
  assign new_n21343_ = new_n21339_ & new_n21344_ & ~new_n21331_ & ~new_n21329_ & ~new_n21318_ & ~new_n21328_;
  assign new_n21344_ = ~new_n21320_ & (\all_features[3835]  | \all_features[3836]  | \all_features[3837]  | \all_features[3838]  | \all_features[3839] );
  assign new_n21345_ = new_n21342_ & new_n21339_ & (~new_n21341_ | ~new_n21340_ | (new_n21315_ & new_n21346_));
  assign new_n21346_ = new_n21327_ & new_n21324_ & new_n21337_;
  assign new_n21347_ = ~new_n21051_ & new_n20962_;
  assign new_n21348_ = new_n21355_ ? ((~new_n21353_ | new_n21389_) & (new_n21351_ | new_n21349_ | ~new_n21389_)) : ~new_n21390_;
  assign new_n21349_ = new_n21350_ & new_n9167_;
  assign new_n21350_ = ~new_n8292_ & (~new_n8269_ | new_n18100_);
  assign new_n21351_ = ~new_n9167_ & new_n11164_ & (new_n11161_ | new_n21352_);
  assign new_n21352_ = new_n11132_ & new_n11154_;
  assign new_n21353_ = ~new_n13806_ & (new_n17414_ | ~new_n21354_);
  assign new_n21354_ = ~new_n17392_ & ~new_n19644_;
  assign new_n21355_ = ~new_n21387_ & new_n21356_;
  assign new_n21356_ = ~new_n21357_ & ~new_n21382_;
  assign new_n21357_ = new_n21374_ & (new_n21381_ | new_n21380_ | (~new_n21378_ & ~new_n21379_ & ~new_n21358_));
  assign new_n21358_ = ~new_n21370_ & ~new_n21372_ & (~new_n21359_ | (~new_n21364_ & new_n21366_ & new_n21368_));
  assign new_n21359_ = new_n21360_ & new_n21363_;
  assign new_n21360_ = \all_features[5927]  & (\all_features[5926]  | (\all_features[5925]  & (\all_features[5924]  | ~new_n21362_ | ~new_n21361_)));
  assign new_n21361_ = ~\all_features[5922]  & ~\all_features[5923] ;
  assign new_n21362_ = ~\all_features[5920]  & ~\all_features[5921] ;
  assign new_n21363_ = \all_features[5927]  & (\all_features[5925]  | \all_features[5926]  | \all_features[5924] );
  assign new_n21364_ = \all_features[5927]  & \all_features[5926]  & ~new_n21365_ & \all_features[5925] ;
  assign new_n21365_ = ~\all_features[5923]  & ~\all_features[5924]  & (~\all_features[5922]  | new_n21362_);
  assign new_n21366_ = \all_features[5926]  & \all_features[5927]  & (\all_features[5924]  | \all_features[5925]  | new_n21367_ | ~new_n21361_);
  assign new_n21367_ = \all_features[5920]  & \all_features[5921] ;
  assign new_n21368_ = \all_features[5927]  & (\all_features[5926]  | (new_n21369_ & (\all_features[5922]  | \all_features[5923]  | \all_features[5921] )));
  assign new_n21369_ = \all_features[5924]  & \all_features[5925] ;
  assign new_n21370_ = ~new_n21371_ & ~\all_features[5927] ;
  assign new_n21371_ = \all_features[5925]  & \all_features[5926]  & (\all_features[5924]  | (\all_features[5922]  & \all_features[5923]  & \all_features[5921] ));
  assign new_n21372_ = ~\all_features[5927]  & (~\all_features[5926]  | ~new_n21367_ | ~new_n21369_ | ~new_n21373_);
  assign new_n21373_ = \all_features[5922]  & \all_features[5923] ;
  assign new_n21374_ = ~new_n21375_ & ~new_n21377_;
  assign new_n21375_ = ~\all_features[5925]  & new_n21376_ & ((~\all_features[5922]  & new_n21362_) | ~\all_features[5924]  | ~\all_features[5923] );
  assign new_n21376_ = ~\all_features[5926]  & ~\all_features[5927] ;
  assign new_n21377_ = ~\all_features[5927]  & ~\all_features[5926]  & ~\all_features[5925]  & ~\all_features[5923]  & ~\all_features[5924] ;
  assign new_n21378_ = ~\all_features[5927]  & (~\all_features[5926]  | (~\all_features[5925]  & (new_n21362_ | ~new_n21373_ | ~\all_features[5924] )));
  assign new_n21379_ = ~\all_features[5927]  & (~\all_features[5926]  | (~\all_features[5924]  & ~\all_features[5925]  & ~new_n21373_));
  assign new_n21380_ = new_n21376_ & (~\all_features[5925]  | (~\all_features[5924]  & (~\all_features[5923]  | (~\all_features[5922]  & ~\all_features[5921] ))));
  assign new_n21381_ = new_n21376_ & (~\all_features[5923]  | ~new_n21369_ | (~\all_features[5922]  & ~new_n21367_));
  assign new_n21382_ = ~new_n21377_ & (new_n21375_ | (~new_n21380_ & ~new_n21383_));
  assign new_n21383_ = ~new_n21381_ & (new_n21379_ | (~new_n21378_ & (new_n21370_ | (~new_n21372_ & ~new_n21384_))));
  assign new_n21384_ = new_n21363_ & (~new_n21360_ | (new_n21368_ & (new_n21385_ | ~new_n21366_)));
  assign new_n21385_ = \all_features[5926]  & \all_features[5927]  & (\all_features[5925]  | (~new_n21361_ & \all_features[5924] ));
  assign new_n21387_ = new_n21374_ & ~new_n21380_ & ~new_n21381_;
  assign new_n21388_ = ~new_n21379_ & ~new_n21372_ & ~new_n21378_ & ~new_n21370_;
  assign new_n21389_ = new_n8535_ & new_n18328_ & new_n8533_;
  assign new_n21390_ = new_n16562_ & (new_n16559_ | ~new_n21391_);
  assign new_n21391_ = ~new_n16529_ & ~new_n16550_;
  assign new_n21392_ = ~new_n20806_ & new_n20867_;
  assign new_n21393_ = new_n21394_ ? (~new_n21619_ ^ new_n21686_) : (new_n21619_ ^ new_n21686_);
  assign new_n21394_ = new_n21395_ ? (~new_n21565_ ^ new_n21600_) : (new_n21565_ ^ new_n21600_);
  assign new_n21395_ = new_n21396_ ? (~new_n21446_ ^ new_n21347_) : (new_n21446_ ^ new_n21347_);
  assign new_n21396_ = ~new_n21397_ & new_n21442_;
  assign new_n21397_ = ~new_n21398_ & ~new_n21435_ & new_n21408_ & (new_n21441_ | ~new_n21434_);
  assign new_n21398_ = new_n21399_ & (new_n8927_ ? new_n21400_ : ~new_n21407_);
  assign new_n21399_ = ~new_n13887_ & new_n20967_;
  assign new_n21400_ = ~new_n21401_ & new_n21406_;
  assign new_n21401_ = new_n19673_ & new_n21402_;
  assign new_n21402_ = ~new_n21403_ & (\all_features[2115]  | \all_features[2116]  | \all_features[2117]  | \all_features[2118]  | \all_features[2119] );
  assign new_n21403_ = ~new_n19654_ & (new_n19657_ | (~new_n19658_ & (new_n19667_ | (~new_n19662_ & ~new_n21404_))));
  assign new_n21404_ = ~new_n19664_ & (new_n19666_ | (new_n19672_ & (~new_n19668_ | (~new_n21405_ & new_n19670_))));
  assign new_n21405_ = ~\all_features[2117]  & \all_features[2118]  & \all_features[2119]  & (\all_features[2116]  ? new_n19669_ : (new_n19660_ | ~new_n19669_));
  assign new_n21406_ = ~new_n19651_ & ~new_n19677_;
  assign new_n21407_ = new_n14416_ & (new_n14394_ | new_n17766_);
  assign new_n21408_ = (~new_n21409_ | new_n21433_) & (new_n21412_ | new_n20967_ | ~new_n16659_);
  assign new_n21409_ = new_n20967_ & new_n13887_ & new_n21410_;
  assign new_n21410_ = new_n21411_ & new_n15157_;
  assign new_n21411_ = new_n11446_ & new_n11468_;
  assign new_n21412_ = (new_n21413_ & ~new_n18990_) | (new_n21414_ & new_n21422_ & new_n21430_ & new_n18990_);
  assign new_n21413_ = ~new_n14679_ & (~new_n14686_ | ~new_n14656_);
  assign new_n21414_ = ~new_n21415_ & (\all_features[5747]  | \all_features[5748]  | \all_features[5749]  | \all_features[5750]  | \all_features[5751] );
  assign new_n21415_ = ~new_n21178_ & (new_n21173_ | (~new_n21175_ & (new_n21180_ | (~new_n21181_ & ~new_n21416_))));
  assign new_n21416_ = ~new_n21176_ & (new_n21168_ | (new_n21421_ & (~new_n21417_ | (~new_n21420_ & new_n21419_))));
  assign new_n21417_ = \all_features[5751]  & (\all_features[5750]  | (\all_features[5749]  & (\all_features[5748]  | ~new_n21418_ | ~new_n21179_)));
  assign new_n21418_ = ~\all_features[5746]  & ~\all_features[5747] ;
  assign new_n21419_ = \all_features[5751]  & (\all_features[5750]  | (new_n21171_ & (\all_features[5746]  | \all_features[5747]  | \all_features[5745] )));
  assign new_n21420_ = ~\all_features[5749]  & \all_features[5750]  & \all_features[5751]  & (\all_features[5748]  ? new_n21418_ : (new_n21169_ | ~new_n21418_));
  assign new_n21421_ = \all_features[5751]  & (\all_features[5749]  | \all_features[5750]  | \all_features[5748] );
  assign new_n21422_ = new_n21429_ & (~new_n21172_ | (~new_n21423_ & new_n21428_));
  assign new_n21423_ = new_n21426_ & ((~new_n21424_ & new_n21419_ & new_n21427_) | ~new_n21421_ | ~new_n21417_);
  assign new_n21424_ = \all_features[5751]  & \all_features[5750]  & ~new_n21425_ & \all_features[5749] ;
  assign new_n21425_ = ~\all_features[5747]  & ~\all_features[5748]  & (~\all_features[5746]  | new_n21179_);
  assign new_n21426_ = ~new_n21176_ & ~new_n21168_;
  assign new_n21427_ = \all_features[5750]  & \all_features[5751]  & (\all_features[5748]  | \all_features[5749]  | new_n21169_ | ~new_n21418_);
  assign new_n21428_ = ~new_n21180_ & ~new_n21181_;
  assign new_n21429_ = ~new_n21178_ & (\all_features[5747]  | \all_features[5748]  | \all_features[5749]  | \all_features[5750]  | \all_features[5751] );
  assign new_n21430_ = new_n21166_ & new_n21431_;
  assign new_n21431_ = new_n21172_ & new_n21429_ & (~new_n21426_ | ~new_n21428_ | (new_n21432_ & new_n21417_));
  assign new_n21432_ = new_n21421_ & new_n21419_ & new_n21427_;
  assign new_n21433_ = new_n7513_ & (new_n7510_ | ~new_n12759_);
  assign new_n21434_ = new_n20967_ & ~new_n21410_ & new_n13887_;
  assign new_n21435_ = ~new_n16659_ & ~new_n20967_ & (new_n21436_ ? new_n16103_ : new_n14293_);
  assign new_n21436_ = new_n15086_ & (~new_n21437_ | (~new_n11807_ & (new_n11811_ | (~new_n21438_ & ~new_n11810_))));
  assign new_n21437_ = new_n11794_ & (\all_features[1443]  | \all_features[1444]  | \all_features[1445]  | \all_features[1446]  | \all_features[1447] );
  assign new_n21438_ = ~new_n11813_ & (new_n11815_ | (~new_n11818_ & (new_n11817_ | new_n21439_)));
  assign new_n21439_ = \all_features[1447]  & ((~new_n21440_ & \all_features[1446]  & new_n11802_) | (~new_n11800_ & ((~new_n21440_ & new_n11802_) | (~new_n11797_ & ~\all_features[1446] ))));
  assign new_n21440_ = ~\all_features[1445]  & \all_features[1446]  & \all_features[1447]  & (\all_features[1444]  ? new_n11799_ : (new_n11804_ | ~new_n11799_));
  assign new_n21441_ = ~new_n20790_ & new_n20118_;
  assign new_n21442_ = new_n21444_ & new_n21443_ & (~new_n21441_ | ~new_n21434_);
  assign new_n21443_ = (new_n21400_ | ~new_n21399_ | ~new_n8927_) & (~new_n21433_ | ~new_n21409_);
  assign new_n21444_ = (new_n21445_ | new_n20967_) & (new_n13887_ | new_n8927_ | ~new_n21407_ | ~new_n20967_);
  assign new_n21445_ = (new_n14293_ | new_n21436_ | new_n16659_) & (new_n18990_ | ~new_n21413_ | ~new_n16659_);
  assign new_n21446_ = new_n21447_ ? (new_n21488_ ^ new_n21532_) : (~new_n21488_ ^ new_n21532_);
  assign new_n21447_ = new_n21448_ & (~new_n17326_ | (~new_n21487_ & new_n6804_ & new_n10608_) | (~new_n21486_ & ~new_n10608_));
  assign new_n21448_ = (new_n21449_ | new_n17326_) & (new_n10608_ | new_n21485_ | ~new_n12408_ | ~new_n14810_ | ~new_n17326_);
  assign new_n21449_ = (~new_n21450_ | new_n6919_) & (new_n21484_ | new_n8097_ | ~new_n14883_);
  assign new_n21450_ = ~new_n14883_ & ~new_n21483_ & ~new_n21478_ & (new_n21471_ | new_n21480_ | ~new_n21451_);
  assign new_n21451_ = new_n21468_ & (~new_n21472_ | (~new_n21452_ & new_n21475_));
  assign new_n21452_ = new_n21453_ & ((~new_n21460_ & new_n21465_ & new_n21466_) | ~new_n21467_ | ~new_n21463_);
  assign new_n21453_ = ~new_n21454_ & ~new_n21456_;
  assign new_n21454_ = ~new_n21455_ & ~\all_features[1607] ;
  assign new_n21455_ = \all_features[1605]  & \all_features[1606]  & (\all_features[1604]  | (\all_features[1602]  & \all_features[1603]  & \all_features[1601] ));
  assign new_n21456_ = ~\all_features[1607]  & (~\all_features[1606]  | ~new_n21457_ | ~new_n21458_ | ~new_n21459_);
  assign new_n21457_ = \all_features[1600]  & \all_features[1601] ;
  assign new_n21458_ = \all_features[1604]  & \all_features[1605] ;
  assign new_n21459_ = \all_features[1602]  & \all_features[1603] ;
  assign new_n21460_ = \all_features[1607]  & \all_features[1606]  & ~new_n21461_ & \all_features[1605] ;
  assign new_n21461_ = ~\all_features[1603]  & ~\all_features[1604]  & (~\all_features[1602]  | new_n21462_);
  assign new_n21462_ = ~\all_features[1600]  & ~\all_features[1601] ;
  assign new_n21463_ = \all_features[1607]  & (\all_features[1606]  | (\all_features[1605]  & (\all_features[1604]  | ~new_n21464_ | ~new_n21462_)));
  assign new_n21464_ = ~\all_features[1602]  & ~\all_features[1603] ;
  assign new_n21465_ = \all_features[1607]  & (\all_features[1606]  | (new_n21458_ & (\all_features[1602]  | \all_features[1603]  | \all_features[1601] )));
  assign new_n21466_ = \all_features[1606]  & \all_features[1607]  & (\all_features[1604]  | \all_features[1605]  | new_n21457_ | ~new_n21464_);
  assign new_n21467_ = \all_features[1607]  & (\all_features[1605]  | \all_features[1606]  | \all_features[1604] );
  assign new_n21468_ = ~new_n21469_ & ~new_n21471_;
  assign new_n21469_ = ~\all_features[1605]  & new_n21470_ & ((~\all_features[1602]  & new_n21462_) | ~\all_features[1604]  | ~\all_features[1603] );
  assign new_n21470_ = ~\all_features[1606]  & ~\all_features[1607] ;
  assign new_n21471_ = ~\all_features[1607]  & ~\all_features[1606]  & ~\all_features[1605]  & ~\all_features[1603]  & ~\all_features[1604] ;
  assign new_n21472_ = ~new_n21473_ & ~new_n21474_;
  assign new_n21473_ = new_n21470_ & (~\all_features[1605]  | (~\all_features[1604]  & (~\all_features[1603]  | (~\all_features[1602]  & ~\all_features[1601] ))));
  assign new_n21474_ = new_n21470_ & (~\all_features[1603]  | ~new_n21458_ | (~\all_features[1602]  & ~new_n21457_));
  assign new_n21475_ = ~new_n21476_ & ~new_n21477_;
  assign new_n21476_ = ~\all_features[1607]  & (~\all_features[1606]  | (~\all_features[1604]  & ~\all_features[1605]  & ~new_n21459_));
  assign new_n21477_ = ~\all_features[1607]  & (~\all_features[1606]  | (~\all_features[1605]  & (new_n21462_ | ~new_n21459_ | ~\all_features[1604] )));
  assign new_n21478_ = ~new_n21471_ & ~new_n21474_ & ~new_n21473_ & ~new_n21479_ & ~new_n21469_;
  assign new_n21479_ = new_n21475_ & new_n21453_ & (~new_n21466_ | ~new_n21467_ | ~new_n21463_ | ~new_n21465_);
  assign new_n21480_ = ~new_n21469_ & (new_n21473_ | (~new_n21474_ & (new_n21476_ | (~new_n21481_ & ~new_n21477_))));
  assign new_n21481_ = ~new_n21454_ & (new_n21456_ | (new_n21467_ & (~new_n21463_ | (~new_n21482_ & new_n21465_))));
  assign new_n21482_ = ~\all_features[1605]  & \all_features[1606]  & \all_features[1607]  & (\all_features[1604]  ? new_n21464_ : (new_n21457_ | ~new_n21464_));
  assign new_n21483_ = new_n21472_ & new_n21468_ & ~new_n21456_ & ~new_n21454_ & ~new_n21476_ & ~new_n21477_;
  assign new_n21484_ = new_n9100_ & new_n16648_;
  assign new_n21485_ = ~new_n14787_ & ~new_n18086_;
  assign new_n21486_ = ~new_n12408_ & (~new_n16455_ | new_n19426_);
  assign new_n21487_ = ~new_n7104_ & ~new_n7126_;
  assign new_n21488_ = ~new_n21489_ & ~new_n21531_;
  assign new_n21489_ = ~new_n21528_ & new_n21490_;
  assign new_n21490_ = new_n21527_ ? ((new_n21525_ & new_n17388_ & ~new_n21492_) | (new_n21491_ & new_n21492_)) : new_n20851_;
  assign new_n21491_ = ~new_n15674_ & (new_n14545_ | ~new_n15828_);
  assign new_n21492_ = ~new_n21493_ & new_n21524_;
  assign new_n21493_ = ~new_n21494_ & ~new_n21521_;
  assign new_n21494_ = new_n21506_ & (~new_n21510_ | (new_n21513_ & (~new_n21517_ | new_n21495_)));
  assign new_n21495_ = new_n21496_ & (~new_n21500_ | (~new_n21505_ & \all_features[1269]  & \all_features[1270]  & \all_features[1271] ));
  assign new_n21496_ = \all_features[1271]  & (\all_features[1270]  | (~new_n21497_ & \all_features[1269] ));
  assign new_n21497_ = new_n21498_ & ~\all_features[1268]  & new_n21499_;
  assign new_n21498_ = ~\all_features[1264]  & ~\all_features[1265] ;
  assign new_n21499_ = ~\all_features[1266]  & ~\all_features[1267] ;
  assign new_n21500_ = \all_features[1271]  & \all_features[1270]  & ~new_n21503_ & new_n21501_;
  assign new_n21501_ = \all_features[1271]  & (\all_features[1270]  | (new_n21502_ & (\all_features[1266]  | \all_features[1267]  | \all_features[1265] )));
  assign new_n21502_ = \all_features[1268]  & \all_features[1269] ;
  assign new_n21503_ = new_n21499_ & ~\all_features[1269]  & ~new_n21504_ & ~\all_features[1268] ;
  assign new_n21504_ = \all_features[1264]  & \all_features[1265] ;
  assign new_n21505_ = ~\all_features[1267]  & ~\all_features[1268]  & (~\all_features[1266]  | new_n21498_);
  assign new_n21506_ = ~new_n21507_ & ~new_n21509_;
  assign new_n21507_ = ~\all_features[1269]  & new_n21508_ & ((~\all_features[1266]  & new_n21498_) | ~\all_features[1268]  | ~\all_features[1267] );
  assign new_n21508_ = ~\all_features[1270]  & ~\all_features[1271] ;
  assign new_n21509_ = ~\all_features[1271]  & ~\all_features[1270]  & ~\all_features[1269]  & ~\all_features[1267]  & ~\all_features[1268] ;
  assign new_n21510_ = ~new_n21511_ & ~new_n21512_;
  assign new_n21511_ = new_n21508_ & (~\all_features[1267]  | ~new_n21502_ | (~\all_features[1266]  & ~new_n21504_));
  assign new_n21512_ = new_n21508_ & (~\all_features[1269]  | (~\all_features[1268]  & (~\all_features[1267]  | (~\all_features[1266]  & ~\all_features[1265] ))));
  assign new_n21513_ = ~new_n21514_ & ~new_n21516_;
  assign new_n21514_ = ~\all_features[1271]  & (~\all_features[1270]  | (~\all_features[1268]  & ~\all_features[1269]  & ~new_n21515_));
  assign new_n21515_ = \all_features[1266]  & \all_features[1267] ;
  assign new_n21516_ = ~\all_features[1271]  & (~\all_features[1270]  | (~\all_features[1269]  & (new_n21498_ | ~new_n21515_ | ~\all_features[1268] )));
  assign new_n21517_ = ~new_n21518_ & ~new_n21519_;
  assign new_n21518_ = ~\all_features[1271]  & (~\all_features[1270]  | ~new_n21504_ | ~new_n21502_ | ~new_n21515_);
  assign new_n21519_ = ~new_n21520_ & ~\all_features[1271] ;
  assign new_n21520_ = \all_features[1269]  & \all_features[1270]  & (\all_features[1268]  | (\all_features[1266]  & \all_features[1267]  & \all_features[1265] ));
  assign new_n21521_ = new_n21522_ & (new_n21516_ | new_n21519_ | ~new_n21523_ | (new_n21500_ & new_n21496_));
  assign new_n21522_ = new_n21506_ & new_n21510_;
  assign new_n21523_ = ~new_n21514_ & ~new_n21518_;
  assign new_n21524_ = new_n21517_ & new_n21522_ & new_n21513_;
  assign new_n21525_ = ~new_n7832_ & (~new_n7830_ | ~new_n21526_);
  assign new_n21526_ = new_n7805_ & new_n16901_;
  assign new_n21527_ = new_n13409_ & new_n13437_;
  assign new_n21528_ = ~new_n21527_ & new_n20851_ & (new_n21529_ | (new_n14042_ & (new_n14039_ | ~new_n20114_)));
  assign new_n21529_ = new_n21530_ & ~new_n8705_ & ~new_n8725_;
  assign new_n21530_ = ~new_n8736_ & ~new_n8739_;
  assign new_n21531_ = new_n17388_ & new_n21527_ & ~new_n21492_ & new_n21525_;
  assign new_n21532_ = new_n21561_ ? new_n21533_ : ((new_n21563_ & new_n19702_) ? new_n21560_ : new_n21564_);
  assign new_n21533_ = (~new_n16190_ & (~new_n16158_ | ~new_n16188_)) ? new_n21534_ : ~new_n20787_;
  assign new_n21534_ = new_n21535_ ? new_n21536_ : (~new_n17480_ | (new_n17472_ & new_n17485_));
  assign new_n21535_ = ~new_n6908_ & (~new_n6910_ | ~new_n6886_);
  assign new_n21536_ = ~new_n21537_ & ~new_n21559_;
  assign new_n21537_ = new_n21538_ & (~new_n21547_ | (new_n21557_ & new_n21558_ & new_n21554_ & new_n21556_));
  assign new_n21538_ = new_n21539_ & ~new_n21543_ & ~new_n21544_;
  assign new_n21539_ = ~new_n21540_ & (\all_features[4635]  | \all_features[4636]  | \all_features[4637]  | \all_features[4638]  | \all_features[4639] );
  assign new_n21540_ = ~\all_features[4637]  & new_n21542_ & ((~\all_features[4634]  & new_n21541_) | ~\all_features[4636]  | ~\all_features[4635] );
  assign new_n21541_ = ~\all_features[4632]  & ~\all_features[4633] ;
  assign new_n21542_ = ~\all_features[4638]  & ~\all_features[4639] ;
  assign new_n21543_ = new_n21542_ & (~\all_features[4637]  | (~\all_features[4636]  & (~\all_features[4635]  | (~\all_features[4634]  & ~\all_features[4633] ))));
  assign new_n21544_ = new_n21542_ & (~\all_features[4635]  | ~new_n21545_ | (~\all_features[4634]  & ~new_n21546_));
  assign new_n21545_ = \all_features[4636]  & \all_features[4637] ;
  assign new_n21546_ = \all_features[4632]  & \all_features[4633] ;
  assign new_n21547_ = ~new_n21553_ & ~new_n21552_ & ~new_n21548_ & ~new_n21550_;
  assign new_n21548_ = ~\all_features[4639]  & (~\all_features[4638]  | (~\all_features[4637]  & (new_n21541_ | ~new_n21549_ | ~\all_features[4636] )));
  assign new_n21549_ = \all_features[4634]  & \all_features[4635] ;
  assign new_n21550_ = ~new_n21551_ & ~\all_features[4639] ;
  assign new_n21551_ = \all_features[4637]  & \all_features[4638]  & (\all_features[4636]  | (\all_features[4634]  & \all_features[4635]  & \all_features[4633] ));
  assign new_n21552_ = ~\all_features[4639]  & (~\all_features[4638]  | ~new_n21545_ | ~new_n21546_ | ~new_n21549_);
  assign new_n21553_ = ~\all_features[4639]  & (~\all_features[4638]  | (~\all_features[4636]  & ~\all_features[4637]  & ~new_n21549_));
  assign new_n21554_ = \all_features[4639]  & (\all_features[4638]  | (\all_features[4637]  & (\all_features[4636]  | ~new_n21541_ | ~new_n21555_)));
  assign new_n21555_ = ~\all_features[4634]  & ~\all_features[4635] ;
  assign new_n21556_ = \all_features[4639]  & (\all_features[4638]  | (new_n21545_ & (\all_features[4634]  | \all_features[4635]  | \all_features[4633] )));
  assign new_n21557_ = \all_features[4638]  & \all_features[4639]  & (\all_features[4636]  | \all_features[4637]  | new_n21546_ | ~new_n21555_);
  assign new_n21558_ = \all_features[4639]  & (\all_features[4637]  | \all_features[4638]  | \all_features[4636] );
  assign new_n21559_ = new_n21538_ & new_n21547_;
  assign new_n21560_ = new_n16565_ & new_n13095_ & (new_n13067_ | ~new_n13517_);
  assign new_n21561_ = new_n19534_ & new_n21562_ & new_n19510_;
  assign new_n21562_ = new_n19538_ & new_n19541_;
  assign new_n21563_ = ~new_n19720_ & new_n19679_;
  assign new_n21564_ = (new_n20978_ & new_n21001_ & ~new_n18893_) | (~new_n16101_ & new_n18893_ & (~new_n16098_ | ~new_n16067_));
  assign new_n21565_ = ~new_n21566_ & new_n21597_;
  assign new_n21566_ = ~new_n21567_ & new_n21587_ & (~new_n21586_ | (~new_n19197_ & new_n20579_));
  assign new_n21567_ = new_n21568_ & (new_n21571_ ? new_n21572_ : ~new_n21569_);
  assign new_n21568_ = new_n9725_ & new_n20695_;
  assign new_n21569_ = ~new_n21211_ & new_n21570_;
  assign new_n21570_ = new_n21242_ & new_n21245_;
  assign new_n21571_ = ~new_n8619_ & (~new_n8622_ | ~new_n8626_ | ~new_n8596_);
  assign new_n21572_ = new_n13329_ & new_n21573_ & new_n21584_;
  assign new_n21573_ = new_n21583_ & (~new_n13336_ | (~new_n21574_ & ~new_n13342_ & ~new_n13345_));
  assign new_n21574_ = ~new_n13340_ & ~new_n13331_ & (~new_n21575_ | (~new_n21578_ & new_n21580_));
  assign new_n21575_ = \all_features[1735]  & (\all_features[1734]  | (~new_n21576_ & \all_features[1733] ));
  assign new_n21576_ = new_n13344_ & ~\all_features[1732]  & new_n21577_;
  assign new_n21577_ = ~\all_features[1730]  & ~\all_features[1731] ;
  assign new_n21578_ = \all_features[1735]  & \all_features[1734]  & ~new_n21579_ & \all_features[1733] ;
  assign new_n21579_ = ~\all_features[1731]  & ~\all_features[1732]  & (~\all_features[1730]  | new_n13344_);
  assign new_n21580_ = \all_features[1735]  & \all_features[1734]  & ~new_n21582_ & new_n21581_;
  assign new_n21581_ = \all_features[1735]  & (\all_features[1734]  | (new_n13333_ & (\all_features[1730]  | \all_features[1731]  | \all_features[1729] )));
  assign new_n21582_ = new_n21577_ & ~\all_features[1733]  & ~new_n13332_ & ~\all_features[1732] ;
  assign new_n21583_ = ~new_n13343_ & ~new_n13335_;
  assign new_n21584_ = new_n21583_ & ~new_n21585_ & new_n13336_;
  assign new_n21585_ = ~new_n13340_ & ~new_n13331_ & ~new_n13342_ & ~new_n13345_ & (~new_n21580_ | ~new_n21575_);
  assign new_n21586_ = ~new_n9725_ & new_n20695_;
  assign new_n21587_ = new_n20695_ | ((~new_n21590_ | ~new_n21596_ | new_n21589_) & (new_n21588_ | ~new_n19719_ | ~new_n21589_));
  assign new_n21588_ = ~new_n12798_ & (~new_n14920_ | ~new_n12793_);
  assign new_n21589_ = new_n10455_ & new_n10481_;
  assign new_n21590_ = new_n21591_ & ~new_n13758_ & ~new_n21592_;
  assign new_n21591_ = ~new_n13736_ & ~new_n13765_;
  assign new_n21592_ = ~new_n21593_ & (\all_features[5547]  | \all_features[5548]  | \all_features[5549]  | \all_features[5550]  | \all_features[5551] );
  assign new_n21593_ = ~new_n13754_ & (new_n13756_ | (~new_n13757_ & (new_n13747_ | (~new_n13739_ & ~new_n21594_))));
  assign new_n21594_ = ~new_n13742_ & (new_n13744_ | (new_n13752_ & (~new_n13748_ | (~new_n21595_ & new_n13750_))));
  assign new_n21595_ = ~\all_features[5549]  & \all_features[5550]  & \all_features[5551]  & (\all_features[5548]  ? new_n13749_ : (new_n13746_ | ~new_n13749_));
  assign new_n21596_ = ~new_n19704_ & ~new_n8188_;
  assign new_n21597_ = new_n21598_ & (~new_n21568_ | (new_n21572_ & new_n21571_) | (~new_n21569_ & ~new_n21571_));
  assign new_n21598_ = ~new_n21599_ & (new_n19197_ | ~new_n20579_ | ~new_n21586_);
  assign new_n21599_ = ~new_n20695_ & (new_n21589_ ? (new_n21588_ | ~new_n19719_) : ~new_n21590_);
  assign new_n21600_ = (new_n21603_ | ~new_n21617_) & (new_n21601_ | ~new_n16997_ | ~new_n21616_ | new_n21617_);
  assign new_n21601_ = ~new_n6532_ | (~new_n6529_ & new_n21602_);
  assign new_n21602_ = ~new_n6499_ & ~new_n6521_;
  assign new_n21603_ = new_n21614_ ? ~new_n21604_ : (new_n21615_ | (~new_n14848_ & new_n7987_));
  assign new_n21604_ = ~new_n18385_ & (~new_n21610_ | ~new_n21605_);
  assign new_n21605_ = new_n10308_ & new_n10285_ & new_n21606_;
  assign new_n21606_ = new_n10303_ & (~new_n10309_ | (~new_n21607_ & ~new_n10297_ & ~new_n10301_));
  assign new_n21607_ = ~new_n10302_ & ~new_n10295_ & (~new_n10293_ | ~new_n10299_ | new_n21608_);
  assign new_n21608_ = new_n10288_ & new_n10290_ & (new_n21609_ | ~\all_features[5469]  | ~\all_features[5470]  | ~\all_features[5471] );
  assign new_n21609_ = ~\all_features[5467]  & ~\all_features[5468]  & (~\all_features[5466]  | new_n10300_);
  assign new_n21610_ = ~new_n21611_ & (\all_features[5467]  | \all_features[5468]  | \all_features[5469]  | \all_features[5470]  | \all_features[5471] );
  assign new_n21611_ = ~new_n10304_ & (new_n10306_ | (~new_n10307_ & (new_n10297_ | (~new_n10301_ & ~new_n21612_))));
  assign new_n21612_ = ~new_n10295_ & (new_n10302_ | (new_n10293_ & (~new_n10299_ | (~new_n21613_ & new_n10288_))));
  assign new_n21613_ = ~\all_features[5469]  & \all_features[5470]  & \all_features[5471]  & (\all_features[5468]  ? new_n10291_ : (new_n10292_ | ~new_n10291_));
  assign new_n21614_ = ~new_n8344_ & (~new_n8346_ | ~new_n10774_);
  assign new_n21615_ = new_n13368_ & (~new_n13397_ | ~new_n13393_);
  assign new_n21616_ = ~new_n6591_ & (~new_n6569_ | ~new_n6592_);
  assign new_n21617_ = new_n15702_ & (new_n15676_ | new_n21618_);
  assign new_n21618_ = new_n15703_ & new_n17850_;
  assign new_n21619_ = ~new_n21620_ & new_n21681_;
  assign new_n21620_ = new_n21621_ & new_n21674_;
  assign new_n21621_ = ~new_n21622_ & (~new_n20844_ | ((new_n21640_ | ~new_n11824_) & (new_n21638_ | ~new_n21639_ | new_n11824_)));
  assign new_n21622_ = new_n21623_ & new_n21624_ & (new_n15315_ | ~new_n15283_);
  assign new_n21623_ = ~new_n18175_ & ~new_n20844_;
  assign new_n21624_ = ~new_n21625_ & new_n15265_;
  assign new_n21625_ = ~new_n21626_ & ~new_n21636_;
  assign new_n21626_ = new_n21635_ & (~new_n15271_ | (~new_n21627_ & ~new_n15269_ & ~new_n15280_));
  assign new_n21627_ = ~new_n15275_ & ~new_n15279_ & (~new_n21628_ | (~new_n21630_ & new_n21632_));
  assign new_n21628_ = \all_features[1047]  & (\all_features[1046]  | (~new_n21629_ & \all_features[1045] ));
  assign new_n21629_ = new_n15278_ & ~\all_features[1044]  & ~\all_features[1042]  & ~\all_features[1043] ;
  assign new_n21630_ = \all_features[1047]  & \all_features[1046]  & ~new_n21631_ & \all_features[1045] ;
  assign new_n21631_ = ~\all_features[1043]  & ~\all_features[1044]  & (~\all_features[1042]  | new_n15278_);
  assign new_n21632_ = \all_features[1047]  & \all_features[1046]  & ~new_n21634_ & new_n21633_;
  assign new_n21633_ = \all_features[1047]  & (\all_features[1046]  | (new_n15273_ & (\all_features[1042]  | \all_features[1043]  | \all_features[1041] )));
  assign new_n21634_ = ~\all_features[1042]  & ~\all_features[1043]  & ~\all_features[1044]  & ~\all_features[1045]  & (~\all_features[1041]  | ~\all_features[1040] );
  assign new_n21635_ = ~new_n15267_ & ~new_n15277_;
  assign new_n21636_ = new_n21635_ & ~new_n21637_ & new_n15271_;
  assign new_n21637_ = ~new_n15275_ & ~new_n15269_ & ~new_n15279_ & ~new_n15280_ & (~new_n21632_ | ~new_n21628_);
  assign new_n21638_ = new_n20464_ & (~new_n20478_ | ~new_n20474_);
  assign new_n21639_ = ~new_n16269_ & new_n14626_;
  assign new_n21640_ = ~new_n14985_ & new_n21641_;
  assign new_n21641_ = ~new_n21642_ & new_n21669_;
  assign new_n21642_ = ~new_n21668_ & (~new_n21661_ | (~new_n21666_ & (new_n21659_ | new_n21667_ | ~new_n21643_)));
  assign new_n21643_ = ~new_n21655_ & ~new_n21653_ & ((~new_n21650_ & new_n21644_) | ~new_n21658_ | ~new_n21657_);
  assign new_n21644_ = \all_features[3967]  & \all_features[3966]  & ~new_n21647_ & new_n21645_;
  assign new_n21645_ = \all_features[3967]  & (\all_features[3966]  | (new_n21646_ & (\all_features[3962]  | \all_features[3963]  | \all_features[3961] )));
  assign new_n21646_ = \all_features[3964]  & \all_features[3965] ;
  assign new_n21647_ = new_n21649_ & ~\all_features[3965]  & ~new_n21648_ & ~\all_features[3964] ;
  assign new_n21648_ = \all_features[3960]  & \all_features[3961] ;
  assign new_n21649_ = ~\all_features[3962]  & ~\all_features[3963] ;
  assign new_n21650_ = \all_features[3967]  & \all_features[3966]  & ~new_n21651_ & \all_features[3965] ;
  assign new_n21651_ = ~\all_features[3963]  & ~\all_features[3964]  & (~\all_features[3962]  | new_n21652_);
  assign new_n21652_ = ~\all_features[3960]  & ~\all_features[3961] ;
  assign new_n21653_ = ~new_n21654_ & ~\all_features[3967] ;
  assign new_n21654_ = \all_features[3965]  & \all_features[3966]  & (\all_features[3964]  | (\all_features[3962]  & \all_features[3963]  & \all_features[3961] ));
  assign new_n21655_ = ~\all_features[3967]  & (~\all_features[3966]  | ~new_n21656_ | ~new_n21648_ | ~new_n21646_);
  assign new_n21656_ = \all_features[3962]  & \all_features[3963] ;
  assign new_n21657_ = \all_features[3967]  & (\all_features[3966]  | (\all_features[3965]  & (\all_features[3964]  | ~new_n21649_ | ~new_n21652_)));
  assign new_n21658_ = \all_features[3967]  & (\all_features[3965]  | \all_features[3966]  | \all_features[3964] );
  assign new_n21659_ = ~new_n21653_ & (new_n21655_ | (new_n21658_ & (~new_n21657_ | (~new_n21660_ & new_n21645_))));
  assign new_n21660_ = ~\all_features[3965]  & \all_features[3966]  & \all_features[3967]  & (\all_features[3964]  ? new_n21649_ : (new_n21648_ | ~new_n21649_));
  assign new_n21661_ = ~new_n21665_ & ~new_n21662_ & ~new_n21664_;
  assign new_n21662_ = new_n21663_ & (~\all_features[3965]  | (~\all_features[3964]  & (~\all_features[3963]  | (~\all_features[3962]  & ~\all_features[3961] ))));
  assign new_n21663_ = ~\all_features[3966]  & ~\all_features[3967] ;
  assign new_n21664_ = ~\all_features[3965]  & new_n21663_ & ((~\all_features[3962]  & new_n21652_) | ~\all_features[3964]  | ~\all_features[3963] );
  assign new_n21665_ = new_n21663_ & (~\all_features[3963]  | ~new_n21646_ | (~\all_features[3962]  & ~new_n21648_));
  assign new_n21666_ = ~\all_features[3967]  & (~\all_features[3966]  | (~\all_features[3964]  & ~\all_features[3965]  & ~new_n21656_));
  assign new_n21667_ = ~\all_features[3967]  & (~\all_features[3966]  | (~\all_features[3965]  & (new_n21652_ | ~\all_features[3964]  | ~new_n21656_)));
  assign new_n21668_ = ~\all_features[3967]  & ~\all_features[3966]  & ~\all_features[3965]  & ~\all_features[3963]  & ~\all_features[3964] ;
  assign new_n21669_ = new_n21662_ | ~new_n21672_ | ((new_n21653_ | ~new_n21673_) & (new_n21670_ | new_n21665_));
  assign new_n21670_ = new_n21671_ & (~new_n21644_ | ~new_n21657_ | ~new_n21658_);
  assign new_n21671_ = ~new_n21655_ & ~new_n21653_ & ~new_n21666_ & ~new_n21667_;
  assign new_n21672_ = ~new_n21664_ & ~new_n21668_;
  assign new_n21673_ = ~new_n21665_ & ~new_n21655_ & ~new_n21666_ & ~new_n21667_;
  assign new_n21674_ = (~new_n21680_ | ~new_n21675_) & (~new_n21676_ | (new_n21678_ ? ~new_n21677_ : ~new_n21679_));
  assign new_n21675_ = ~new_n21624_ & new_n21623_;
  assign new_n21676_ = ~new_n20844_ & new_n18175_;
  assign new_n21677_ = new_n19584_ & (new_n19581_ | ~new_n19552_);
  assign new_n21678_ = ~new_n20838_ & ~new_n20812_ & ~new_n20842_;
  assign new_n21679_ = new_n20977_ & (~new_n21007_ | ~new_n21003_);
  assign new_n21680_ = new_n17734_ & (new_n21194_ | new_n21190_ | new_n17711_);
  assign new_n21681_ = new_n21682_ & new_n21683_;
  assign new_n21682_ = (~new_n21675_ | new_n21680_) & (~new_n21676_ | (new_n21678_ ? new_n21677_ : new_n21679_));
  assign new_n21683_ = ~new_n20844_ | (new_n11824_ ? ~new_n21640_ : (new_n21639_ ? ~new_n21638_ : new_n21684_));
  assign new_n21684_ = new_n12304_ & new_n21685_;
  assign new_n21685_ = ~new_n12334_ & ~new_n12337_;
  assign new_n21686_ = new_n21687_ & (~new_n21697_ | ~new_n21696_);
  assign new_n21687_ = new_n21688_ & (~new_n21691_ | (~new_n12190_ & new_n21695_) | (new_n21692_ & ~new_n21695_));
  assign new_n21688_ = new_n21689_ | ((new_n12228_ | new_n8225_ | new_n15592_) & (~new_n15592_ | (~new_n21690_ & ~new_n16758_)));
  assign new_n21689_ = ~new_n20474_ & new_n20464_;
  assign new_n21690_ = ~new_n19737_ & new_n19766_;
  assign new_n21691_ = ~new_n17415_ & new_n21689_;
  assign new_n21692_ = ~new_n19384_ & new_n21693_;
  assign new_n21693_ = ~new_n19405_ & new_n21694_;
  assign new_n21694_ = ~new_n19412_ & ~new_n19414_;
  assign new_n21695_ = ~new_n13158_ & (~new_n13136_ | new_n13159_);
  assign new_n21696_ = new_n21689_ & new_n17415_;
  assign new_n21697_ = new_n12373_ ? new_n19767_ : ~new_n11025_;
  assign new_n21698_ = ~new_n21699_ & new_n21757_;
  assign new_n21699_ = ~new_n21721_ & new_n21700_ & (~new_n21755_ | (~new_n16810_ & new_n19883_) | (new_n21756_ & ~new_n19883_));
  assign new_n21700_ = (~new_n21714_ | ~new_n17709_) & (new_n16758_ | ~new_n21701_);
  assign new_n21701_ = new_n21705_ & ~new_n21704_ & new_n21702_;
  assign new_n21702_ = ~new_n21703_ & ~new_n11201_;
  assign new_n21703_ = ~new_n14279_ & new_n11199_;
  assign new_n21704_ = new_n7869_ & new_n16647_;
  assign new_n21705_ = new_n21706_ & (new_n20221_ | (~new_n21711_ & ~new_n20219_));
  assign new_n21706_ = ~new_n20232_ & ~new_n20207_ & (~new_n20218_ | new_n21707_);
  assign new_n21707_ = new_n20226_ & (new_n20225_ | new_n20231_ | (~new_n20229_ & ~new_n21708_ & ~new_n20223_));
  assign new_n21708_ = new_n20217_ & ~new_n21709_ & new_n20209_;
  assign new_n21709_ = ~new_n20213_ & new_n20215_ & \all_features[1006]  & \all_features[1007]  & (~\all_features[1005]  | new_n21710_);
  assign new_n21710_ = ~\all_features[1003]  & ~\all_features[1004]  & (~\all_features[1002]  | new_n20211_);
  assign new_n21711_ = ~new_n20227_ & (new_n20228_ | (~new_n20225_ & (new_n20231_ | (~new_n20229_ & ~new_n21712_))));
  assign new_n21712_ = ~new_n20223_ & (~new_n20217_ | (new_n20209_ & (~new_n20215_ | (~new_n21713_ & new_n20212_))));
  assign new_n21713_ = \all_features[1006]  & \all_features[1007]  & (\all_features[1005]  | (\all_features[1004]  & (\all_features[1003]  | \all_features[1002] )));
  assign new_n21714_ = new_n21716_ & ~new_n21702_ & new_n21715_;
  assign new_n21715_ = ~new_n12001_ & (~new_n14086_ | ~new_n17935_);
  assign new_n21716_ = ~new_n21717_ & new_n19469_;
  assign new_n21717_ = ~new_n21718_ & (\all_features[2275]  | \all_features[2276]  | \all_features[2277]  | \all_features[2278]  | \all_features[2279] );
  assign new_n21718_ = ~new_n19486_ & (new_n19492_ | (~new_n19491_ & (new_n19493_ | (~new_n19488_ & ~new_n21719_))));
  assign new_n21719_ = ~new_n19482_ & (new_n19481_ | (new_n19484_ & (~new_n19480_ | (~new_n21720_ & new_n19473_))));
  assign new_n21720_ = ~\all_features[2277]  & \all_features[2278]  & \all_features[2279]  & (\all_features[2276]  ? new_n19478_ : (new_n19479_ | ~new_n19478_));
  assign new_n21721_ = new_n21702_ & (new_n21704_ ? (new_n21722_ ? ~new_n19767_ : new_n14038_) : ~new_n21705_);
  assign new_n21722_ = ~new_n21723_ & new_n21750_;
  assign new_n21723_ = ~new_n21749_ & (~new_n21742_ | (~new_n21747_ & (new_n21740_ | new_n21748_ | ~new_n21724_)));
  assign new_n21724_ = ~new_n21736_ & ~new_n21734_ & ((~new_n21731_ & new_n21725_) | ~new_n21739_ | ~new_n21738_);
  assign new_n21725_ = \all_features[1175]  & \all_features[1174]  & ~new_n21728_ & new_n21726_;
  assign new_n21726_ = \all_features[1175]  & (\all_features[1174]  | (new_n21727_ & (\all_features[1170]  | \all_features[1171]  | \all_features[1169] )));
  assign new_n21727_ = \all_features[1172]  & \all_features[1173] ;
  assign new_n21728_ = new_n21730_ & ~\all_features[1173]  & ~new_n21729_ & ~\all_features[1172] ;
  assign new_n21729_ = \all_features[1168]  & \all_features[1169] ;
  assign new_n21730_ = ~\all_features[1170]  & ~\all_features[1171] ;
  assign new_n21731_ = \all_features[1175]  & \all_features[1174]  & ~new_n21732_ & \all_features[1173] ;
  assign new_n21732_ = ~\all_features[1171]  & ~\all_features[1172]  & (~\all_features[1170]  | new_n21733_);
  assign new_n21733_ = ~\all_features[1168]  & ~\all_features[1169] ;
  assign new_n21734_ = ~new_n21735_ & ~\all_features[1175] ;
  assign new_n21735_ = \all_features[1173]  & \all_features[1174]  & (\all_features[1172]  | (\all_features[1170]  & \all_features[1171]  & \all_features[1169] ));
  assign new_n21736_ = ~\all_features[1175]  & (~\all_features[1174]  | ~new_n21737_ | ~new_n21729_ | ~new_n21727_);
  assign new_n21737_ = \all_features[1170]  & \all_features[1171] ;
  assign new_n21738_ = \all_features[1175]  & (\all_features[1174]  | (\all_features[1173]  & (\all_features[1172]  | ~new_n21730_ | ~new_n21733_)));
  assign new_n21739_ = \all_features[1175]  & (\all_features[1173]  | \all_features[1174]  | \all_features[1172] );
  assign new_n21740_ = ~new_n21734_ & (new_n21736_ | (new_n21739_ & (~new_n21738_ | (~new_n21741_ & new_n21726_))));
  assign new_n21741_ = ~\all_features[1173]  & \all_features[1174]  & \all_features[1175]  & (\all_features[1172]  ? new_n21730_ : (new_n21729_ | ~new_n21730_));
  assign new_n21742_ = ~new_n21746_ & ~new_n21743_ & ~new_n21745_;
  assign new_n21743_ = new_n21744_ & (~\all_features[1173]  | (~\all_features[1172]  & (~\all_features[1171]  | (~\all_features[1170]  & ~\all_features[1169] ))));
  assign new_n21744_ = ~\all_features[1174]  & ~\all_features[1175] ;
  assign new_n21745_ = ~\all_features[1173]  & new_n21744_ & ((~\all_features[1170]  & new_n21733_) | ~\all_features[1172]  | ~\all_features[1171] );
  assign new_n21746_ = new_n21744_ & (~\all_features[1171]  | ~new_n21727_ | (~\all_features[1170]  & ~new_n21729_));
  assign new_n21747_ = ~\all_features[1175]  & (~\all_features[1174]  | (~\all_features[1172]  & ~\all_features[1173]  & ~new_n21737_));
  assign new_n21748_ = ~\all_features[1175]  & (~\all_features[1174]  | (~\all_features[1173]  & (new_n21733_ | ~\all_features[1172]  | ~new_n21737_)));
  assign new_n21749_ = ~\all_features[1175]  & ~\all_features[1174]  & ~\all_features[1173]  & ~\all_features[1171]  & ~\all_features[1172] ;
  assign new_n21750_ = new_n21743_ | ~new_n21753_ | ((new_n21734_ | ~new_n21754_) & (new_n21751_ | new_n21746_));
  assign new_n21751_ = new_n21752_ & (~new_n21725_ | ~new_n21738_ | ~new_n21739_);
  assign new_n21752_ = ~new_n21736_ & ~new_n21734_ & ~new_n21747_ & ~new_n21748_;
  assign new_n21753_ = ~new_n21745_ & ~new_n21749_;
  assign new_n21754_ = ~new_n21746_ & ~new_n21736_ & ~new_n21747_ & ~new_n21748_;
  assign new_n21755_ = ~new_n21702_ & ~new_n21715_;
  assign new_n21756_ = ~new_n8927_ & (~new_n8924_ | ~new_n12733_);
  assign new_n21757_ = ~new_n21760_ & ~new_n21759_ & new_n21758_ & (~new_n19883_ | new_n16810_ | ~new_n21755_);
  assign new_n21758_ = (new_n17709_ | ~new_n21714_) & (~new_n21701_ | ~new_n16758_);
  assign new_n21759_ = ~new_n21702_ & ((~new_n19883_ & new_n21756_ & ~new_n21715_) | (~new_n9547_ & ~new_n21716_ & new_n21715_));
  assign new_n21760_ = new_n21722_ & new_n19767_ & new_n21702_ & new_n21704_;
  assign new_n21761_ = ~new_n21762_ & new_n21843_;
  assign new_n21762_ = ~new_n21763_ & ~new_n21839_ & new_n21805_ & (~new_n21840_ | (~new_n21841_ & new_n16026_));
  assign new_n21763_ = ~new_n17676_ & new_n21764_;
  assign new_n21764_ = ~new_n21770_ & new_n21765_;
  assign new_n21765_ = ~new_n21766_ & new_n21767_;
  assign new_n21766_ = ~new_n21563_ & ~new_n19702_;
  assign new_n21767_ = new_n21768_ & new_n21769_;
  assign new_n21768_ = ~new_n8545_ & ~new_n6955_;
  assign new_n21769_ = ~new_n8554_ & ~new_n19233_;
  assign new_n21770_ = ~new_n21771_ & new_n21800_;
  assign new_n21771_ = new_n21772_ & new_n21793_;
  assign new_n21772_ = ~new_n21773_ & (\all_features[2299]  | \all_features[2300]  | \all_features[2301]  | \all_features[2302]  | \all_features[2303] );
  assign new_n21773_ = ~new_n21787_ & (new_n21792_ | (~new_n21789_ & (new_n21790_ | (~new_n21791_ & ~new_n21774_))));
  assign new_n21774_ = ~new_n21775_ & (new_n21777_ | (new_n21786_ & (~new_n21781_ | (~new_n21785_ & new_n21784_))));
  assign new_n21775_ = ~new_n21776_ & ~\all_features[2303] ;
  assign new_n21776_ = \all_features[2301]  & \all_features[2302]  & (\all_features[2300]  | (\all_features[2298]  & \all_features[2299]  & \all_features[2297] ));
  assign new_n21777_ = ~\all_features[2303]  & (~\all_features[2302]  | ~new_n21778_ | ~new_n21779_ | ~new_n21780_);
  assign new_n21778_ = \all_features[2296]  & \all_features[2297] ;
  assign new_n21779_ = \all_features[2300]  & \all_features[2301] ;
  assign new_n21780_ = \all_features[2298]  & \all_features[2299] ;
  assign new_n21781_ = \all_features[2303]  & (\all_features[2302]  | (\all_features[2301]  & (\all_features[2300]  | ~new_n21783_ | ~new_n21782_)));
  assign new_n21782_ = ~\all_features[2296]  & ~\all_features[2297] ;
  assign new_n21783_ = ~\all_features[2298]  & ~\all_features[2299] ;
  assign new_n21784_ = \all_features[2303]  & (\all_features[2302]  | (new_n21779_ & (\all_features[2298]  | \all_features[2299]  | \all_features[2297] )));
  assign new_n21785_ = ~\all_features[2301]  & \all_features[2302]  & \all_features[2303]  & (\all_features[2300]  ? new_n21783_ : (new_n21778_ | ~new_n21783_));
  assign new_n21786_ = \all_features[2303]  & (\all_features[2301]  | \all_features[2302]  | \all_features[2300] );
  assign new_n21787_ = ~\all_features[2301]  & new_n21788_ & ((~\all_features[2298]  & new_n21782_) | ~\all_features[2300]  | ~\all_features[2299] );
  assign new_n21788_ = ~\all_features[2302]  & ~\all_features[2303] ;
  assign new_n21789_ = new_n21788_ & (~\all_features[2299]  | ~new_n21779_ | (~\all_features[2298]  & ~new_n21778_));
  assign new_n21790_ = ~\all_features[2303]  & (~\all_features[2302]  | (~\all_features[2300]  & ~\all_features[2301]  & ~new_n21780_));
  assign new_n21791_ = ~\all_features[2303]  & (~\all_features[2302]  | (~\all_features[2301]  & (new_n21782_ | ~new_n21780_ | ~\all_features[2300] )));
  assign new_n21792_ = new_n21788_ & (~\all_features[2301]  | (~\all_features[2300]  & (~\all_features[2299]  | (~\all_features[2298]  & ~\all_features[2297] ))));
  assign new_n21793_ = new_n21799_ & (~new_n21798_ | (~new_n21794_ & ~new_n21790_ & ~new_n21791_));
  assign new_n21794_ = ~new_n21775_ & ~new_n21777_ & (~new_n21786_ | ~new_n21781_ | new_n21795_);
  assign new_n21795_ = new_n21784_ & new_n21796_ & (new_n21797_ | ~\all_features[2301]  | ~\all_features[2302]  | ~\all_features[2303] );
  assign new_n21796_ = \all_features[2302]  & \all_features[2303]  & (\all_features[2300]  | \all_features[2301]  | new_n21778_ | ~new_n21783_);
  assign new_n21797_ = ~\all_features[2299]  & ~\all_features[2300]  & (~\all_features[2298]  | new_n21782_);
  assign new_n21798_ = ~new_n21789_ & ~new_n21792_;
  assign new_n21799_ = ~new_n21787_ & (\all_features[2299]  | \all_features[2300]  | \all_features[2301]  | \all_features[2302]  | \all_features[2303] );
  assign new_n21800_ = ~new_n21801_ & ~new_n21804_;
  assign new_n21801_ = new_n21802_ & (~new_n21803_ | (new_n21796_ & new_n21786_ & new_n21781_ & new_n21784_));
  assign new_n21802_ = new_n21798_ & new_n21799_;
  assign new_n21803_ = ~new_n21777_ & ~new_n21775_ & ~new_n21790_ & ~new_n21791_;
  assign new_n21804_ = new_n21802_ & new_n21803_;
  assign new_n21805_ = (~new_n20536_ | ~new_n21807_ | ~new_n15672_) & (~new_n21806_ | ~new_n19160_ | ~new_n21808_);
  assign new_n21806_ = new_n21766_ & new_n21767_;
  assign new_n21807_ = ~new_n21767_ & ~new_n14292_;
  assign new_n21808_ = ~new_n21836_ & ~new_n21809_ & ~new_n21834_;
  assign new_n21809_ = new_n21825_ & (~new_n21829_ | (~new_n21810_ & ~new_n21832_ & ~new_n21833_));
  assign new_n21810_ = ~new_n21821_ & ~new_n21823_ & (~new_n21814_ | (~new_n21811_ & new_n21817_ & new_n21819_));
  assign new_n21811_ = \all_features[1415]  & \all_features[1414]  & ~new_n21812_ & \all_features[1413] ;
  assign new_n21812_ = ~\all_features[1411]  & ~\all_features[1412]  & (~\all_features[1410]  | new_n21813_);
  assign new_n21813_ = ~\all_features[1408]  & ~\all_features[1409] ;
  assign new_n21814_ = \all_features[1415]  & (\all_features[1414]  | (~new_n21816_ & new_n21815_));
  assign new_n21815_ = \all_features[1413]  & (\all_features[1410]  | \all_features[1411]  | \all_features[1412]  | ~new_n21813_);
  assign new_n21816_ = ~\all_features[1412]  & ~\all_features[1413] ;
  assign new_n21817_ = \all_features[1415]  & (\all_features[1414]  | (new_n21818_ & (\all_features[1410]  | \all_features[1411]  | \all_features[1409] )));
  assign new_n21818_ = \all_features[1412]  & \all_features[1413] ;
  assign new_n21819_ = \all_features[1414]  & \all_features[1415]  & (\all_features[1410]  | \all_features[1411]  | new_n21820_ | ~new_n21816_);
  assign new_n21820_ = \all_features[1408]  & \all_features[1409] ;
  assign new_n21821_ = ~\all_features[1415]  & (~\all_features[1414]  | ~new_n21820_ | ~new_n21818_ | ~new_n21822_);
  assign new_n21822_ = \all_features[1410]  & \all_features[1411] ;
  assign new_n21823_ = ~new_n21824_ & ~\all_features[1415] ;
  assign new_n21824_ = \all_features[1413]  & \all_features[1414]  & (\all_features[1412]  | (\all_features[1410]  & \all_features[1411]  & \all_features[1409] ));
  assign new_n21825_ = ~new_n21826_ & ~new_n21828_;
  assign new_n21826_ = ~\all_features[1413]  & new_n21827_ & ((~\all_features[1410]  & new_n21813_) | ~\all_features[1412]  | ~\all_features[1411] );
  assign new_n21827_ = ~\all_features[1414]  & ~\all_features[1415] ;
  assign new_n21828_ = ~\all_features[1415]  & ~\all_features[1414]  & ~\all_features[1413]  & ~\all_features[1411]  & ~\all_features[1412] ;
  assign new_n21829_ = ~new_n21830_ & ~new_n21831_;
  assign new_n21830_ = new_n21827_ & (~\all_features[1411]  | ~new_n21818_ | (~\all_features[1410]  & ~new_n21820_));
  assign new_n21831_ = new_n21827_ & (~\all_features[1413]  | (~\all_features[1412]  & (~\all_features[1411]  | (~\all_features[1410]  & ~\all_features[1409] ))));
  assign new_n21832_ = ~\all_features[1415]  & (~\all_features[1414]  | (~\all_features[1413]  & (new_n21813_ | ~new_n21822_ | ~\all_features[1412] )));
  assign new_n21833_ = ~\all_features[1415]  & (~\all_features[1414]  | (~new_n21822_ & new_n21816_));
  assign new_n21834_ = new_n21835_ & ~new_n21833_ & ~new_n21832_ & ~new_n21826_ & ~new_n21830_;
  assign new_n21835_ = ~new_n21828_ & ~new_n21823_ & ~new_n21831_ & ~new_n21821_;
  assign new_n21836_ = new_n21825_ & new_n21829_ & (new_n21837_ | new_n21823_ | new_n21832_ | ~new_n21838_);
  assign new_n21837_ = new_n21819_ & new_n21817_ & \all_features[1415]  & (\all_features[1414]  | (~new_n21816_ & new_n21815_));
  assign new_n21838_ = ~new_n21821_ & ~new_n21833_;
  assign new_n21839_ = new_n21806_ & (new_n21808_ ? ~new_n19160_ : new_n15022_);
  assign new_n21840_ = ~new_n21767_ & new_n14292_;
  assign new_n21841_ = ~new_n11901_ & (~new_n21842_ | new_n6534_);
  assign new_n21842_ = ~new_n6563_ & new_n6566_;
  assign new_n21843_ = new_n21844_ & (~new_n17676_ | ~new_n21764_);
  assign new_n21844_ = ~new_n21846_ & ~new_n21845_ & (~new_n21807_ | (new_n10241_ & ~new_n20536_) | (new_n15672_ & new_n20536_));
  assign new_n21845_ = ~new_n11094_ & new_n21770_ & new_n21765_ & (~new_n11092_ | ~new_n11083_);
  assign new_n21846_ = new_n21840_ & ~new_n21841_ & new_n16026_;
  assign new_n21847_ = ~new_n21914_ & new_n21848_;
  assign new_n21848_ = new_n21849_ & (new_n21854_ | ((~new_n21890_ | new_n21853_) & (new_n17709_ | new_n21892_ | ~new_n21853_)));
  assign new_n21849_ = (new_n14690_ | new_n19835_ | new_n12562_ | ~new_n21854_) & (~new_n21853_ | ~new_n21850_ | new_n21854_);
  assign new_n21850_ = ~new_n21851_ & new_n17709_;
  assign new_n21851_ = new_n21852_ & new_n6388_;
  assign new_n21852_ = new_n6385_ & new_n6378_;
  assign new_n21853_ = ~new_n7475_ & (~new_n7477_ | ~new_n7446_);
  assign new_n21854_ = new_n21855_ & (~new_n21886_ | ~new_n21882_);
  assign new_n21855_ = ~new_n21856_ & ~new_n21880_;
  assign new_n21856_ = new_n21874_ & ~new_n21879_ & ~new_n21857_ & ~new_n21878_;
  assign new_n21857_ = new_n21863_ & (~new_n21858_ | ~new_n21872_ | ~new_n21873_);
  assign new_n21858_ = new_n21859_ & new_n21862_;
  assign new_n21859_ = \all_features[2983]  & (\all_features[2982]  | (\all_features[2981]  & (\all_features[2980]  | ~new_n21861_ | ~new_n21860_)));
  assign new_n21860_ = ~\all_features[2978]  & ~\all_features[2979] ;
  assign new_n21861_ = ~\all_features[2976]  & ~\all_features[2977] ;
  assign new_n21862_ = \all_features[2983]  & (\all_features[2981]  | \all_features[2982]  | \all_features[2980] );
  assign new_n21863_ = ~new_n21871_ & ~new_n21868_ & ~new_n21864_ & ~new_n21866_;
  assign new_n21864_ = ~\all_features[2983]  & (~\all_features[2982]  | (~\all_features[2981]  & (new_n21861_ | ~new_n21865_ | ~\all_features[2980] )));
  assign new_n21865_ = \all_features[2978]  & \all_features[2979] ;
  assign new_n21866_ = ~new_n21867_ & ~\all_features[2983] ;
  assign new_n21867_ = \all_features[2981]  & \all_features[2982]  & (\all_features[2980]  | (\all_features[2978]  & \all_features[2979]  & \all_features[2977] ));
  assign new_n21868_ = ~\all_features[2983]  & (~\all_features[2982]  | ~new_n21869_ | ~new_n21870_ | ~new_n21865_);
  assign new_n21869_ = \all_features[2976]  & \all_features[2977] ;
  assign new_n21870_ = \all_features[2980]  & \all_features[2981] ;
  assign new_n21871_ = ~\all_features[2983]  & (~\all_features[2982]  | (~\all_features[2980]  & ~\all_features[2981]  & ~new_n21865_));
  assign new_n21872_ = \all_features[2982]  & \all_features[2983]  & (\all_features[2980]  | \all_features[2981]  | new_n21869_ | ~new_n21860_);
  assign new_n21873_ = \all_features[2983]  & (\all_features[2982]  | (new_n21870_ & (\all_features[2978]  | \all_features[2979]  | \all_features[2977] )));
  assign new_n21874_ = ~new_n21875_ & ~new_n21877_;
  assign new_n21875_ = ~\all_features[2981]  & new_n21876_ & ((~\all_features[2978]  & new_n21861_) | ~\all_features[2980]  | ~\all_features[2979] );
  assign new_n21876_ = ~\all_features[2982]  & ~\all_features[2983] ;
  assign new_n21877_ = ~\all_features[2983]  & ~\all_features[2982]  & ~\all_features[2981]  & ~\all_features[2979]  & ~\all_features[2980] ;
  assign new_n21878_ = new_n21876_ & (~\all_features[2981]  | (~\all_features[2980]  & (~\all_features[2979]  | (~\all_features[2978]  & ~\all_features[2977] ))));
  assign new_n21879_ = new_n21876_ & (~\all_features[2979]  | ~new_n21870_ | (~\all_features[2978]  & ~new_n21869_));
  assign new_n21880_ = new_n21881_ & new_n21874_ & ~new_n21866_ & ~new_n21878_;
  assign new_n21881_ = ~new_n21879_ & ~new_n21871_ & ~new_n21864_ & ~new_n21868_;
  assign new_n21882_ = new_n21874_ & (new_n21879_ | new_n21878_ | (~new_n21864_ & ~new_n21871_ & ~new_n21883_));
  assign new_n21883_ = ~new_n21866_ & ~new_n21868_ & (~new_n21858_ | (~new_n21884_ & new_n21872_ & new_n21873_));
  assign new_n21884_ = \all_features[2983]  & \all_features[2982]  & ~new_n21885_ & \all_features[2981] ;
  assign new_n21885_ = ~\all_features[2979]  & ~\all_features[2980]  & (~\all_features[2978]  | new_n21861_);
  assign new_n21886_ = ~new_n21877_ & (new_n21875_ | (~new_n21878_ & ~new_n21887_));
  assign new_n21887_ = ~new_n21879_ & (new_n21871_ | (~new_n21864_ & (new_n21866_ | (~new_n21868_ & ~new_n21888_))));
  assign new_n21888_ = new_n21862_ & (~new_n21859_ | (new_n21873_ & (new_n21889_ | ~new_n21872_)));
  assign new_n21889_ = \all_features[2982]  & \all_features[2983]  & (\all_features[2981]  | (~new_n21860_ & \all_features[2980] ));
  assign new_n21890_ = (new_n16744_ | (~new_n19457_ & (~new_n19435_ | ~new_n19463_))) & (new_n21891_ | ~new_n16377_ | new_n19457_ | (new_n19435_ & new_n19463_));
  assign new_n21891_ = new_n16406_ & new_n16402_;
  assign new_n21892_ = ~new_n21893_ & ~new_n21911_ & (new_n21913_ | \all_features[1381]  | \all_features[1382]  | \all_features[1383] );
  assign new_n21893_ = new_n21894_ & (~new_n21909_ | (~new_n21907_ & ~new_n21910_ & ~new_n21904_ & new_n21911_));
  assign new_n21894_ = ~new_n21895_ & ~new_n21898_ & ~new_n21904_ & new_n21906_ & (~new_n21903_ | ~new_n21901_);
  assign new_n21895_ = ~\all_features[1383]  & ~new_n21896_ & ~\all_features[1382] ;
  assign new_n21896_ = \all_features[1379]  & \all_features[1380]  & \all_features[1381]  & (\all_features[1378]  | new_n21897_);
  assign new_n21897_ = \all_features[1376]  & \all_features[1377] ;
  assign new_n21898_ = ~\all_features[1383]  & (~\all_features[1382]  | (~\all_features[1381]  & (new_n21900_ | ~\all_features[1380]  | ~new_n21899_)));
  assign new_n21899_ = \all_features[1378]  & \all_features[1379] ;
  assign new_n21900_ = ~\all_features[1376]  & ~\all_features[1377] ;
  assign new_n21901_ = \all_features[1383]  & (\all_features[1382]  | (\all_features[1381]  & (\all_features[1380]  | ~new_n21902_ | ~new_n21900_)));
  assign new_n21902_ = ~\all_features[1378]  & ~\all_features[1379] ;
  assign new_n21903_ = \all_features[1382]  & \all_features[1383]  & (\all_features[1380]  | \all_features[1381]  | new_n21897_ | ~new_n21902_);
  assign new_n21904_ = ~new_n21905_ & ~\all_features[1383] ;
  assign new_n21905_ = \all_features[1381]  & \all_features[1382]  & (\all_features[1380]  | (\all_features[1378]  & \all_features[1379]  & \all_features[1377] ));
  assign new_n21906_ = \all_features[1383]  | (new_n21897_ & \all_features[1380]  & \all_features[1381]  & \all_features[1382]  & new_n21899_);
  assign new_n21907_ = new_n21901_ & (~new_n21903_ | (~new_n21908_ & \all_features[1381]  & \all_features[1382]  & \all_features[1383] ));
  assign new_n21908_ = ~\all_features[1379]  & ~\all_features[1380]  & (~\all_features[1378]  | new_n21900_);
  assign new_n21909_ = \all_features[1383]  | (\all_features[1382]  & (\all_features[1381]  | (~new_n21900_ & \all_features[1380]  & new_n21899_)));
  assign new_n21910_ = ~\all_features[1383]  & (~new_n21897_ | ~\all_features[1380]  | ~\all_features[1381]  | ~\all_features[1382]  | ~new_n21899_);
  assign new_n21911_ = ~\all_features[1383]  & ~\all_features[1382]  & ~\all_features[1381]  & ~\all_features[1379]  & ~\all_features[1380] ;
  assign new_n21913_ = \all_features[1379]  & \all_features[1380]  & (\all_features[1378]  | ~new_n21900_);
  assign new_n21914_ = new_n21915_ & (new_n21854_ | ((new_n17709_ | ~new_n21892_ | ~new_n21853_) & (new_n21890_ | new_n21853_)));
  assign new_n21915_ = ~new_n21854_ | ((new_n21916_ | ~new_n12562_) & (new_n18594_ | ~new_n19835_ | new_n12562_));
  assign new_n21916_ = ~new_n21944_ & new_n21917_ & (new_n21936_ | ~new_n21918_);
  assign new_n21917_ = ~new_n15819_ & (~new_n16338_ | ~new_n15797_);
  assign new_n21918_ = new_n21936_ & (new_n21940_ | (~new_n21941_ & new_n21919_ & (new_n21928_ | new_n21934_)));
  assign new_n21919_ = ~new_n21928_ & ~new_n21930_ & (~new_n21933_ | ~new_n21932_ | new_n21920_);
  assign new_n21920_ = new_n21921_ & ~new_n21926_ & new_n21923_;
  assign new_n21921_ = \all_features[4287]  & (\all_features[4286]  | (new_n21922_ & (\all_features[4282]  | \all_features[4283]  | \all_features[4281] )));
  assign new_n21922_ = \all_features[4284]  & \all_features[4285] ;
  assign new_n21923_ = new_n21925_ & (\all_features[4284]  | \all_features[4285]  | ~new_n21924_ | (\all_features[4281]  & \all_features[4280] ));
  assign new_n21924_ = ~\all_features[4282]  & ~\all_features[4283] ;
  assign new_n21925_ = \all_features[4286]  & \all_features[4287] ;
  assign new_n21926_ = new_n21925_ & \all_features[4285]  & ((~new_n21927_ & \all_features[4282] ) | \all_features[4284]  | \all_features[4283] );
  assign new_n21927_ = ~\all_features[4280]  & ~\all_features[4281] ;
  assign new_n21928_ = ~new_n21929_ & ~\all_features[4287] ;
  assign new_n21929_ = \all_features[4285]  & \all_features[4286]  & (\all_features[4284]  | (\all_features[4282]  & \all_features[4283]  & \all_features[4281] ));
  assign new_n21930_ = ~\all_features[4287]  & (~new_n21922_ | ~\all_features[4280]  | ~\all_features[4281]  | ~\all_features[4286]  | ~new_n21931_);
  assign new_n21931_ = \all_features[4282]  & \all_features[4283] ;
  assign new_n21932_ = \all_features[4287]  & (\all_features[4286]  | (\all_features[4285]  & (\all_features[4284]  | ~new_n21924_ | ~new_n21927_)));
  assign new_n21933_ = \all_features[4287]  & (\all_features[4285]  | \all_features[4286]  | \all_features[4284] );
  assign new_n21934_ = ~new_n21930_ & (~new_n21933_ | (new_n21932_ & (~new_n21921_ | (~new_n21935_ & new_n21923_))));
  assign new_n21935_ = new_n21925_ & (\all_features[4285]  | (~new_n21924_ & \all_features[4284] ));
  assign new_n21936_ = \all_features[4286]  | \all_features[4287]  | (~new_n21939_ & new_n21937_ & \all_features[4285] );
  assign new_n21937_ = new_n21922_ & \all_features[4283]  & (\all_features[4282]  | (\all_features[4280]  & \all_features[4281] ));
  assign new_n21939_ = ~\all_features[4284]  & (~\all_features[4283]  | (~\all_features[4282]  & ~\all_features[4281] ));
  assign new_n21940_ = ~\all_features[4287]  & (~\all_features[4286]  | (~\all_features[4284]  & ~\all_features[4285]  & ~new_n21931_));
  assign new_n21941_ = ~\all_features[4287]  & (~\all_features[4286]  | (~\all_features[4285]  & (new_n21927_ | ~\all_features[4284]  | ~new_n21931_)));
  assign new_n21944_ = ~\all_features[4287]  & ~\all_features[4286]  & ~\all_features[4285]  & ~\all_features[4283]  & ~\all_features[4284] ;
  assign new_n21945_ = ~new_n21946_ & new_n22043_;
  assign new_n21946_ = new_n21947_ & ((~new_n22041_ & new_n21952_) | (~new_n22040_ & new_n19597_ & new_n16106_ & ~new_n21952_));
  assign new_n21947_ = new_n22038_ & new_n21948_ & (~new_n10247_ | ~new_n22037_);
  assign new_n21948_ = new_n21949_ & (~new_n22035_ | ~new_n14337_ | ~new_n22036_);
  assign new_n21949_ = ~new_n21950_ & (new_n22002_ | ~new_n21997_ | ~new_n21962_);
  assign new_n21950_ = ~new_n8956_ & new_n21961_ & new_n21951_ & (~new_n15869_ | ~new_n8930_ | ~new_n8957_);
  assign new_n21951_ = ~new_n21952_ & ~new_n16106_;
  assign new_n21952_ = new_n14759_ & ~new_n21953_ & ~new_n21957_;
  assign new_n21953_ = ~new_n21954_ & (\all_features[1427]  | \all_features[1428]  | \all_features[1429]  | \all_features[1430]  | \all_features[1431] );
  assign new_n21954_ = ~new_n14763_ & (new_n14766_ | (~new_n14767_ & (new_n14776_ | (~new_n14771_ & ~new_n21955_))));
  assign new_n21955_ = ~new_n14773_ & (new_n14775_ | (new_n14781_ & (~new_n14777_ | (~new_n21956_ & new_n14779_))));
  assign new_n21956_ = ~\all_features[1429]  & \all_features[1430]  & \all_features[1431]  & (\all_features[1428]  ? new_n14778_ : (new_n14769_ | ~new_n14778_));
  assign new_n21957_ = new_n14762_ & (new_n14767_ | new_n14766_ | (~new_n14771_ & ~new_n14776_ & ~new_n21958_));
  assign new_n21958_ = ~new_n14775_ & ~new_n14773_ & (~new_n14781_ | ~new_n14777_ | new_n21959_);
  assign new_n21959_ = new_n14779_ & new_n14780_ & (new_n21960_ | ~\all_features[1429]  | ~\all_features[1430]  | ~\all_features[1431] );
  assign new_n21960_ = ~\all_features[1427]  & ~\all_features[1428]  & (~\all_features[1426]  | new_n14764_);
  assign new_n21961_ = new_n15040_ & new_n6806_;
  assign new_n21962_ = new_n21952_ & new_n21963_;
  assign new_n21963_ = new_n21964_ & (new_n21987_ | (~new_n21994_ & ~new_n21985_));
  assign new_n21964_ = ~new_n21983_ & (~new_n21984_ | (~new_n21965_ & ~new_n21990_ & ~new_n21989_ & new_n21991_));
  assign new_n21965_ = ~new_n21977_ & ~new_n21979_ & (new_n21982_ | new_n21980_ | new_n21966_);
  assign new_n21966_ = new_n21976_ & ~new_n21970_ & new_n21967_;
  assign new_n21967_ = \all_features[4983]  & (\all_features[4982]  | new_n21968_);
  assign new_n21968_ = \all_features[4981]  & (\all_features[4978]  | \all_features[4979]  | \all_features[4980]  | ~new_n21969_);
  assign new_n21969_ = ~\all_features[4976]  & ~\all_features[4977] ;
  assign new_n21970_ = ~new_n21973_ & new_n21971_ & \all_features[4982]  & \all_features[4983]  & (~\all_features[4981]  | new_n21975_);
  assign new_n21971_ = \all_features[4983]  & (\all_features[4982]  | (new_n21972_ & (\all_features[4978]  | \all_features[4979]  | \all_features[4977] )));
  assign new_n21972_ = \all_features[4980]  & \all_features[4981] ;
  assign new_n21973_ = ~\all_features[4981]  & ~\all_features[4980]  & ~\all_features[4979]  & ~new_n21974_ & ~\all_features[4978] ;
  assign new_n21974_ = \all_features[4976]  & \all_features[4977] ;
  assign new_n21975_ = ~\all_features[4979]  & ~\all_features[4980]  & (~\all_features[4978]  | new_n21969_);
  assign new_n21976_ = \all_features[4983]  & (\all_features[4981]  | \all_features[4982]  | \all_features[4980] );
  assign new_n21977_ = ~\all_features[4983]  & (~\all_features[4982]  | (~\all_features[4980]  & ~\all_features[4981]  & ~new_n21978_));
  assign new_n21978_ = \all_features[4978]  & \all_features[4979] ;
  assign new_n21979_ = ~\all_features[4983]  & (~\all_features[4982]  | (~\all_features[4981]  & (new_n21969_ | ~new_n21978_ | ~\all_features[4980] )));
  assign new_n21980_ = ~new_n21981_ & ~\all_features[4983] ;
  assign new_n21981_ = \all_features[4981]  & \all_features[4982]  & (\all_features[4980]  | (\all_features[4978]  & \all_features[4979]  & \all_features[4977] ));
  assign new_n21982_ = ~\all_features[4983]  & (~\all_features[4982]  | ~new_n21974_ | ~new_n21972_ | ~new_n21978_);
  assign new_n21983_ = new_n21988_ & new_n21984_ & ~new_n21990_ & ~new_n21980_;
  assign new_n21984_ = ~new_n21985_ & ~new_n21987_;
  assign new_n21985_ = ~\all_features[4981]  & new_n21986_ & ((~\all_features[4978]  & new_n21969_) | ~\all_features[4980]  | ~\all_features[4979] );
  assign new_n21986_ = ~\all_features[4982]  & ~\all_features[4983] ;
  assign new_n21987_ = ~\all_features[4983]  & ~\all_features[4982]  & ~\all_features[4981]  & ~\all_features[4979]  & ~\all_features[4980] ;
  assign new_n21988_ = ~new_n21982_ & ~new_n21979_ & ~new_n21989_ & ~new_n21977_;
  assign new_n21989_ = new_n21986_ & (~\all_features[4979]  | ~new_n21972_ | (~\all_features[4978]  & ~new_n21974_));
  assign new_n21990_ = new_n21986_ & (~\all_features[4981]  | (~\all_features[4980]  & (~\all_features[4979]  | (~\all_features[4978]  & ~\all_features[4977] ))));
  assign new_n21991_ = new_n21993_ & (~new_n21971_ | ~new_n21976_ | ~new_n21992_ | ~new_n21967_);
  assign new_n21992_ = \all_features[4983]  & ~new_n21973_ & \all_features[4982] ;
  assign new_n21993_ = ~new_n21982_ & ~new_n21980_ & ~new_n21977_ & ~new_n21979_;
  assign new_n21994_ = ~new_n21990_ & (new_n21989_ | (~new_n21977_ & (new_n21979_ | (~new_n21995_ & ~new_n21980_))));
  assign new_n21995_ = ~new_n21982_ & (~new_n21976_ | (new_n21967_ & (~new_n21971_ | (~new_n21996_ & new_n21992_))));
  assign new_n21996_ = \all_features[4982]  & \all_features[4983]  & (\all_features[4981]  | (\all_features[4980]  & (\all_features[4979]  | \all_features[4978] )));
  assign new_n21997_ = ~new_n21998_ & new_n16336_;
  assign new_n21998_ = ~new_n21999_ & (\all_features[987]  | \all_features[988]  | \all_features[989]  | \all_features[990]  | \all_features[991] );
  assign new_n21999_ = ~new_n15815_ & (new_n15817_ | (~new_n15818_ & (new_n15805_ | (~new_n15800_ & ~new_n22000_))));
  assign new_n22000_ = ~new_n15803_ & (new_n15806_ | (new_n15813_ & (~new_n15809_ | (~new_n22001_ & new_n15811_))));
  assign new_n22001_ = ~\all_features[989]  & \all_features[990]  & \all_features[991]  & (\all_features[988]  ? new_n15810_ : (new_n15808_ | ~new_n15810_));
  assign new_n22002_ = ~new_n22003_ & new_n22030_;
  assign new_n22003_ = ~new_n22029_ & (~new_n22022_ | (~new_n22027_ & (new_n22020_ | new_n22028_ | ~new_n22004_)));
  assign new_n22004_ = ~new_n22016_ & ~new_n22014_ & ((~new_n22011_ & new_n22005_) | ~new_n22019_ | ~new_n22018_);
  assign new_n22005_ = \all_features[4063]  & \all_features[4062]  & ~new_n22008_ & new_n22006_;
  assign new_n22006_ = \all_features[4063]  & (\all_features[4062]  | (new_n22007_ & (\all_features[4058]  | \all_features[4059]  | \all_features[4057] )));
  assign new_n22007_ = \all_features[4060]  & \all_features[4061] ;
  assign new_n22008_ = new_n22010_ & ~\all_features[4061]  & ~new_n22009_ & ~\all_features[4060] ;
  assign new_n22009_ = \all_features[4056]  & \all_features[4057] ;
  assign new_n22010_ = ~\all_features[4058]  & ~\all_features[4059] ;
  assign new_n22011_ = \all_features[4063]  & \all_features[4062]  & ~new_n22012_ & \all_features[4061] ;
  assign new_n22012_ = ~\all_features[4059]  & ~\all_features[4060]  & (~\all_features[4058]  | new_n22013_);
  assign new_n22013_ = ~\all_features[4056]  & ~\all_features[4057] ;
  assign new_n22014_ = ~new_n22015_ & ~\all_features[4063] ;
  assign new_n22015_ = \all_features[4061]  & \all_features[4062]  & (\all_features[4060]  | (\all_features[4058]  & \all_features[4059]  & \all_features[4057] ));
  assign new_n22016_ = ~\all_features[4063]  & (~\all_features[4062]  | ~new_n22017_ | ~new_n22009_ | ~new_n22007_);
  assign new_n22017_ = \all_features[4058]  & \all_features[4059] ;
  assign new_n22018_ = \all_features[4063]  & (\all_features[4062]  | (\all_features[4061]  & (\all_features[4060]  | ~new_n22010_ | ~new_n22013_)));
  assign new_n22019_ = \all_features[4063]  & (\all_features[4061]  | \all_features[4062]  | \all_features[4060] );
  assign new_n22020_ = ~new_n22014_ & (new_n22016_ | (new_n22019_ & (~new_n22018_ | (~new_n22021_ & new_n22006_))));
  assign new_n22021_ = ~\all_features[4061]  & \all_features[4062]  & \all_features[4063]  & (\all_features[4060]  ? new_n22010_ : (new_n22009_ | ~new_n22010_));
  assign new_n22022_ = ~new_n22026_ & ~new_n22023_ & ~new_n22025_;
  assign new_n22023_ = new_n22024_ & (~\all_features[4061]  | (~\all_features[4060]  & (~\all_features[4059]  | (~\all_features[4058]  & ~\all_features[4057] ))));
  assign new_n22024_ = ~\all_features[4062]  & ~\all_features[4063] ;
  assign new_n22025_ = ~\all_features[4061]  & new_n22024_ & ((~\all_features[4058]  & new_n22013_) | ~\all_features[4060]  | ~\all_features[4059] );
  assign new_n22026_ = new_n22024_ & (~\all_features[4059]  | ~new_n22007_ | (~\all_features[4058]  & ~new_n22009_));
  assign new_n22027_ = ~\all_features[4063]  & (~\all_features[4062]  | (~\all_features[4060]  & ~\all_features[4061]  & ~new_n22017_));
  assign new_n22028_ = ~\all_features[4063]  & (~\all_features[4062]  | (~\all_features[4061]  & (new_n22013_ | ~\all_features[4060]  | ~new_n22017_)));
  assign new_n22029_ = ~\all_features[4063]  & ~\all_features[4062]  & ~\all_features[4061]  & ~\all_features[4059]  & ~\all_features[4060] ;
  assign new_n22030_ = new_n22023_ | ~new_n22033_ | ((new_n22014_ | ~new_n22034_) & (new_n22031_ | new_n22026_));
  assign new_n22031_ = new_n22032_ & (~new_n22005_ | ~new_n22018_ | ~new_n22019_);
  assign new_n22032_ = ~new_n22016_ & ~new_n22014_ & ~new_n22027_ & ~new_n22028_;
  assign new_n22033_ = ~new_n22025_ & ~new_n22029_;
  assign new_n22034_ = ~new_n22026_ & ~new_n22016_ & ~new_n22027_ & ~new_n22028_;
  assign new_n22035_ = ~new_n21963_ & new_n21952_;
  assign new_n22036_ = ~new_n10099_ & ~new_n10072_ & ~new_n10097_;
  assign new_n22037_ = ~new_n21961_ & new_n21951_;
  assign new_n22038_ = ~new_n22039_ | (new_n19597_ ? ~new_n22040_ : ~new_n14159_);
  assign new_n22039_ = ~new_n21952_ & new_n16106_;
  assign new_n22040_ = new_n17699_ & (new_n17705_ | new_n17677_);
  assign new_n22041_ = (new_n21997_ | new_n14317_ | ~new_n21963_) & (new_n14337_ | ~new_n22042_ | new_n21963_);
  assign new_n22042_ = ~new_n6734_ & new_n8478_;
  assign new_n22043_ = new_n22044_ & (new_n10247_ | ~new_n22037_) & (new_n19597_ | new_n14159_ | ~new_n22039_);
  assign new_n22044_ = ~new_n22045_ & (~new_n21962_ | (~new_n22002_ & new_n21997_) | (~new_n14317_ & ~new_n21997_));
  assign new_n22045_ = new_n22035_ & (new_n14337_ ? ~new_n22036_ : ~new_n22042_);
  assign new_n22046_ = (new_n22047_ & ~new_n18221_ & (~new_n18194_ | ~new_n18217_)) | (~new_n13560_ & ~new_n8765_ & (new_n18221_ | (new_n18194_ & new_n18217_)));
  assign new_n22047_ = (new_n22049_ | new_n22050_ | (new_n22083_ & new_n22052_)) & (new_n22051_ | new_n22048_ | ~new_n22050_);
  assign new_n22048_ = new_n10876_ & new_n20881_;
  assign new_n22049_ = ~new_n15860_ & (~new_n15862_ | ~new_n16105_);
  assign new_n22050_ = ~new_n20405_ & new_n20376_;
  assign new_n22051_ = ~new_n14045_ & new_n12977_;
  assign new_n22052_ = new_n22053_ & new_n22080_;
  assign new_n22053_ = new_n22065_ & (~new_n22069_ | (new_n22072_ & (~new_n22076_ | new_n22054_)));
  assign new_n22054_ = new_n22055_ & (~new_n22059_ | (~new_n22064_ & \all_features[5229]  & \all_features[5230]  & \all_features[5231] ));
  assign new_n22055_ = \all_features[5231]  & (\all_features[5230]  | (~new_n22056_ & \all_features[5229] ));
  assign new_n22056_ = new_n22057_ & ~\all_features[5228]  & new_n22058_;
  assign new_n22057_ = ~\all_features[5224]  & ~\all_features[5225] ;
  assign new_n22058_ = ~\all_features[5226]  & ~\all_features[5227] ;
  assign new_n22059_ = \all_features[5231]  & \all_features[5230]  & ~new_n22062_ & new_n22060_;
  assign new_n22060_ = \all_features[5231]  & (\all_features[5230]  | (new_n22061_ & (\all_features[5226]  | \all_features[5227]  | \all_features[5225] )));
  assign new_n22061_ = \all_features[5228]  & \all_features[5229] ;
  assign new_n22062_ = new_n22058_ & ~\all_features[5229]  & ~new_n22063_ & ~\all_features[5228] ;
  assign new_n22063_ = \all_features[5224]  & \all_features[5225] ;
  assign new_n22064_ = ~\all_features[5227]  & ~\all_features[5228]  & (~\all_features[5226]  | new_n22057_);
  assign new_n22065_ = ~new_n22066_ & ~new_n22068_;
  assign new_n22066_ = ~\all_features[5229]  & new_n22067_ & ((~\all_features[5226]  & new_n22057_) | ~\all_features[5228]  | ~\all_features[5227] );
  assign new_n22067_ = ~\all_features[5230]  & ~\all_features[5231] ;
  assign new_n22068_ = ~\all_features[5231]  & ~\all_features[5230]  & ~\all_features[5229]  & ~\all_features[5227]  & ~\all_features[5228] ;
  assign new_n22069_ = ~new_n22070_ & ~new_n22071_;
  assign new_n22070_ = new_n22067_ & (~\all_features[5227]  | ~new_n22061_ | (~\all_features[5226]  & ~new_n22063_));
  assign new_n22071_ = new_n22067_ & (~\all_features[5229]  | (~\all_features[5228]  & (~\all_features[5227]  | (~\all_features[5226]  & ~\all_features[5225] ))));
  assign new_n22072_ = ~new_n22073_ & ~new_n22075_;
  assign new_n22073_ = ~\all_features[5231]  & (~\all_features[5230]  | (~\all_features[5228]  & ~\all_features[5229]  & ~new_n22074_));
  assign new_n22074_ = \all_features[5226]  & \all_features[5227] ;
  assign new_n22075_ = ~\all_features[5231]  & (~\all_features[5230]  | (~\all_features[5229]  & (new_n22057_ | ~new_n22074_ | ~\all_features[5228] )));
  assign new_n22076_ = ~new_n22077_ & ~new_n22078_;
  assign new_n22077_ = ~\all_features[5231]  & (~\all_features[5230]  | ~new_n22063_ | ~new_n22061_ | ~new_n22074_);
  assign new_n22078_ = ~new_n22079_ & ~\all_features[5231] ;
  assign new_n22079_ = \all_features[5229]  & \all_features[5230]  & (\all_features[5228]  | (\all_features[5226]  & \all_features[5227]  & \all_features[5225] ));
  assign new_n22080_ = new_n22081_ & (new_n22075_ | new_n22078_ | ~new_n22082_ | (new_n22059_ & new_n22055_));
  assign new_n22081_ = new_n22065_ & new_n22069_;
  assign new_n22082_ = ~new_n22073_ & ~new_n22077_;
  assign new_n22083_ = new_n22076_ & new_n22081_ & new_n22072_;
  assign \o[22]  = ~new_n22085_ ^ new_n22086_;
  assign new_n22085_ = (new_n21945_ & new_n22046_) | (~new_n20027_ & (new_n21945_ | new_n22046_));
  assign new_n22086_ = new_n22087_ ? (~new_n22088_ ^ new_n22188_) : (new_n22088_ ^ new_n22188_);
  assign new_n22087_ = (new_n21761_ & new_n21847_) | (~new_n20028_ & (new_n21761_ | new_n21847_));
  assign new_n22088_ = new_n22089_ ? (~new_n22090_ ^ new_n22187_) : (new_n22090_ ^ new_n22187_);
  assign new_n22089_ = (~new_n21393_ & new_n21698_) | (~new_n20029_ & (~new_n21393_ | new_n21698_));
  assign new_n22090_ = new_n22091_ ? (new_n22092_ ^ new_n22133_) : (~new_n22092_ ^ new_n22133_);
  assign new_n22091_ = (~new_n20873_ & new_n21392_) | (~new_n20030_ & (~new_n20873_ | new_n21392_));
  assign new_n22092_ = new_n22093_ ? (new_n22110_ ^ new_n22111_) : (~new_n22110_ ^ new_n22111_);
  assign new_n22093_ = new_n22094_ ? (~new_n22108_ ^ new_n22109_) : (new_n22108_ ^ new_n22109_);
  assign new_n22094_ = new_n22095_ ? (new_n22099_ ^ new_n22107_) : (~new_n22099_ ^ new_n22107_);
  assign new_n22095_ = new_n22096_ ? (new_n22097_ ^ new_n22098_) : (~new_n22097_ ^ new_n22098_);
  assign new_n22096_ = new_n20034_ & new_n20089_;
  assign new_n22097_ = new_n21053_ & new_n21182_;
  assign new_n22098_ = new_n21566_ & new_n21597_;
  assign new_n22099_ = new_n22100_ ? (new_n22101_ ^ new_n22102_) : (~new_n22101_ ^ new_n22102_);
  assign new_n22100_ = new_n21620_ & new_n21681_;
  assign new_n22101_ = ~new_n20147_ & new_n20093_;
  assign new_n22102_ = new_n22103_ & ~new_n21696_ & new_n21687_;
  assign new_n22103_ = ~new_n22106_ & ~new_n22104_ & (~new_n21691_ | (new_n12190_ & new_n21695_) | (~new_n21692_ & ~new_n21695_));
  assign new_n22104_ = ~new_n21689_ & ~new_n22105_ & ~new_n15592_;
  assign new_n22105_ = new_n12228_ ? (new_n8854_ | (~new_n8819_ & new_n8851_)) : ~new_n8225_;
  assign new_n22106_ = new_n15592_ & ~new_n21690_ & ~new_n16758_ & ~new_n21689_;
  assign new_n22107_ = (new_n20961_ & new_n21052_) | (new_n20876_ & (new_n20961_ | new_n21052_));
  assign new_n22108_ = (new_n20236_ & new_n20269_) | (~new_n20032_ & (new_n20236_ | new_n20269_));
  assign new_n22109_ = (~new_n21184_ & new_n21347_) | (new_n20875_ & (~new_n21184_ | new_n21347_));
  assign new_n22110_ = (~new_n20451_ & new_n20805_) | (~new_n20031_ & (~new_n20451_ | new_n20805_));
  assign new_n22111_ = new_n22112_ ? (new_n22119_ ^ new_n22132_) : (~new_n22119_ ^ new_n22132_);
  assign new_n22112_ = new_n22113_ ? (~new_n22114_ ^ new_n22115_) : (new_n22114_ ^ new_n22115_);
  assign new_n22113_ = (new_n20092_ & new_n20148_) | (new_n20033_ & (new_n20092_ | new_n20148_));
  assign new_n22114_ = (new_n20490_ & new_n20574_) | (new_n20453_ & (new_n20490_ | new_n20574_));
  assign new_n22115_ = new_n22116_ ? (new_n22117_ ^ new_n22118_) : (~new_n22117_ ^ new_n22118_);
  assign new_n22116_ = new_n21699_ & new_n21757_;
  assign new_n22117_ = new_n20455_ & new_n20487_;
  assign new_n22118_ = new_n20575_ & new_n20625_;
  assign new_n22119_ = new_n22120_ ? (~new_n22127_ ^ new_n22131_) : (new_n22127_ ^ new_n22131_);
  assign new_n22120_ = new_n22121_ ? (new_n22122_ ^ new_n22124_) : (~new_n22122_ ^ new_n22124_);
  assign new_n22121_ = new_n21947_ & new_n22043_;
  assign new_n22122_ = new_n20629_ & ~new_n22123_ & new_n20772_;
  assign new_n22123_ = (~new_n20729_ | ~new_n20728_) & (~new_n20774_ | (new_n20777_ ? ~new_n6532_ : ~new_n20775_));
  assign new_n22124_ = ~new_n22125_ & new_n22126_;
  assign new_n22125_ = ~new_n20795_ & new_n20802_;
  assign new_n22126_ = ~new_n20796_ & new_n20780_;
  assign new_n22127_ = new_n22128_ ? (new_n22129_ ^ new_n22130_) : (~new_n22129_ ^ new_n22130_);
  assign new_n22128_ = new_n21762_ & new_n21843_;
  assign new_n22129_ = new_n21848_ & new_n21914_;
  assign new_n22130_ = new_n20491_ & new_n20571_;
  assign new_n22131_ = ~new_n20628_ & ~new_n20779_;
  assign new_n22132_ = (~new_n20627_ & new_n20236_) | (~new_n20452_ & (~new_n20627_ | new_n20236_));
  assign new_n22133_ = new_n22134_ ? (~new_n22185_ ^ new_n22186_) : (new_n22185_ ^ new_n22186_);
  assign new_n22134_ = new_n22135_ ? (~new_n22183_ ^ new_n22184_) : (new_n22183_ ^ new_n22184_);
  assign new_n22135_ = new_n22136_ ? (~new_n22181_ ^ new_n22182_) : (new_n22181_ ^ new_n22182_);
  assign new_n22136_ = new_n22137_ ? (new_n22141_ ^ new_n22180_) : (~new_n22141_ ^ new_n22180_);
  assign new_n22137_ = ~new_n22140_ & new_n20876_ & new_n22138_ & (~new_n20887_ | ~new_n20878_);
  assign new_n22138_ = new_n22139_ & (new_n20960_ | ~new_n20892_) & (~new_n20958_ | ~new_n20890_);
  assign new_n22139_ = (~new_n20894_ | ~new_n20893_) & (~new_n20885_ | (new_n11614_ ? ~new_n14618_ : ~new_n20888_));
  assign new_n22140_ = ~new_n19340_ & new_n20891_ & (new_n16222_ | (new_n19158_ & new_n16216_));
  assign new_n22141_ = ~new_n22142_ & ~new_n22144_ & new_n21348_ & (~new_n22143_ | (~new_n21349_ & ~new_n21351_));
  assign new_n22142_ = new_n21355_ & ~new_n21353_ & ~new_n21389_;
  assign new_n22143_ = new_n21355_ & new_n21389_;
  assign new_n22144_ = ~new_n21355_ & ~new_n21390_ & (~new_n22175_ | new_n22145_);
  assign new_n22145_ = new_n22146_ & new_n22167_;
  assign new_n22146_ = ~new_n22147_ & (\all_features[5475]  | \all_features[5476]  | \all_features[5477]  | \all_features[5478]  | \all_features[5479] );
  assign new_n22147_ = ~new_n22161_ & (new_n22166_ | (~new_n22163_ & (new_n22164_ | (~new_n22165_ & ~new_n22148_))));
  assign new_n22148_ = ~new_n22149_ & (new_n22158_ | (new_n22160_ & (~new_n22151_ | (~new_n22156_ & new_n22154_))));
  assign new_n22149_ = ~new_n22150_ & ~\all_features[5479] ;
  assign new_n22150_ = \all_features[5477]  & \all_features[5478]  & (\all_features[5476]  | (\all_features[5474]  & \all_features[5475]  & \all_features[5473] ));
  assign new_n22151_ = \all_features[5479]  & (\all_features[5478]  | (\all_features[5477]  & (\all_features[5476]  | ~new_n22153_ | ~new_n22152_)));
  assign new_n22152_ = ~\all_features[5472]  & ~\all_features[5473] ;
  assign new_n22153_ = ~\all_features[5474]  & ~\all_features[5475] ;
  assign new_n22154_ = \all_features[5479]  & (\all_features[5478]  | (new_n22155_ & (\all_features[5474]  | \all_features[5475]  | \all_features[5473] )));
  assign new_n22155_ = \all_features[5476]  & \all_features[5477] ;
  assign new_n22156_ = ~\all_features[5477]  & \all_features[5478]  & \all_features[5479]  & (\all_features[5476]  ? new_n22153_ : (new_n22157_ | ~new_n22153_));
  assign new_n22157_ = \all_features[5472]  & \all_features[5473] ;
  assign new_n22158_ = ~\all_features[5479]  & (~\all_features[5478]  | ~new_n22157_ | ~new_n22155_ | ~new_n22159_);
  assign new_n22159_ = \all_features[5474]  & \all_features[5475] ;
  assign new_n22160_ = \all_features[5479]  & (\all_features[5477]  | \all_features[5478]  | \all_features[5476] );
  assign new_n22161_ = ~\all_features[5477]  & new_n22162_ & ((~\all_features[5474]  & new_n22152_) | ~\all_features[5476]  | ~\all_features[5475] );
  assign new_n22162_ = ~\all_features[5478]  & ~\all_features[5479] ;
  assign new_n22163_ = new_n22162_ & (~\all_features[5475]  | ~new_n22155_ | (~\all_features[5474]  & ~new_n22157_));
  assign new_n22164_ = ~\all_features[5479]  & (~\all_features[5478]  | (~\all_features[5476]  & ~\all_features[5477]  & ~new_n22159_));
  assign new_n22165_ = ~\all_features[5479]  & (~\all_features[5478]  | (~\all_features[5477]  & (new_n22152_ | ~new_n22159_ | ~\all_features[5476] )));
  assign new_n22166_ = new_n22162_ & (~\all_features[5477]  | (~\all_features[5476]  & (~\all_features[5475]  | (~\all_features[5474]  & ~\all_features[5473] ))));
  assign new_n22167_ = new_n22173_ & (~new_n22174_ | (~new_n22168_ & ~new_n22164_ & ~new_n22165_));
  assign new_n22168_ = new_n22171_ & ((~new_n22169_ & new_n22154_ & new_n22172_) | ~new_n22160_ | ~new_n22151_);
  assign new_n22169_ = \all_features[5479]  & \all_features[5478]  & ~new_n22170_ & \all_features[5477] ;
  assign new_n22170_ = ~\all_features[5475]  & ~\all_features[5476]  & (~\all_features[5474]  | new_n22152_);
  assign new_n22171_ = ~new_n22149_ & ~new_n22158_;
  assign new_n22172_ = \all_features[5478]  & \all_features[5479]  & (\all_features[5476]  | \all_features[5477]  | new_n22157_ | ~new_n22153_);
  assign new_n22173_ = ~new_n22161_ & (\all_features[5475]  | \all_features[5476]  | \all_features[5477]  | \all_features[5478]  | \all_features[5479] );
  assign new_n22174_ = ~new_n22163_ & ~new_n22166_;
  assign new_n22175_ = ~new_n22176_ & ~new_n22179_;
  assign new_n22176_ = new_n22174_ & ~new_n22177_ & new_n22173_;
  assign new_n22177_ = new_n22178_ & (~new_n22172_ | ~new_n22160_ | ~new_n22151_ | ~new_n22154_);
  assign new_n22178_ = ~new_n22158_ & ~new_n22149_ & ~new_n22164_ & ~new_n22165_;
  assign new_n22179_ = new_n22171_ & new_n22173_ & ~new_n22166_ & ~new_n22165_ & ~new_n22163_ & ~new_n22164_;
  assign new_n22180_ = new_n21186_ & new_n21246_;
  assign new_n22181_ = (new_n21488_ & new_n21532_) | (new_n21447_ & (new_n21488_ | new_n21532_));
  assign new_n22182_ = (~new_n21247_ & new_n21185_) | (new_n20237_ & (~new_n21247_ | new_n21185_));
  assign new_n22183_ = (~new_n21446_ & new_n21347_) | (new_n21396_ & (~new_n21446_ | new_n21347_));
  assign new_n22184_ = new_n21397_ & new_n21442_;
  assign new_n22185_ = (new_n20805_ & new_n21348_) | (~new_n20874_ & (new_n20805_ | new_n21348_));
  assign new_n22186_ = (new_n21565_ & new_n21600_) | (~new_n21395_ & (new_n21565_ | new_n21600_));
  assign new_n22187_ = (new_n21619_ & new_n21686_) | (~new_n21394_ & (new_n21619_ | new_n21686_));
  assign new_n22188_ = ~new_n21531_ & new_n21489_;
  assign \o[23]  = ~new_n22190_ ^ new_n22191_;
  assign new_n22190_ = ~new_n22086_ & new_n22085_;
  assign new_n22191_ = new_n22192_ ^ new_n22193_;
  assign new_n22192_ = (~new_n22088_ & new_n22188_) | (new_n22087_ & (~new_n22088_ | new_n22188_));
  assign new_n22193_ = ~new_n22194_ ^ new_n22195_;
  assign new_n22194_ = (~new_n22090_ & new_n22187_) | (new_n22089_ & (~new_n22090_ | new_n22187_));
  assign new_n22195_ = new_n22196_ ? (new_n22197_ ^ new_n22223_) : (~new_n22197_ ^ new_n22223_);
  assign new_n22196_ = (~new_n22092_ & ~new_n22133_) | (new_n22091_ & (~new_n22092_ | ~new_n22133_));
  assign new_n22197_ = new_n22198_ ? (new_n22206_ ^ new_n22207_) : (~new_n22206_ ^ new_n22207_);
  assign new_n22198_ = new_n22199_ ? (~new_n22204_ ^ new_n22205_) : (new_n22204_ ^ new_n22205_);
  assign new_n22199_ = ~new_n22200_ ^ new_n22203_;
  assign new_n22200_ = new_n22201_ ^ new_n22202_;
  assign new_n22201_ = (new_n22097_ & new_n22098_) | (new_n22096_ & (new_n22097_ | new_n22098_));
  assign new_n22202_ = (new_n22141_ & new_n22180_) | (new_n22137_ & (new_n22141_ | new_n22180_));
  assign new_n22203_ = (new_n22181_ & new_n22182_) | (~new_n22136_ & (new_n22181_ | new_n22182_));
  assign new_n22204_ = (new_n22108_ & new_n22109_) | (~new_n22094_ & (new_n22108_ | new_n22109_));
  assign new_n22205_ = (new_n22183_ & new_n22184_) | (~new_n22135_ & (new_n22183_ | new_n22184_));
  assign new_n22206_ = (~new_n22111_ & new_n22110_) | (~new_n22093_ & (~new_n22111_ | new_n22110_));
  assign new_n22207_ = new_n22208_ ? (new_n22212_ ^ new_n22213_) : (~new_n22212_ ^ new_n22213_);
  assign new_n22208_ = new_n22209_ ? (new_n22210_ ^ new_n22211_) : (~new_n22210_ ^ new_n22211_);
  assign new_n22209_ = (~new_n22099_ & new_n22107_) | (~new_n22095_ & (~new_n22099_ | new_n22107_));
  assign new_n22210_ = (~new_n22115_ & new_n22114_) | (new_n22113_ & (~new_n22115_ | new_n22114_));
  assign new_n22211_ = (new_n22101_ & new_n22102_) | (new_n22100_ & (new_n22101_ | new_n22102_));
  assign new_n22212_ = (~new_n22119_ & new_n22132_) | (~new_n22112_ & (~new_n22119_ | new_n22132_));
  assign new_n22213_ = new_n22214_ ? (new_n22217_ ^ new_n22218_) : (~new_n22217_ ^ new_n22218_);
  assign new_n22214_ = ~new_n22215_ ^ new_n22216_;
  assign new_n22215_ = (new_n22129_ & new_n22130_) | (new_n22128_ & (new_n22129_ | new_n22130_));
  assign new_n22216_ = (new_n22117_ & new_n22118_) | (new_n22116_ & (new_n22117_ | new_n22118_));
  assign new_n22217_ = (~new_n22127_ & ~new_n22131_) | (~new_n22120_ & (~new_n22127_ | ~new_n22131_));
  assign new_n22218_ = new_n22219_ ^ new_n22220_;
  assign new_n22219_ = (new_n22122_ & new_n22124_) | (new_n22121_ & (new_n22122_ | new_n22124_));
  assign new_n22220_ = new_n22221_ ^ new_n22222_;
  assign new_n22221_ = new_n22123_ & new_n20629_ & new_n20772_;
  assign new_n22222_ = new_n22125_ & new_n22126_;
  assign new_n22223_ = (new_n22185_ & new_n22186_) | (~new_n22134_ & (new_n22185_ | new_n22186_));
  assign \o[24]  = ((new_n22225_ | new_n22226_) & (new_n22227_ ^ new_n22228_)) | (~new_n22225_ & ~new_n22226_ & (~new_n22227_ ^ new_n22228_));
  assign new_n22225_ = ~new_n22191_ & new_n22190_;
  assign new_n22226_ = ~new_n22193_ & new_n22192_;
  assign new_n22227_ = new_n22194_ & new_n22195_;
  assign new_n22228_ = ~new_n22229_ ^ new_n22230_;
  assign new_n22229_ = (~new_n22197_ & new_n22223_) | (new_n22196_ & (~new_n22197_ | new_n22223_));
  assign new_n22230_ = new_n22231_ ? (new_n22232_ ^ new_n22244_) : (~new_n22232_ ^ new_n22244_);
  assign new_n22231_ = (~new_n22207_ & new_n22206_) | (~new_n22198_ & (~new_n22207_ | new_n22206_));
  assign new_n22232_ = new_n22233_ ? (new_n22237_ ^ new_n22238_) : (~new_n22237_ ^ new_n22238_);
  assign new_n22233_ = new_n22234_ ? (new_n22235_ ^ new_n22236_) : (~new_n22235_ ^ new_n22236_);
  assign new_n22234_ = new_n22200_ & new_n22203_;
  assign new_n22235_ = (new_n22210_ & new_n22211_) | (new_n22209_ & (new_n22210_ | new_n22211_));
  assign new_n22236_ = new_n22201_ & new_n22202_;
  assign new_n22237_ = (~new_n22213_ & new_n22212_) | (~new_n22208_ & (~new_n22213_ | new_n22212_));
  assign new_n22238_ = new_n22239_ ? (~new_n22240_ ^ new_n22243_) : (new_n22240_ ^ new_n22243_);
  assign new_n22239_ = (~new_n22218_ & new_n22217_) | (~new_n22214_ & (~new_n22218_ | new_n22217_));
  assign new_n22240_ = new_n22241_ ^ new_n22242_;
  assign new_n22241_ = ~new_n22220_ & new_n22219_;
  assign new_n22242_ = ~new_n22221_ & ~new_n22222_;
  assign new_n22243_ = new_n22215_ & new_n22216_;
  assign new_n22244_ = (new_n22204_ & new_n22205_) | (~new_n22199_ & (new_n22204_ | new_n22205_));
  assign \o[25]  = ~new_n22246_ ^ new_n22247_;
  assign new_n22246_ = (new_n22227_ | (~new_n22228_ & (new_n22226_ | new_n22225_))) & (new_n22226_ | new_n22225_ | ~new_n22228_);
  assign new_n22247_ = new_n22248_ ^ new_n22249_;
  assign new_n22248_ = new_n22229_ & new_n22230_;
  assign new_n22249_ = ~new_n22250_ ^ new_n22251_;
  assign new_n22250_ = (~new_n22232_ & new_n22244_) | (new_n22231_ & (~new_n22232_ | new_n22244_));
  assign new_n22251_ = new_n22252_ ? (new_n22253_ ^ new_n22254_) : (~new_n22253_ ^ new_n22254_);
  assign new_n22252_ = (~new_n22238_ & new_n22237_) | (~new_n22233_ & (~new_n22238_ | new_n22237_));
  assign new_n22253_ = (new_n22235_ & new_n22236_) | (new_n22234_ & (new_n22235_ | new_n22236_));
  assign new_n22254_ = ~new_n22255_ ^ new_n22256_;
  assign new_n22255_ = (~new_n22240_ & new_n22243_) | (new_n22239_ & (~new_n22240_ | new_n22243_));
  assign new_n22256_ = ~new_n22242_ & new_n22241_;
  assign \o[26]  = ((new_n22261_ ^ new_n22262_) & ((~new_n22258_ & ~new_n22259_ & ~new_n22260_) | (new_n22260_ & (new_n22258_ | new_n22259_)))) | (((~new_n22260_ & (new_n22258_ | new_n22259_)) | (~new_n22258_ & ~new_n22259_ & new_n22260_)) & (new_n22261_ ^ ~new_n22262_));
  assign new_n22258_ = ~new_n22247_ & new_n22246_;
  assign new_n22259_ = ~new_n22249_ & new_n22248_;
  assign new_n22260_ = new_n22250_ & new_n22251_;
  assign new_n22261_ = (~new_n22254_ & new_n22253_) | (new_n22252_ & (~new_n22254_ | new_n22253_));
  assign new_n22262_ = new_n22255_ & new_n22256_;
  assign \o[27]  = (~new_n22260_ | ~new_n22261_ | ~new_n22262_ | (~new_n22258_ & ~new_n22259_)) & (new_n22260_ | new_n22261_ | new_n22262_) & (new_n22258_ | new_n22259_ | ((new_n22261_ | new_n22262_) & (new_n22260_ | (new_n22261_ & new_n22262_))));
  assign \o[28]  = new_n22265_ ? (new_n23275_ ^ new_n23325_) : (~new_n23275_ ^ new_n23325_);
  assign new_n22265_ = new_n22266_ ? (~new_n23181_ ^ new_n23197_) : (new_n23181_ ^ new_n23197_);
  assign new_n22266_ = new_n22267_ ? (new_n23126_ ^ new_n23165_) : (~new_n23126_ ^ new_n23165_);
  assign new_n22267_ = new_n22268_ ? (new_n22830_ ^ new_n23082_) : (~new_n22830_ ^ new_n23082_);
  assign new_n22268_ = new_n22269_ ? (new_n22535_ ^ new_n22792_) : (~new_n22535_ ^ new_n22792_);
  assign new_n22269_ = new_n22270_ ? (~new_n22434_ ^ new_n22463_) : (new_n22434_ ^ new_n22463_);
  assign new_n22270_ = new_n22271_ ? (new_n22350_ ^ new_n22377_) : (~new_n22350_ ^ new_n22377_);
  assign new_n22271_ = new_n22348_ & (new_n22349_ | ~new_n22272_);
  assign new_n22272_ = ~new_n22273_ & ~new_n22284_ & (~new_n22275_ | (new_n22324_ & new_n22320_) | (new_n22322_ & ~new_n22320_));
  assign new_n22273_ = new_n22274_ & new_n22283_;
  assign new_n22274_ = ~new_n22278_ & ~new_n22275_ & ~new_n22277_;
  assign new_n22275_ = ~new_n22276_ & ~new_n8854_;
  assign new_n22276_ = new_n11634_ & new_n8851_;
  assign new_n22277_ = ~new_n10368_ & new_n13406_;
  assign new_n22278_ = ~new_n20921_ & ~new_n20896_ & (~new_n20915_ | new_n22279_);
  assign new_n22279_ = new_n20922_ & (new_n20913_ | new_n20911_ | (~new_n20909_ & ~new_n22280_ & ~new_n20914_));
  assign new_n22280_ = new_n20904_ & ~new_n22281_ & new_n20905_;
  assign new_n22281_ = ~new_n20900_ & new_n20902_ & \all_features[782]  & \all_features[783]  & (~\all_features[781]  | new_n22282_);
  assign new_n22282_ = ~\all_features[779]  & ~\all_features[780]  & (~\all_features[778]  | new_n20907_);
  assign new_n22283_ = new_n20846_ & ~new_n19764_ & ~new_n19766_;
  assign new_n22284_ = new_n22285_ & ~new_n22286_ & ~new_n22319_;
  assign new_n22285_ = ~new_n22275_ & new_n22278_;
  assign new_n22286_ = ~new_n22287_ & new_n10773_;
  assign new_n22287_ = ~new_n22317_ & (new_n22314_ | new_n22288_ | new_n22308_ | new_n22311_ | ~new_n22318_);
  assign new_n22288_ = new_n22307_ & (new_n22313_ | (~new_n22312_ & new_n22302_ & (new_n22305_ | new_n22289_)));
  assign new_n22289_ = ~new_n22296_ & (~new_n22300_ | (new_n22290_ & (~new_n22299_ | (~new_n22301_ & new_n22293_))));
  assign new_n22290_ = \all_features[743]  & (\all_features[742]  | new_n22291_);
  assign new_n22291_ = \all_features[741]  & (\all_features[738]  | \all_features[739]  | \all_features[740]  | ~new_n22292_);
  assign new_n22292_ = ~\all_features[736]  & ~\all_features[737] ;
  assign new_n22293_ = \all_features[743]  & ~new_n22294_ & \all_features[742] ;
  assign new_n22294_ = ~\all_features[741]  & ~\all_features[740]  & ~\all_features[739]  & ~new_n22295_ & ~\all_features[738] ;
  assign new_n22295_ = \all_features[736]  & \all_features[737] ;
  assign new_n22296_ = ~\all_features[743]  & (~\all_features[742]  | ~new_n22297_ | ~new_n22295_ | ~new_n22298_);
  assign new_n22297_ = \all_features[738]  & \all_features[739] ;
  assign new_n22298_ = \all_features[740]  & \all_features[741] ;
  assign new_n22299_ = \all_features[743]  & (\all_features[742]  | (new_n22298_ & (\all_features[738]  | \all_features[739]  | \all_features[737] )));
  assign new_n22300_ = \all_features[743]  & (\all_features[741]  | \all_features[742]  | \all_features[740] );
  assign new_n22301_ = \all_features[742]  & \all_features[743]  & (\all_features[741]  | (\all_features[740]  & (\all_features[739]  | \all_features[738] )));
  assign new_n22302_ = ~new_n22296_ & ~new_n22305_ & (~new_n22300_ | new_n22303_ | ~new_n22290_);
  assign new_n22303_ = ~new_n22294_ & new_n22299_ & \all_features[742]  & \all_features[743]  & (~\all_features[741]  | new_n22304_);
  assign new_n22304_ = ~\all_features[739]  & ~\all_features[740]  & (~\all_features[738]  | new_n22292_);
  assign new_n22305_ = ~new_n22306_ & ~\all_features[743] ;
  assign new_n22306_ = \all_features[741]  & \all_features[742]  & (\all_features[740]  | (\all_features[738]  & \all_features[739]  & \all_features[737] ));
  assign new_n22307_ = ~new_n22311_ & ~new_n22308_ & ~new_n22310_;
  assign new_n22308_ = new_n22309_ & (~\all_features[741]  | (~\all_features[740]  & (~\all_features[739]  | (~\all_features[738]  & ~\all_features[737] ))));
  assign new_n22309_ = ~\all_features[742]  & ~\all_features[743] ;
  assign new_n22310_ = ~\all_features[741]  & new_n22309_ & ((~\all_features[738]  & new_n22292_) | ~\all_features[740]  | ~\all_features[739] );
  assign new_n22311_ = new_n22309_ & (~\all_features[739]  | ~new_n22298_ | (~\all_features[738]  & ~new_n22295_));
  assign new_n22312_ = ~\all_features[743]  & (~\all_features[742]  | (~\all_features[741]  & (new_n22292_ | ~new_n22297_ | ~\all_features[740] )));
  assign new_n22313_ = ~\all_features[743]  & (~\all_features[742]  | (~\all_features[740]  & ~\all_features[741]  & ~new_n22297_));
  assign new_n22314_ = ~new_n22305_ & ~new_n22312_ & new_n22316_ & (~new_n22290_ | ~new_n22315_);
  assign new_n22315_ = new_n22300_ & new_n22293_ & new_n22299_;
  assign new_n22316_ = ~new_n22296_ & ~new_n22313_;
  assign new_n22317_ = new_n22316_ & new_n22318_ & ~new_n22311_ & ~new_n22312_ & ~new_n22305_ & ~new_n22308_;
  assign new_n22318_ = ~new_n22310_ & (\all_features[739]  | \all_features[740]  | \all_features[741]  | \all_features[742]  | \all_features[743] );
  assign new_n22319_ = ~new_n10773_ & new_n21400_;
  assign new_n22320_ = ~new_n22321_ & new_n17588_;
  assign new_n22321_ = new_n17450_ & new_n8055_;
  assign new_n22322_ = new_n22323_ & new_n18109_ & new_n22321_;
  assign new_n22323_ = new_n17699_ & new_n20798_ & new_n17677_;
  assign new_n22324_ = ~new_n22341_ | ~new_n22345_ | ~new_n22346_ | (~new_n22344_ & new_n22335_);
  assign new_n22326_ = \all_features[3775]  & (\all_features[3774]  | new_n22327_);
  assign new_n22327_ = \all_features[3773]  & (\all_features[3770]  | \all_features[3771]  | \all_features[3772]  | ~new_n22328_);
  assign new_n22328_ = ~\all_features[3768]  & ~\all_features[3769] ;
  assign new_n22329_ = \all_features[3775]  & (\all_features[3774]  | (new_n22330_ & (\all_features[3770]  | \all_features[3771]  | \all_features[3769] )));
  assign new_n22330_ = \all_features[3772]  & \all_features[3773] ;
  assign new_n22331_ = new_n22333_ & (new_n22332_ | \all_features[3770]  | \all_features[3771]  | \all_features[3772]  | \all_features[3773] );
  assign new_n22332_ = \all_features[3768]  & \all_features[3769] ;
  assign new_n22333_ = \all_features[3774]  & \all_features[3775] ;
  assign new_n22335_ = new_n22336_ & (~new_n22326_ | ~new_n22329_ | ~new_n22331_);
  assign new_n22336_ = new_n22339_ & (\all_features[3775]  | (new_n22340_ & new_n22337_));
  assign new_n22337_ = \all_features[3774]  & (\all_features[3773]  | (~new_n22328_ & \all_features[3772]  & new_n22338_));
  assign new_n22338_ = \all_features[3770]  & \all_features[3771] ;
  assign new_n22339_ = \all_features[3775]  | (new_n22338_ & \all_features[3772]  & \all_features[3773]  & \all_features[3774]  & new_n22332_);
  assign new_n22340_ = \all_features[3773]  & \all_features[3774]  & (\all_features[3772]  | (\all_features[3770]  & \all_features[3771]  & \all_features[3769] ));
  assign new_n22341_ = \all_features[3774]  | \all_features[3775]  | (new_n22343_ & new_n22342_);
  assign new_n22342_ = new_n22330_ & \all_features[3771]  & (\all_features[3770]  | new_n22332_);
  assign new_n22343_ = \all_features[3773]  & (\all_features[3772]  | (\all_features[3771]  & (\all_features[3770]  | \all_features[3769] )));
  assign new_n22344_ = \all_features[3775]  | (new_n22330_ & new_n22340_ & new_n22338_ & \all_features[3774]  & new_n22332_);
  assign new_n22345_ = \all_features[3775]  | (\all_features[3774]  & (\all_features[3773]  | (~new_n22328_ & new_n22338_ & \all_features[3772] )));
  assign new_n22346_ = ~new_n22347_ | (\all_features[3771]  & \all_features[3772]  & (\all_features[3770]  | ~new_n22328_));
  assign new_n22347_ = ~\all_features[3775]  & ~\all_features[3773]  & ~\all_features[3774] ;
  assign new_n22348_ = (new_n22283_ | ~new_n22274_) & (~new_n22285_ | ~new_n22286_);
  assign new_n22349_ = (~new_n22324_ | ~new_n22320_ | ~new_n22275_) & (new_n22275_ | (new_n22278_ ? ~new_n22319_ : ~new_n22277_));
  assign new_n22350_ = ~new_n22351_ & new_n22375_;
  assign new_n22351_ = new_n22352_ & new_n22368_ & (new_n22370_ | new_n22373_ | new_n22364_ | new_n22365_);
  assign new_n22352_ = (new_n19338_ | new_n22366_ | ~new_n22364_) & (new_n22353_ | ~new_n22365_ | new_n22364_);
  assign new_n22353_ = (~new_n22354_ | ~new_n22362_) & (~new_n19708_ | ~new_n19712_ | ~new_n22363_ | new_n22362_);
  assign new_n22354_ = new_n22355_ & new_n22361_;
  assign new_n22355_ = ~new_n22356_ & ~new_n12984_;
  assign new_n22356_ = (new_n22357_ | (new_n13008_ & (~\all_features[1451]  | ~\all_features[1452]  | (~\all_features[1450]  & new_n12988_)))) & (~new_n13008_ | \all_features[1451]  | \all_features[1452] );
  assign new_n22357_ = ~new_n12997_ & (new_n12996_ | (~new_n13000_ & (new_n13002_ | (~new_n22358_ & ~new_n13005_))));
  assign new_n22358_ = ~new_n13004_ & (~\all_features[1455]  | new_n22359_ | (~\all_features[1452]  & ~\all_features[1453]  & ~\all_features[1454] ));
  assign new_n22359_ = \all_features[1455]  & ((~new_n22360_ & ~\all_features[1453]  & \all_features[1454] ) | (~new_n12990_ & (\all_features[1454]  | (~new_n12987_ & \all_features[1453] ))));
  assign new_n22360_ = (\all_features[1452]  & (\all_features[1450]  | \all_features[1451] )) | (~new_n12993_ & ~\all_features[1450]  & ~\all_features[1451]  & ~\all_features[1452] );
  assign new_n22361_ = ~new_n13009_ & ~new_n13012_;
  assign new_n22362_ = ~new_n6495_ & (~new_n6484_ | ~new_n6491_);
  assign new_n22363_ = new_n18396_ & new_n18412_;
  assign new_n22364_ = new_n13158_ & (new_n13136_ | ~new_n13159_);
  assign new_n22365_ = ~new_n9275_ & new_n9248_;
  assign new_n22366_ = new_n22367_ & (~new_n18985_ | (~new_n18962_ & ~new_n20442_));
  assign new_n22367_ = new_n18069_ & (new_n18046_ | (new_n18071_ & new_n18075_));
  assign new_n22368_ = ~new_n22369_ & (~new_n19338_ | ~new_n22364_ | (new_n22371_ ? new_n15873_ : new_n22372_));
  assign new_n22369_ = new_n22370_ & ~new_n22364_ & ~new_n22365_;
  assign new_n22370_ = new_n17012_ & new_n7126_;
  assign new_n22371_ = new_n6955_ & (new_n8545_ | new_n19232_);
  assign new_n22372_ = ~new_n13329_ & ~new_n21573_ & ~new_n21584_;
  assign new_n22373_ = ~new_n17012_ & new_n22374_;
  assign new_n22374_ = new_n6532_ & (new_n6529_ | new_n6521_);
  assign new_n22375_ = new_n22376_ & (~new_n22364_ | ((new_n22371_ | ~new_n22372_ | ~new_n19338_) & (~new_n22366_ | new_n19338_)));
  assign new_n22376_ = new_n22364_ | (new_n22365_ ? ~new_n22353_ : ~new_n22373_);
  assign new_n22377_ = ~new_n22378_ & new_n22430_;
  assign new_n22378_ = new_n22379_ & (~new_n22428_ | (new_n18632_ & ~new_n22429_) | (~new_n20116_ & new_n22429_));
  assign new_n22379_ = ~new_n22380_ & ~new_n22388_ & (~new_n22425_ | (new_n22426_ & new_n22427_) | (~new_n21853_ & ~new_n22427_));
  assign new_n22380_ = new_n22381_ & (new_n22385_ ? new_n22386_ : new_n22384_);
  assign new_n22381_ = ~new_n22382_ & ~new_n22383_;
  assign new_n22382_ = ~new_n8188_ & (~new_n8166_ | new_n15495_);
  assign new_n22383_ = new_n13009_ & new_n13012_;
  assign new_n22384_ = new_n7672_ & new_n7905_;
  assign new_n22385_ = ~new_n11378_ & new_n13845_;
  assign new_n22386_ = ~new_n22387_ & new_n6604_;
  assign new_n22387_ = new_n6630_ & new_n6634_;
  assign new_n22388_ = new_n22424_ & new_n16519_ & new_n22389_;
  assign new_n22389_ = new_n22390_ & new_n22419_;
  assign new_n22390_ = ~new_n22391_ & ~new_n22415_;
  assign new_n22391_ = new_n22412_ & (~new_n22406_ | (~new_n22392_ & ~new_n22410_ & ~new_n22414_));
  assign new_n22392_ = ~new_n22404_ & ~new_n22402_ & (~new_n22405_ | ~new_n22401_ | new_n22393_);
  assign new_n22393_ = new_n22394_ & new_n22398_ & (new_n22396_ | ~\all_features[2197]  | ~\all_features[2198]  | ~\all_features[2199] );
  assign new_n22394_ = \all_features[2199]  & (\all_features[2198]  | (new_n22395_ & (\all_features[2194]  | \all_features[2195]  | \all_features[2193] )));
  assign new_n22395_ = \all_features[2196]  & \all_features[2197] ;
  assign new_n22396_ = ~\all_features[2195]  & ~\all_features[2196]  & (~\all_features[2194]  | new_n22397_);
  assign new_n22397_ = ~\all_features[2192]  & ~\all_features[2193] ;
  assign new_n22398_ = \all_features[2198]  & \all_features[2199]  & (\all_features[2196]  | \all_features[2197]  | new_n22399_ | ~new_n22400_);
  assign new_n22399_ = \all_features[2192]  & \all_features[2193] ;
  assign new_n22400_ = ~\all_features[2194]  & ~\all_features[2195] ;
  assign new_n22401_ = \all_features[2199]  & (\all_features[2198]  | (\all_features[2197]  & (\all_features[2196]  | ~new_n22400_ | ~new_n22397_)));
  assign new_n22402_ = ~new_n22403_ & ~\all_features[2199] ;
  assign new_n22403_ = \all_features[2197]  & \all_features[2198]  & (\all_features[2196]  | (\all_features[2194]  & \all_features[2195]  & \all_features[2193] ));
  assign new_n22404_ = ~\all_features[2199]  & (~new_n22395_ | ~\all_features[2194]  | ~\all_features[2195]  | ~\all_features[2198]  | ~new_n22399_);
  assign new_n22405_ = \all_features[2199]  & (\all_features[2197]  | \all_features[2198]  | \all_features[2196] );
  assign new_n22406_ = ~new_n22407_ & ~new_n22409_;
  assign new_n22407_ = new_n22408_ & (~\all_features[2195]  | ~new_n22395_ | (~\all_features[2194]  & ~new_n22399_));
  assign new_n22408_ = ~\all_features[2198]  & ~\all_features[2199] ;
  assign new_n22409_ = new_n22408_ & (~\all_features[2197]  | (~\all_features[2196]  & (~\all_features[2195]  | (~\all_features[2194]  & ~\all_features[2193] ))));
  assign new_n22410_ = ~\all_features[2199]  & (~\all_features[2198]  | new_n22411_);
  assign new_n22411_ = ~\all_features[2197]  & (new_n22397_ | ~\all_features[2195]  | ~\all_features[2196]  | ~\all_features[2194] );
  assign new_n22412_ = ~new_n22413_ & (\all_features[2195]  | \all_features[2196]  | \all_features[2197]  | \all_features[2198]  | \all_features[2199] );
  assign new_n22413_ = ~\all_features[2197]  & new_n22408_ & ((~\all_features[2194]  & new_n22397_) | ~\all_features[2196]  | ~\all_features[2195] );
  assign new_n22414_ = ~\all_features[2199]  & (~\all_features[2198]  | (~\all_features[2197]  & ~\all_features[2196]  & (~\all_features[2195]  | ~\all_features[2194] )));
  assign new_n22415_ = ~new_n22416_ & (\all_features[2195]  | \all_features[2196]  | \all_features[2197]  | \all_features[2198]  | \all_features[2199] );
  assign new_n22416_ = ~new_n22413_ & (new_n22409_ | (~new_n22407_ & (new_n22414_ | (~new_n22410_ & ~new_n22417_))));
  assign new_n22417_ = ~new_n22402_ & (new_n22404_ | (new_n22405_ & (~new_n22401_ | (~new_n22418_ & new_n22394_))));
  assign new_n22418_ = ~\all_features[2197]  & \all_features[2198]  & \all_features[2199]  & (\all_features[2196]  ? new_n22400_ : (new_n22399_ | ~new_n22400_));
  assign new_n22419_ = ~new_n22420_ & ~new_n22423_;
  assign new_n22420_ = new_n22422_ & (~new_n22421_ | (new_n22401_ & new_n22405_ & new_n22394_ & new_n22398_));
  assign new_n22421_ = ~new_n22414_ & ~new_n22404_ & ~new_n22410_ & ~new_n22402_;
  assign new_n22422_ = new_n22406_ & new_n22412_;
  assign new_n22423_ = new_n22421_ & new_n22422_;
  assign new_n22424_ = new_n19844_ & new_n22383_;
  assign new_n22425_ = ~new_n22383_ & new_n22382_;
  assign new_n22426_ = new_n10970_ & (new_n10949_ | ~new_n15321_);
  assign new_n22427_ = ~new_n7869_ & new_n15319_;
  assign new_n22428_ = ~new_n19844_ & new_n22383_;
  assign new_n22429_ = new_n10726_ & (new_n10729_ | new_n10703_);
  assign new_n22430_ = new_n22431_ & (~new_n22428_ | (new_n20116_ & new_n22429_) | (~new_n18632_ & ~new_n22429_));
  assign new_n22431_ = new_n22432_ & (~new_n22425_ | (~new_n22426_ & new_n22427_) | (new_n21853_ & ~new_n22427_));
  assign new_n22432_ = ~new_n22433_ & (~new_n22381_ | (new_n22384_ & ~new_n22385_) | (new_n22386_ & new_n22385_));
  assign new_n22433_ = new_n22424_ & (new_n22389_ ? ~new_n16519_ : ~new_n6884_);
  assign new_n22434_ = ~new_n22435_ & new_n22453_;
  assign new_n22435_ = ~new_n15673_ & ((~new_n22436_ & ~new_n18579_) | (~new_n22452_ & new_n15873_ & new_n22387_ & new_n18579_));
  assign new_n22436_ = (new_n22437_ & ~new_n16453_) | (new_n22443_ & new_n16453_ & (~new_n22448_ | ~new_n22444_));
  assign new_n22437_ = ~new_n17357_ & (~new_n17353_ | ~new_n22438_ | ~new_n17330_);
  assign new_n22438_ = ~new_n17349_ & (new_n17346_ | (~new_n17352_ & (new_n17351_ | (~new_n17339_ & ~new_n22439_))));
  assign new_n22439_ = ~new_n17341_ & (new_n17342_ | (~new_n17344_ & (~new_n22442_ | new_n22440_)));
  assign new_n22440_ = \all_features[5047]  & ((~new_n22441_ & ~\all_features[5045]  & \all_features[5046] ) | (~new_n17336_ & (\all_features[5046]  | (~new_n17333_ & \all_features[5045] ))));
  assign new_n22441_ = (~\all_features[5042]  & ~\all_features[5043]  & ~\all_features[5044]  & (~\all_features[5041]  | ~\all_features[5040] )) | (\all_features[5044]  & (\all_features[5042]  | \all_features[5043] ));
  assign new_n22442_ = \all_features[5047]  & (\all_features[5045]  | \all_features[5046]  | \all_features[5044] );
  assign new_n22443_ = ~new_n20103_ & ~new_n15247_;
  assign new_n22444_ = ~new_n22445_ & ~new_n15260_;
  assign new_n22445_ = ~new_n15262_ & (new_n15256_ | (~new_n15252_ & (new_n15261_ | (~new_n15248_ & ~new_n22446_))));
  assign new_n22446_ = ~new_n15257_ & (new_n15263_ | (new_n20110_ & (~new_n20106_ | (~new_n22447_ & new_n20108_))));
  assign new_n22447_ = ~\all_features[1229]  & \all_features[1230]  & \all_features[1231]  & (\all_features[1228]  ? new_n20107_ : (new_n15254_ | ~new_n20107_));
  assign new_n22448_ = ~new_n15260_ & ~new_n15262_ & (~new_n15251_ | (~new_n15248_ & ~new_n22449_ & ~new_n15261_));
  assign new_n22449_ = ~new_n15257_ & ~new_n15263_ & (~new_n20110_ | ~new_n20106_ | new_n22450_);
  assign new_n22450_ = new_n20108_ & new_n20109_ & (new_n22451_ | ~\all_features[1229]  | ~\all_features[1230]  | ~\all_features[1231] );
  assign new_n22451_ = ~\all_features[1227]  & ~\all_features[1228]  & (~\all_features[1226]  | new_n15250_);
  assign new_n22452_ = ~new_n9686_ & (~new_n9679_ | new_n15023_);
  assign new_n22453_ = (~new_n22452_ | ~new_n22462_ | new_n15673_) & (~new_n15673_ | (new_n22459_ ? ~new_n22460_ : new_n22454_));
  assign new_n22454_ = (new_n22457_ & new_n7334_) ? (~new_n15477_ & new_n22458_) : new_n22455_;
  assign new_n22455_ = new_n14210_ & (new_n14207_ | ~new_n22456_);
  assign new_n22456_ = ~new_n15107_ & ~new_n14182_;
  assign new_n22457_ = new_n7305_ & new_n7327_;
  assign new_n22458_ = ~new_n15473_ & ~new_n15445_;
  assign new_n22459_ = new_n11612_ & (new_n11609_ | ~new_n11903_);
  assign new_n22460_ = ~new_n22461_ & new_n20308_;
  assign new_n22461_ = ~new_n13933_ & new_n13923_;
  assign new_n22462_ = new_n18579_ & new_n15308_ & (new_n15284_ | ~new_n15311_);
  assign new_n22463_ = new_n22531_ ? new_n22464_ : ((~new_n22533_ | new_n15282_) & (new_n17675_ | new_n22532_ | ~new_n15282_));
  assign new_n22464_ = ~new_n22465_ & (new_n17848_ | new_n22501_ | new_n22528_ | new_n22530_ | ~new_n10726_);
  assign new_n22465_ = ~new_n10726_ & new_n22500_ & (~new_n22466_ | new_n22498_) & (~new_n18626_ | new_n18619_);
  assign new_n22466_ = ~new_n22467_ & ~new_n22494_;
  assign new_n22467_ = new_n22491_ & (~new_n22487_ | (~new_n22468_ & new_n22484_));
  assign new_n22468_ = new_n22469_ & ((~new_n22476_ & new_n22481_ & new_n22482_) | ~new_n22483_ | ~new_n22479_);
  assign new_n22469_ = ~new_n22470_ & ~new_n22474_;
  assign new_n22470_ = ~\all_features[1703]  & (~\all_features[1702]  | ~new_n22471_ | ~new_n22472_ | ~new_n22473_);
  assign new_n22471_ = \all_features[1700]  & \all_features[1701] ;
  assign new_n22472_ = \all_features[1696]  & \all_features[1697] ;
  assign new_n22473_ = \all_features[1698]  & \all_features[1699] ;
  assign new_n22474_ = ~new_n22475_ & ~\all_features[1703] ;
  assign new_n22475_ = \all_features[1701]  & \all_features[1702]  & (\all_features[1700]  | (\all_features[1698]  & \all_features[1699]  & \all_features[1697] ));
  assign new_n22476_ = \all_features[1703]  & \all_features[1702]  & ~new_n22477_ & \all_features[1701] ;
  assign new_n22477_ = ~\all_features[1699]  & ~\all_features[1700]  & (~\all_features[1698]  | new_n22478_);
  assign new_n22478_ = ~\all_features[1696]  & ~\all_features[1697] ;
  assign new_n22479_ = \all_features[1703]  & (\all_features[1702]  | (\all_features[1701]  & (\all_features[1700]  | ~new_n22478_ | ~new_n22480_)));
  assign new_n22480_ = ~\all_features[1698]  & ~\all_features[1699] ;
  assign new_n22481_ = \all_features[1703]  & (\all_features[1702]  | (new_n22471_ & (\all_features[1698]  | \all_features[1699]  | \all_features[1697] )));
  assign new_n22482_ = \all_features[1702]  & \all_features[1703]  & (\all_features[1700]  | \all_features[1701]  | new_n22472_ | ~new_n22480_);
  assign new_n22483_ = \all_features[1703]  & (\all_features[1701]  | \all_features[1702]  | \all_features[1700] );
  assign new_n22484_ = ~new_n22485_ & ~new_n22486_;
  assign new_n22485_ = ~\all_features[1703]  & (~\all_features[1702]  | (~\all_features[1700]  & ~\all_features[1701]  & ~new_n22473_));
  assign new_n22486_ = ~\all_features[1703]  & (~\all_features[1702]  | (~\all_features[1701]  & (new_n22478_ | ~new_n22473_ | ~\all_features[1700] )));
  assign new_n22487_ = ~new_n22488_ & ~new_n22490_;
  assign new_n22488_ = new_n22489_ & (~\all_features[1699]  | ~new_n22471_ | (~\all_features[1698]  & ~new_n22472_));
  assign new_n22489_ = ~\all_features[1702]  & ~\all_features[1703] ;
  assign new_n22490_ = new_n22489_ & (~\all_features[1701]  | (~\all_features[1700]  & (~\all_features[1699]  | (~\all_features[1698]  & ~\all_features[1697] ))));
  assign new_n22491_ = ~new_n22492_ & ~new_n22493_;
  assign new_n22492_ = ~\all_features[1701]  & new_n22489_ & ((~\all_features[1698]  & new_n22478_) | ~\all_features[1700]  | ~\all_features[1699] );
  assign new_n22493_ = ~\all_features[1703]  & ~\all_features[1702]  & ~\all_features[1701]  & ~\all_features[1699]  & ~\all_features[1700] ;
  assign new_n22494_ = ~new_n22493_ & (new_n22492_ | new_n22495_);
  assign new_n22495_ = ~new_n22490_ & (new_n22488_ | (~new_n22485_ & (new_n22486_ | (~new_n22474_ & ~new_n22496_))));
  assign new_n22496_ = ~new_n22470_ & (~new_n22483_ | (new_n22479_ & (~new_n22481_ | (~new_n22497_ & new_n22482_))));
  assign new_n22497_ = \all_features[1702]  & \all_features[1703]  & (\all_features[1701]  | (~new_n22480_ & \all_features[1700] ));
  assign new_n22498_ = new_n22491_ & new_n22487_ & (~new_n22469_ | ~new_n22484_ | (new_n22499_ & new_n22479_));
  assign new_n22499_ = new_n22483_ & new_n22481_ & new_n22482_;
  assign new_n22500_ = new_n22491_ & new_n22487_ & new_n22484_ & new_n22469_;
  assign new_n22501_ = new_n22518_ & (~new_n22522_ | (~new_n22502_ & new_n22525_));
  assign new_n22502_ = new_n22503_ & ((~new_n22510_ & new_n22514_ & new_n22513_) | ~new_n22517_ | ~new_n22516_);
  assign new_n22503_ = ~new_n22504_ & ~new_n22506_;
  assign new_n22504_ = ~new_n22505_ & ~\all_features[2423] ;
  assign new_n22505_ = \all_features[2421]  & \all_features[2422]  & (\all_features[2420]  | (\all_features[2418]  & \all_features[2419]  & \all_features[2417] ));
  assign new_n22506_ = ~\all_features[2423]  & (~\all_features[2422]  | ~new_n22507_ | ~new_n22508_ | ~new_n22509_);
  assign new_n22507_ = \all_features[2416]  & \all_features[2417] ;
  assign new_n22508_ = \all_features[2420]  & \all_features[2421] ;
  assign new_n22509_ = \all_features[2418]  & \all_features[2419] ;
  assign new_n22510_ = \all_features[2423]  & \all_features[2422]  & ~new_n22511_ & \all_features[2421] ;
  assign new_n22511_ = ~\all_features[2419]  & ~\all_features[2420]  & (~\all_features[2418]  | new_n22512_);
  assign new_n22512_ = ~\all_features[2416]  & ~\all_features[2417] ;
  assign new_n22513_ = \all_features[2423]  & (\all_features[2422]  | (new_n22508_ & (\all_features[2418]  | \all_features[2419]  | \all_features[2417] )));
  assign new_n22514_ = \all_features[2422]  & \all_features[2423]  & (\all_features[2420]  | \all_features[2421]  | new_n22507_ | ~new_n22515_);
  assign new_n22515_ = ~\all_features[2418]  & ~\all_features[2419] ;
  assign new_n22516_ = \all_features[2423]  & (\all_features[2422]  | (\all_features[2421]  & (\all_features[2420]  | ~new_n22515_ | ~new_n22512_)));
  assign new_n22517_ = \all_features[2423]  & (\all_features[2421]  | \all_features[2422]  | \all_features[2420] );
  assign new_n22518_ = ~new_n22519_ & ~new_n22521_;
  assign new_n22519_ = ~\all_features[2421]  & new_n22520_ & ((~\all_features[2418]  & new_n22512_) | ~\all_features[2420]  | ~\all_features[2419] );
  assign new_n22520_ = ~\all_features[2422]  & ~\all_features[2423] ;
  assign new_n22521_ = ~\all_features[2423]  & ~\all_features[2422]  & ~\all_features[2421]  & ~\all_features[2419]  & ~\all_features[2420] ;
  assign new_n22522_ = ~new_n22523_ & ~new_n22524_;
  assign new_n22523_ = new_n22520_ & (~\all_features[2421]  | (~\all_features[2420]  & (~\all_features[2419]  | (~\all_features[2418]  & ~\all_features[2417] ))));
  assign new_n22524_ = new_n22520_ & (~\all_features[2419]  | ~new_n22508_ | (~\all_features[2418]  & ~new_n22507_));
  assign new_n22525_ = ~new_n22526_ & ~new_n22527_;
  assign new_n22526_ = ~\all_features[2423]  & (~\all_features[2422]  | (~\all_features[2420]  & ~\all_features[2421]  & ~new_n22509_));
  assign new_n22527_ = ~\all_features[2423]  & (~\all_features[2422]  | (~\all_features[2421]  & (new_n22512_ | ~new_n22509_ | ~\all_features[2420] )));
  assign new_n22528_ = new_n22518_ & new_n22522_ & (~new_n22503_ | ~new_n22525_ | (new_n22529_ & new_n22516_));
  assign new_n22529_ = new_n22517_ & new_n22513_ & new_n22514_;
  assign new_n22530_ = new_n22503_ & new_n22525_ & new_n22518_ & new_n22522_;
  assign new_n22531_ = ~new_n10775_ & (~new_n10776_ | new_n8298_);
  assign new_n22532_ = new_n9246_ & new_n15593_;
  assign new_n22533_ = ~new_n14681_ & new_n22534_ & (new_n11784_ | ~new_n11757_);
  assign new_n22534_ = new_n14656_ & new_n14679_;
  assign new_n22535_ = new_n22536_ ? (new_n22649_ ^ new_n22781_) : (~new_n22649_ ^ new_n22781_);
  assign new_n22536_ = new_n22537_ ^ new_n22598_;
  assign new_n22537_ = ~new_n22538_ & new_n22595_;
  assign new_n22538_ = new_n22539_ & ((~new_n22562_ & (new_n22551_ | (~new_n22547_ & ~new_n10910_ & new_n22541_))) | (new_n22551_ & (new_n10910_ | ~new_n22541_)));
  assign new_n22539_ = ~new_n22540_ & (new_n13887_ | ~new_n22544_ | ~new_n22545_);
  assign new_n22540_ = new_n22541_ & new_n10910_ & (~new_n18324_ | new_n8320_);
  assign new_n22541_ = ~new_n18099_ & new_n22542_;
  assign new_n22542_ = new_n20172_ & new_n22543_;
  assign new_n22543_ = ~new_n20202_ & ~new_n20205_;
  assign new_n22544_ = ~new_n21702_ & ~new_n22542_;
  assign new_n22545_ = new_n22466_ & new_n22546_;
  assign new_n22546_ = ~new_n22498_ & ~new_n22500_;
  assign new_n22547_ = new_n22548_ & new_n22544_ & new_n13887_;
  assign new_n22548_ = new_n22549_ & new_n22550_;
  assign new_n22549_ = ~new_n19782_ & ~new_n19802_;
  assign new_n22550_ = ~new_n19811_ & ~new_n19813_;
  assign new_n22551_ = new_n22542_ & ~new_n22552_ & new_n18099_;
  assign new_n22552_ = (~new_n17415_ | new_n17765_) & (new_n22553_ | ~new_n10610_ | ~new_n17765_);
  assign new_n22553_ = ~new_n22554_ & ~new_n22558_;
  assign new_n22554_ = ~new_n22555_ & (\all_features[3411]  | \all_features[3412]  | \all_features[3413]  | \all_features[3414]  | \all_features[3415] );
  assign new_n22555_ = ~new_n10630_ & (new_n10632_ | (~new_n10633_ & (new_n10623_ | (~new_n10627_ & ~new_n22556_))));
  assign new_n22556_ = ~new_n10621_ & (new_n10628_ | (new_n10619_ & (~new_n10625_ | (~new_n22557_ & new_n10614_))));
  assign new_n22557_ = ~\all_features[3413]  & \all_features[3414]  & \all_features[3415]  & (\all_features[3412]  ? new_n10617_ : (new_n10618_ | ~new_n10617_));
  assign new_n22558_ = new_n10629_ & (~new_n10635_ | (~new_n22559_ & ~new_n10623_ & ~new_n10627_));
  assign new_n22559_ = ~new_n10628_ & ~new_n10621_ & (~new_n10619_ | ~new_n10625_ | new_n22560_);
  assign new_n22560_ = new_n10614_ & new_n10616_ & (new_n22561_ | ~\all_features[3413]  | ~\all_features[3414]  | ~\all_features[3415] );
  assign new_n22561_ = ~\all_features[3411]  & ~\all_features[3412]  & (~\all_features[3410]  | new_n10626_);
  assign new_n22562_ = ~new_n22563_ & new_n22590_;
  assign new_n22563_ = ~new_n22589_ & (~new_n22582_ | (~new_n22587_ & (new_n22580_ | new_n22588_ | ~new_n22564_)));
  assign new_n22564_ = ~new_n22576_ & ~new_n22574_ & ((~new_n22571_ & new_n22565_) | ~new_n22579_ | ~new_n22578_);
  assign new_n22565_ = \all_features[1303]  & \all_features[1302]  & ~new_n22568_ & new_n22566_;
  assign new_n22566_ = \all_features[1303]  & (\all_features[1302]  | (new_n22567_ & (\all_features[1298]  | \all_features[1299]  | \all_features[1297] )));
  assign new_n22567_ = \all_features[1300]  & \all_features[1301] ;
  assign new_n22568_ = new_n22570_ & ~\all_features[1301]  & ~new_n22569_ & ~\all_features[1300] ;
  assign new_n22569_ = \all_features[1296]  & \all_features[1297] ;
  assign new_n22570_ = ~\all_features[1298]  & ~\all_features[1299] ;
  assign new_n22571_ = \all_features[1303]  & \all_features[1302]  & ~new_n22572_ & \all_features[1301] ;
  assign new_n22572_ = ~\all_features[1299]  & ~\all_features[1300]  & (~\all_features[1298]  | new_n22573_);
  assign new_n22573_ = ~\all_features[1296]  & ~\all_features[1297] ;
  assign new_n22574_ = ~new_n22575_ & ~\all_features[1303] ;
  assign new_n22575_ = \all_features[1301]  & \all_features[1302]  & (\all_features[1300]  | (\all_features[1298]  & \all_features[1299]  & \all_features[1297] ));
  assign new_n22576_ = ~\all_features[1303]  & (~\all_features[1302]  | ~new_n22577_ | ~new_n22569_ | ~new_n22567_);
  assign new_n22577_ = \all_features[1298]  & \all_features[1299] ;
  assign new_n22578_ = \all_features[1303]  & (\all_features[1302]  | (\all_features[1301]  & (\all_features[1300]  | ~new_n22570_ | ~new_n22573_)));
  assign new_n22579_ = \all_features[1303]  & (\all_features[1301]  | \all_features[1302]  | \all_features[1300] );
  assign new_n22580_ = ~new_n22574_ & (new_n22576_ | (new_n22579_ & (~new_n22578_ | (~new_n22581_ & new_n22566_))));
  assign new_n22581_ = ~\all_features[1301]  & \all_features[1302]  & \all_features[1303]  & (\all_features[1300]  ? new_n22570_ : (new_n22569_ | ~new_n22570_));
  assign new_n22582_ = ~new_n22586_ & ~new_n22583_ & ~new_n22585_;
  assign new_n22583_ = new_n22584_ & (~\all_features[1301]  | (~\all_features[1300]  & (~\all_features[1299]  | (~\all_features[1298]  & ~\all_features[1297] ))));
  assign new_n22584_ = ~\all_features[1302]  & ~\all_features[1303] ;
  assign new_n22585_ = ~\all_features[1301]  & new_n22584_ & ((~\all_features[1298]  & new_n22573_) | ~\all_features[1300]  | ~\all_features[1299] );
  assign new_n22586_ = new_n22584_ & (~\all_features[1299]  | ~new_n22567_ | (~\all_features[1298]  & ~new_n22569_));
  assign new_n22587_ = ~\all_features[1303]  & (~\all_features[1302]  | (~\all_features[1300]  & ~\all_features[1301]  & ~new_n22577_));
  assign new_n22588_ = ~\all_features[1303]  & (~\all_features[1302]  | (~\all_features[1301]  & (new_n22573_ | ~\all_features[1300]  | ~new_n22577_)));
  assign new_n22589_ = ~\all_features[1303]  & ~\all_features[1302]  & ~\all_features[1301]  & ~\all_features[1299]  & ~\all_features[1300] ;
  assign new_n22590_ = new_n22583_ | ~new_n22593_ | ((new_n22574_ | ~new_n22594_) & (new_n22591_ | new_n22586_));
  assign new_n22591_ = new_n22592_ & (~new_n22565_ | ~new_n22578_ | ~new_n22579_);
  assign new_n22592_ = ~new_n22576_ & ~new_n22574_ & ~new_n22587_ & ~new_n22588_;
  assign new_n22593_ = ~new_n22585_ & ~new_n22589_;
  assign new_n22594_ = ~new_n22586_ & ~new_n22576_ & ~new_n22587_ & ~new_n22588_;
  assign new_n22595_ = ~new_n22596_ & new_n22597_;
  assign new_n22596_ = ~new_n22542_ & ((~new_n22545_ & (~new_n13887_ | new_n21702_)) | (new_n13516_ & new_n21702_) | (~new_n22548_ & new_n13887_ & ~new_n21702_));
  assign new_n22597_ = (new_n13516_ | ~new_n21702_ | ~new_n22545_ | new_n22542_) & (~new_n22552_ | ~new_n18099_ | ~new_n22542_);
  assign new_n22598_ = ~new_n22599_ & new_n22646_;
  assign new_n22599_ = ~new_n22643_ & new_n22600_;
  assign new_n22600_ = (~new_n22603_ | ~new_n6698_) & (~new_n22609_ | ~new_n22604_) & (~new_n22601_ | ~new_n22607_);
  assign new_n22601_ = new_n22602_ & new_n12153_ & new_n15022_;
  assign new_n22602_ = ~new_n22448_ & new_n22443_;
  assign new_n22603_ = new_n22602_ & ~new_n9725_ & ~new_n15022_;
  assign new_n22604_ = new_n22605_ & ~new_n12841_ & ~new_n22602_;
  assign new_n22605_ = ~new_n22606_ & new_n18579_;
  assign new_n22606_ = new_n9347_ & new_n9371_;
  assign new_n22607_ = ~new_n6662_ & new_n22608_;
  assign new_n22608_ = ~new_n6640_ & ~new_n6670_;
  assign new_n22609_ = new_n22610_ & new_n22634_;
  assign new_n22610_ = ~new_n22611_ & ~new_n22633_;
  assign new_n22611_ = new_n22612_ & (~new_n22621_ | (new_n22631_ & new_n22632_ & new_n22628_ & new_n22630_));
  assign new_n22612_ = new_n22613_ & ~new_n22617_ & ~new_n22618_;
  assign new_n22613_ = ~new_n22614_ & (\all_features[4419]  | \all_features[4420]  | \all_features[4421]  | \all_features[4422]  | \all_features[4423] );
  assign new_n22614_ = ~\all_features[4421]  & new_n22616_ & ((~\all_features[4418]  & new_n22615_) | ~\all_features[4420]  | ~\all_features[4419] );
  assign new_n22615_ = ~\all_features[4416]  & ~\all_features[4417] ;
  assign new_n22616_ = ~\all_features[4422]  & ~\all_features[4423] ;
  assign new_n22617_ = new_n22616_ & (~\all_features[4421]  | (~\all_features[4420]  & (~\all_features[4419]  | (~\all_features[4418]  & ~\all_features[4417] ))));
  assign new_n22618_ = new_n22616_ & (~\all_features[4419]  | ~new_n22619_ | (~\all_features[4418]  & ~new_n22620_));
  assign new_n22619_ = \all_features[4420]  & \all_features[4421] ;
  assign new_n22620_ = \all_features[4416]  & \all_features[4417] ;
  assign new_n22621_ = ~new_n22627_ & ~new_n22626_ & ~new_n22622_ & ~new_n22624_;
  assign new_n22622_ = ~\all_features[4423]  & (~\all_features[4422]  | (~\all_features[4421]  & (new_n22615_ | ~new_n22623_ | ~\all_features[4420] )));
  assign new_n22623_ = \all_features[4418]  & \all_features[4419] ;
  assign new_n22624_ = ~new_n22625_ & ~\all_features[4423] ;
  assign new_n22625_ = \all_features[4421]  & \all_features[4422]  & (\all_features[4420]  | (\all_features[4418]  & \all_features[4419]  & \all_features[4417] ));
  assign new_n22626_ = ~\all_features[4423]  & (~\all_features[4422]  | ~new_n22619_ | ~new_n22620_ | ~new_n22623_);
  assign new_n22627_ = ~\all_features[4423]  & (~\all_features[4422]  | (~\all_features[4420]  & ~\all_features[4421]  & ~new_n22623_));
  assign new_n22628_ = \all_features[4423]  & (\all_features[4422]  | (\all_features[4421]  & (\all_features[4420]  | ~new_n22615_ | ~new_n22629_)));
  assign new_n22629_ = ~\all_features[4418]  & ~\all_features[4419] ;
  assign new_n22630_ = \all_features[4423]  & (\all_features[4422]  | (new_n22619_ & (\all_features[4418]  | \all_features[4419]  | \all_features[4417] )));
  assign new_n22631_ = \all_features[4422]  & \all_features[4423]  & (\all_features[4420]  | \all_features[4421]  | new_n22620_ | ~new_n22629_);
  assign new_n22632_ = \all_features[4423]  & (\all_features[4421]  | \all_features[4422]  | \all_features[4420] );
  assign new_n22633_ = new_n22612_ & new_n22621_;
  assign new_n22634_ = ~new_n22635_ & ~new_n22639_;
  assign new_n22635_ = new_n22613_ & (new_n22618_ | new_n22617_ | (~new_n22622_ & ~new_n22627_ & ~new_n22636_));
  assign new_n22636_ = ~new_n22626_ & ~new_n22624_ & (~new_n22632_ | ~new_n22628_ | new_n22637_);
  assign new_n22637_ = new_n22630_ & new_n22631_ & (new_n22638_ | ~\all_features[4421]  | ~\all_features[4422]  | ~\all_features[4423] );
  assign new_n22638_ = ~\all_features[4419]  & ~\all_features[4420]  & (~\all_features[4418]  | new_n22615_);
  assign new_n22639_ = ~new_n22640_ & (\all_features[4419]  | \all_features[4420]  | \all_features[4421]  | \all_features[4422]  | \all_features[4423] );
  assign new_n22640_ = ~new_n22614_ & (new_n22617_ | (~new_n22618_ & (new_n22627_ | (~new_n22622_ & ~new_n22641_))));
  assign new_n22641_ = ~new_n22624_ & (new_n22626_ | (new_n22632_ & (~new_n22628_ | (~new_n22642_ & new_n22630_))));
  assign new_n22642_ = ~\all_features[4421]  & \all_features[4422]  & \all_features[4423]  & (\all_features[4420]  ? new_n22629_ : (new_n22620_ | ~new_n22629_));
  assign new_n22643_ = ~new_n22602_ & ((new_n22644_ & ~new_n22605_) | (new_n12841_ & new_n22605_ & (new_n22645_ | ~new_n15762_)));
  assign new_n22644_ = new_n10948_ & new_n13349_;
  assign new_n22645_ = ~new_n15789_ & ~new_n15793_;
  assign new_n22646_ = ~new_n22647_ & new_n22648_ & (~new_n22603_ | new_n6698_) & (~new_n22601_ | new_n22607_);
  assign new_n22647_ = new_n22602_ & ((~new_n12153_ & new_n16479_ & new_n15022_) | (~new_n7409_ & new_n9725_ & ~new_n15022_));
  assign new_n22648_ = new_n22602_ | ((new_n12841_ | new_n22609_ | ~new_n22605_) & (new_n22644_ | new_n22605_));
  assign new_n22649_ = new_n22650_ ? (new_n22704_ ^ new_n22769_) : (~new_n22704_ ^ new_n22769_);
  assign new_n22650_ = ~new_n22651_ & new_n22699_;
  assign new_n22651_ = new_n22652_ & (~new_n22692_ | (~new_n13516_ & new_n22693_) | (~new_n22698_ & ~new_n22693_));
  assign new_n22652_ = new_n22653_ & (~new_n16762_ | ~new_n22655_ | new_n15751_ | new_n22386_);
  assign new_n22653_ = ~new_n22654_ & ((~new_n22691_ & new_n14392_) | ~new_n22655_ | ~new_n15751_);
  assign new_n22654_ = new_n18395_ & new_n22690_ & ~new_n22655_ & ~new_n22656_;
  assign new_n22655_ = ~new_n17178_ & new_n17153_;
  assign new_n22656_ = ~new_n22689_ & (~new_n22685_ | ~new_n22657_ | (~new_n22682_ & ~new_n22670_));
  assign new_n22657_ = new_n22658_ & (\all_features[5643]  | \all_features[5644]  | \all_features[5645]  | \all_features[5646]  | \all_features[5647] );
  assign new_n22658_ = new_n22669_ & new_n22676_ & (new_n22659_ | new_n22679_ | new_n22681_ | ~new_n22672_);
  assign new_n22659_ = new_n22668_ & new_n22666_ & new_n22660_ & new_n22663_;
  assign new_n22660_ = \all_features[5647]  & (\all_features[5646]  | new_n22661_);
  assign new_n22661_ = \all_features[5645]  & (\all_features[5642]  | \all_features[5643]  | \all_features[5644]  | ~new_n22662_);
  assign new_n22662_ = ~\all_features[5640]  & ~\all_features[5641] ;
  assign new_n22663_ = \all_features[5647]  & ~new_n22664_ & \all_features[5646] ;
  assign new_n22664_ = ~\all_features[5645]  & ~\all_features[5644]  & ~\all_features[5643]  & ~new_n22665_ & ~\all_features[5642] ;
  assign new_n22665_ = \all_features[5640]  & \all_features[5641] ;
  assign new_n22666_ = \all_features[5647]  & (\all_features[5646]  | (new_n22667_ & (\all_features[5642]  | \all_features[5643]  | \all_features[5641] )));
  assign new_n22667_ = \all_features[5644]  & \all_features[5645] ;
  assign new_n22668_ = \all_features[5647]  & (\all_features[5645]  | \all_features[5646]  | \all_features[5644] );
  assign new_n22669_ = ~new_n22670_ & (\all_features[5643]  | \all_features[5644]  | \all_features[5645]  | \all_features[5646]  | \all_features[5647] );
  assign new_n22670_ = ~\all_features[5645]  & new_n22671_ & ((~\all_features[5642]  & new_n22662_) | ~\all_features[5644]  | ~\all_features[5643] );
  assign new_n22671_ = ~\all_features[5646]  & ~\all_features[5647] ;
  assign new_n22672_ = ~new_n22673_ & ~new_n22675_;
  assign new_n22673_ = ~\all_features[5647]  & (~\all_features[5646]  | ~new_n22674_ | ~new_n22665_ | ~new_n22667_);
  assign new_n22674_ = \all_features[5642]  & \all_features[5643] ;
  assign new_n22675_ = ~\all_features[5647]  & (~\all_features[5646]  | (~\all_features[5644]  & ~\all_features[5645]  & ~new_n22674_));
  assign new_n22676_ = ~new_n22677_ & ~new_n22678_;
  assign new_n22677_ = new_n22671_ & (~\all_features[5645]  | (~\all_features[5644]  & (~\all_features[5643]  | (~\all_features[5642]  & ~\all_features[5641] ))));
  assign new_n22678_ = new_n22671_ & (~\all_features[5643]  | ~new_n22667_ | (~\all_features[5642]  & ~new_n22665_));
  assign new_n22679_ = ~new_n22680_ & ~\all_features[5647] ;
  assign new_n22680_ = \all_features[5645]  & \all_features[5646]  & (\all_features[5644]  | (\all_features[5642]  & \all_features[5643]  & \all_features[5641] ));
  assign new_n22681_ = ~\all_features[5647]  & (~\all_features[5646]  | (~\all_features[5645]  & (new_n22662_ | ~new_n22674_ | ~\all_features[5644] )));
  assign new_n22682_ = ~new_n22677_ & (new_n22678_ | (~new_n22675_ & (new_n22681_ | (~new_n22679_ & ~new_n22683_))));
  assign new_n22683_ = ~new_n22673_ & (~new_n22668_ | (new_n22660_ & (~new_n22666_ | (~new_n22684_ & new_n22663_))));
  assign new_n22684_ = \all_features[5646]  & \all_features[5647]  & (\all_features[5645]  | (\all_features[5644]  & (\all_features[5643]  | \all_features[5642] )));
  assign new_n22685_ = new_n22669_ & (~new_n22676_ | (~new_n22686_ & ~new_n22681_ & ~new_n22675_));
  assign new_n22686_ = ~new_n22673_ & ~new_n22679_ & (~new_n22668_ | new_n22687_ | ~new_n22660_);
  assign new_n22687_ = ~new_n22664_ & new_n22666_ & \all_features[5646]  & \all_features[5647]  & (~\all_features[5645]  | new_n22688_);
  assign new_n22688_ = ~\all_features[5643]  & ~\all_features[5644]  & (~\all_features[5642]  | new_n22662_);
  assign new_n22689_ = new_n22672_ & new_n22669_ & ~new_n22678_ & ~new_n22681_ & ~new_n22679_ & ~new_n22677_;
  assign new_n22690_ = ~new_n21345_ & ~new_n21334_ & ~new_n21343_;
  assign new_n22691_ = new_n10610_ & new_n22558_;
  assign new_n22692_ = ~new_n22655_ & ~new_n18395_;
  assign new_n22693_ = new_n15531_ & (new_n15093_ | (~new_n15090_ & (new_n15104_ | new_n22694_)));
  assign new_n22694_ = ~new_n15103_ & (new_n15101_ | (~new_n15102_ & (new_n15095_ | (~new_n15097_ & ~new_n22695_))));
  assign new_n22695_ = ~new_n22696_ & \all_features[1503]  & (\all_features[1502]  | \all_features[1501]  | \all_features[1500] );
  assign new_n22696_ = \all_features[1503]  & ((~new_n22697_ & ~\all_features[1501]  & \all_features[1502] ) | (~new_n15358_ & (\all_features[1502]  | (~new_n15355_ & \all_features[1501] ))));
  assign new_n22697_ = (\all_features[1500]  & ~new_n15356_) | (~new_n15099_ & ~\all_features[1500]  & new_n15356_);
  assign new_n22698_ = ~new_n9423_ & new_n21056_;
  assign new_n22699_ = new_n22700_ & new_n22703_ & (~new_n22692_ | (new_n13516_ & new_n22693_) | (new_n22698_ & ~new_n22693_));
  assign new_n22700_ = (~new_n18395_ | new_n22701_ | new_n22655_) & (new_n15751_ | new_n22702_ | ~new_n22386_ | ~new_n22655_);
  assign new_n22701_ = new_n22690_ ? ~new_n22656_ : new_n13837_;
  assign new_n22702_ = ~new_n18951_ & ~new_n18953_;
  assign new_n22703_ = ~new_n22655_ | ((new_n22691_ | ~new_n14392_ | ~new_n15751_) & (new_n16762_ | new_n22386_ | new_n15751_));
  assign new_n22704_ = new_n20882_ ? ((new_n22768_ | ~new_n15479_) & (new_n15481_ | ~new_n19821_ | new_n15479_)) : new_n22705_;
  assign new_n22705_ = new_n22710_ ? new_n22706_ : ~new_n22712_;
  assign new_n22706_ = (~new_n22707_ & new_n22709_) | (new_n18069_ & ~new_n22709_ & (new_n18075_ | new_n18046_));
  assign new_n22707_ = ~new_n7736_ & new_n22708_;
  assign new_n22708_ = ~new_n7722_ & ~new_n7733_;
  assign new_n22709_ = ~new_n7432_ & (~new_n7438_ | ~new_n7410_);
  assign new_n22710_ = new_n14528_ & (new_n14505_ | ~new_n22711_);
  assign new_n22711_ = ~new_n14531_ & ~new_n14535_;
  assign new_n22712_ = ~new_n22713_ & (new_n22767_ | (~new_n22759_ & new_n22741_));
  assign new_n22713_ = new_n22734_ & (new_n22714_ | (~new_n22729_ & ~new_n22733_ & (~new_n22736_ | new_n22737_)));
  assign new_n22714_ = ~new_n22733_ & ~new_n22732_ & ~new_n22731_ & ~new_n22715_ & ~new_n22729_;
  assign new_n22715_ = ~new_n22728_ & ~new_n22727_ & ~new_n22725_ & ~new_n22716_ & ~new_n22723_;
  assign new_n22716_ = \all_features[1775]  & \all_features[1774]  & ~new_n22721_ & new_n22719_;
  assign new_n22717_ = \all_features[1773]  & (\all_features[1770]  | \all_features[1771]  | \all_features[1772]  | ~new_n22718_);
  assign new_n22718_ = ~\all_features[1768]  & ~\all_features[1769] ;
  assign new_n22719_ = \all_features[1775]  & (\all_features[1774]  | (new_n22720_ & (\all_features[1770]  | \all_features[1771]  | \all_features[1769] )));
  assign new_n22720_ = \all_features[1772]  & \all_features[1773] ;
  assign new_n22721_ = ~\all_features[1773]  & ~\all_features[1772]  & ~\all_features[1771]  & ~new_n22722_ & ~\all_features[1770] ;
  assign new_n22722_ = \all_features[1768]  & \all_features[1769] ;
  assign new_n22723_ = ~new_n22724_ & ~\all_features[1775] ;
  assign new_n22724_ = \all_features[1773]  & \all_features[1774]  & (\all_features[1772]  | (\all_features[1770]  & \all_features[1771]  & \all_features[1769] ));
  assign new_n22725_ = ~\all_features[1775]  & (~\all_features[1774]  | ~new_n22722_ | ~new_n22720_ | ~new_n22726_);
  assign new_n22726_ = \all_features[1770]  & \all_features[1771] ;
  assign new_n22727_ = ~\all_features[1775]  & (~\all_features[1774]  | (~\all_features[1772]  & ~\all_features[1773]  & ~new_n22726_));
  assign new_n22728_ = ~\all_features[1775]  & (~\all_features[1774]  | (~\all_features[1773]  & (new_n22718_ | ~\all_features[1772]  | ~new_n22726_)));
  assign new_n22729_ = ~\all_features[1773]  & new_n22730_ & ((~\all_features[1770]  & new_n22718_) | ~\all_features[1772]  | ~\all_features[1771] );
  assign new_n22730_ = ~\all_features[1774]  & ~\all_features[1775] ;
  assign new_n22731_ = new_n22730_ & (~\all_features[1771]  | ~new_n22720_ | (~\all_features[1770]  & ~new_n22722_));
  assign new_n22732_ = new_n22730_ & (~\all_features[1773]  | (~\all_features[1772]  & (~\all_features[1771]  | (~\all_features[1770]  & ~\all_features[1769] ))));
  assign new_n22733_ = ~\all_features[1775]  & ~\all_features[1774]  & ~\all_features[1773]  & ~\all_features[1771]  & ~\all_features[1772] ;
  assign new_n22734_ = new_n22736_ & new_n22735_ & ~new_n22728_ & ~new_n22729_ & ~new_n22723_ & ~new_n22727_;
  assign new_n22735_ = ~new_n22725_ & ~new_n22733_;
  assign new_n22736_ = ~new_n22731_ & ~new_n22732_;
  assign new_n22737_ = ~new_n22727_ & ~new_n22728_ & ((~new_n22739_ & new_n22738_) | new_n22725_ | new_n22723_);
  assign new_n22738_ = \all_features[1775]  & (\all_features[1774]  | new_n22717_);
  assign new_n22739_ = ~new_n22721_ & new_n22719_ & \all_features[1774]  & \all_features[1775]  & (~\all_features[1773]  | new_n22740_);
  assign new_n22740_ = ~\all_features[1771]  & ~\all_features[1772]  & (~\all_features[1770]  | new_n22718_);
  assign new_n22741_ = new_n22759_ & (new_n22763_ | (~new_n22764_ & new_n22742_ & (new_n22751_ | new_n22757_)));
  assign new_n22742_ = ~new_n22751_ & ~new_n22753_ & (~new_n22756_ | ~new_n22755_ | new_n22743_);
  assign new_n22743_ = new_n22744_ & ~new_n22749_ & new_n22746_;
  assign new_n22744_ = \all_features[3567]  & (\all_features[3566]  | (new_n22745_ & (\all_features[3562]  | \all_features[3563]  | \all_features[3561] )));
  assign new_n22745_ = \all_features[3564]  & \all_features[3565] ;
  assign new_n22746_ = new_n22748_ & (\all_features[3564]  | \all_features[3565]  | ~new_n22747_ | (\all_features[3561]  & \all_features[3560] ));
  assign new_n22747_ = ~\all_features[3562]  & ~\all_features[3563] ;
  assign new_n22748_ = \all_features[3566]  & \all_features[3567] ;
  assign new_n22749_ = new_n22748_ & \all_features[3565]  & ((~new_n22750_ & \all_features[3562] ) | \all_features[3564]  | \all_features[3563] );
  assign new_n22750_ = ~\all_features[3560]  & ~\all_features[3561] ;
  assign new_n22751_ = ~new_n22752_ & ~\all_features[3567] ;
  assign new_n22752_ = \all_features[3565]  & \all_features[3566]  & (\all_features[3564]  | (\all_features[3562]  & \all_features[3563]  & \all_features[3561] ));
  assign new_n22753_ = ~\all_features[3567]  & (~new_n22745_ | ~\all_features[3560]  | ~\all_features[3561]  | ~\all_features[3566]  | ~new_n22754_);
  assign new_n22754_ = \all_features[3562]  & \all_features[3563] ;
  assign new_n22755_ = \all_features[3567]  & (\all_features[3566]  | (\all_features[3565]  & (\all_features[3564]  | ~new_n22747_ | ~new_n22750_)));
  assign new_n22756_ = \all_features[3567]  & (\all_features[3565]  | \all_features[3566]  | \all_features[3564] );
  assign new_n22757_ = ~new_n22753_ & (~new_n22756_ | (new_n22755_ & (~new_n22744_ | (~new_n22758_ & new_n22746_))));
  assign new_n22758_ = new_n22748_ & (\all_features[3565]  | (~new_n22747_ & \all_features[3564] ));
  assign new_n22759_ = \all_features[3566]  | \all_features[3567]  | (~new_n22762_ & new_n22761_ & \all_features[3565] );
  assign new_n22761_ = new_n22745_ & \all_features[3563]  & (\all_features[3562]  | (\all_features[3560]  & \all_features[3561] ));
  assign new_n22762_ = ~\all_features[3564]  & (~\all_features[3563]  | (~\all_features[3562]  & ~\all_features[3561] ));
  assign new_n22763_ = ~\all_features[3567]  & (~\all_features[3566]  | (~\all_features[3564]  & ~\all_features[3565]  & ~new_n22754_));
  assign new_n22764_ = ~\all_features[3567]  & (~\all_features[3566]  | (~\all_features[3565]  & (new_n22750_ | ~\all_features[3564]  | ~new_n22754_)));
  assign new_n22767_ = ~\all_features[3567]  & ~\all_features[3566]  & ~\all_features[3565]  & ~\all_features[3563]  & ~\all_features[3564] ;
  assign new_n22768_ = ~new_n13012_ & new_n15328_ & new_n12983_ & (~new_n10972_ | ~new_n15322_);
  assign new_n22769_ = ~new_n22770_ & new_n22777_ & (new_n22776_ | new_n22771_ | new_n19802_ | ~new_n22550_);
  assign new_n22770_ = ~new_n22771_ & ~new_n22773_ & (new_n22774_ ? ~new_n22775_ : (~new_n22734_ | ~new_n22714_));
  assign new_n22771_ = ~new_n12525_ & new_n22772_;
  assign new_n22772_ = ~new_n12514_ & ~new_n12523_;
  assign new_n22773_ = ~new_n19802_ & new_n22550_;
  assign new_n22774_ = ~new_n13505_ & new_n20883_;
  assign new_n22775_ = new_n9340_ & (new_n9314_ | new_n15042_);
  assign new_n22776_ = new_n14013_ ? new_n11905_ : (new_n7832_ | (~new_n16900_ & new_n7830_));
  assign new_n22777_ = ~new_n22771_ | ((~new_n15169_ | ~new_n22778_) & (~new_n22780_ | new_n22778_ | (~new_n6491_ & new_n20242_)));
  assign new_n22778_ = ~new_n22779_ & new_n11615_;
  assign new_n22779_ = new_n7188_ & new_n11617_;
  assign new_n22780_ = ~new_n14416_ & new_n6495_;
  assign new_n22781_ = new_n22783_ & (new_n12187_ | (new_n22782_ & new_n20171_) | (new_n22791_ & ~new_n20171_));
  assign new_n22782_ = new_n19147_ ? new_n15320_ : ~new_n8408_;
  assign new_n22783_ = ~new_n12187_ | ((new_n22784_ | new_n15669_) & (new_n22785_ | ~new_n15669_ | (new_n15745_ & ~new_n22790_)));
  assign new_n22784_ = new_n9547_ ? (new_n11704_ | (new_n18460_ & new_n18470_)) : ~new_n14038_;
  assign new_n22785_ = ~new_n22786_ & new_n21536_;
  assign new_n22786_ = new_n21539_ & (new_n21544_ | new_n21543_ | (~new_n21548_ & ~new_n21553_ & ~new_n22787_));
  assign new_n22787_ = ~new_n21552_ & ~new_n21550_ & (~new_n21558_ | ~new_n21554_ | new_n22788_);
  assign new_n22788_ = new_n21556_ & new_n21557_ & (new_n22789_ | ~\all_features[4637]  | ~\all_features[4638]  | ~\all_features[4639] );
  assign new_n22789_ = ~\all_features[4635]  & ~\all_features[4636]  & (~\all_features[4634]  | new_n21541_);
  assign new_n22790_ = ~new_n15717_ & ~new_n15743_;
  assign new_n22791_ = new_n14655_ ? ~new_n18189_ : ~new_n13064_;
  assign new_n22792_ = new_n22797_ ? (new_n22793_ & (new_n22794_ | new_n10936_ | ~new_n20842_)) : new_n22796_;
  assign new_n22793_ = (new_n19425_ | ~new_n7698_ | ~new_n22794_) & (~new_n19162_ | ~new_n10936_ | new_n22794_);
  assign new_n22794_ = ~new_n14813_ & new_n22795_;
  assign new_n22795_ = new_n14843_ & new_n14845_;
  assign new_n22796_ = new_n20969_ & new_n14923_;
  assign new_n22797_ = ~new_n22798_ & new_n22825_;
  assign new_n22798_ = ~new_n22824_ & (~new_n22817_ | (~new_n22822_ & (new_n22815_ | new_n22823_ | ~new_n22799_)));
  assign new_n22799_ = ~new_n22811_ & ~new_n22809_ & ((~new_n22806_ & new_n22800_) | ~new_n22814_ | ~new_n22813_);
  assign new_n22800_ = \all_features[5919]  & \all_features[5918]  & ~new_n22803_ & new_n22801_;
  assign new_n22801_ = \all_features[5919]  & (\all_features[5918]  | (new_n22802_ & (\all_features[5914]  | \all_features[5915]  | \all_features[5913] )));
  assign new_n22802_ = \all_features[5916]  & \all_features[5917] ;
  assign new_n22803_ = new_n22805_ & ~\all_features[5917]  & ~new_n22804_ & ~\all_features[5916] ;
  assign new_n22804_ = \all_features[5912]  & \all_features[5913] ;
  assign new_n22805_ = ~\all_features[5914]  & ~\all_features[5915] ;
  assign new_n22806_ = \all_features[5919]  & \all_features[5918]  & ~new_n22807_ & \all_features[5917] ;
  assign new_n22807_ = ~\all_features[5915]  & ~\all_features[5916]  & (~\all_features[5914]  | new_n22808_);
  assign new_n22808_ = ~\all_features[5912]  & ~\all_features[5913] ;
  assign new_n22809_ = ~new_n22810_ & ~\all_features[5919] ;
  assign new_n22810_ = \all_features[5917]  & \all_features[5918]  & (\all_features[5916]  | (\all_features[5914]  & \all_features[5915]  & \all_features[5913] ));
  assign new_n22811_ = ~\all_features[5919]  & (~\all_features[5918]  | ~new_n22812_ | ~new_n22804_ | ~new_n22802_);
  assign new_n22812_ = \all_features[5914]  & \all_features[5915] ;
  assign new_n22813_ = \all_features[5919]  & (\all_features[5918]  | (\all_features[5917]  & (\all_features[5916]  | ~new_n22805_ | ~new_n22808_)));
  assign new_n22814_ = \all_features[5919]  & (\all_features[5917]  | \all_features[5918]  | \all_features[5916] );
  assign new_n22815_ = ~new_n22809_ & (new_n22811_ | (new_n22814_ & (~new_n22813_ | (~new_n22816_ & new_n22801_))));
  assign new_n22816_ = ~\all_features[5917]  & \all_features[5918]  & \all_features[5919]  & (\all_features[5916]  ? new_n22805_ : (new_n22804_ | ~new_n22805_));
  assign new_n22817_ = ~new_n22821_ & ~new_n22818_ & ~new_n22820_;
  assign new_n22818_ = new_n22819_ & (~\all_features[5917]  | (~\all_features[5916]  & (~\all_features[5915]  | (~\all_features[5914]  & ~\all_features[5913] ))));
  assign new_n22819_ = ~\all_features[5918]  & ~\all_features[5919] ;
  assign new_n22820_ = ~\all_features[5917]  & new_n22819_ & ((~\all_features[5914]  & new_n22808_) | ~\all_features[5916]  | ~\all_features[5915] );
  assign new_n22821_ = new_n22819_ & (~\all_features[5915]  | ~new_n22802_ | (~\all_features[5914]  & ~new_n22804_));
  assign new_n22822_ = ~\all_features[5919]  & (~\all_features[5918]  | (~\all_features[5916]  & ~\all_features[5917]  & ~new_n22812_));
  assign new_n22823_ = ~\all_features[5919]  & (~\all_features[5918]  | (~\all_features[5917]  & (new_n22808_ | ~\all_features[5916]  | ~new_n22812_)));
  assign new_n22824_ = ~\all_features[5919]  & ~\all_features[5918]  & ~\all_features[5917]  & ~\all_features[5915]  & ~\all_features[5916] ;
  assign new_n22825_ = new_n22818_ | ~new_n22828_ | ((new_n22809_ | ~new_n22829_) & (new_n22826_ | new_n22821_));
  assign new_n22826_ = new_n22827_ & (~new_n22800_ | ~new_n22813_ | ~new_n22814_);
  assign new_n22827_ = ~new_n22811_ & ~new_n22809_ & ~new_n22822_ & ~new_n22823_;
  assign new_n22828_ = ~new_n22820_ & ~new_n22824_;
  assign new_n22829_ = ~new_n22821_ & ~new_n22811_ & ~new_n22822_ & ~new_n22823_;
  assign new_n22830_ = new_n22831_ ? (~new_n23060_ ^ new_n23073_) : (new_n23060_ ^ new_n23073_);
  assign new_n22831_ = new_n22832_ ? (new_n22943_ ^ new_n22999_) : (~new_n22943_ ^ new_n22999_);
  assign new_n22832_ = new_n22833_ ? (new_n22895_ ^ new_n22935_) : (~new_n22895_ ^ new_n22935_);
  assign new_n22833_ = new_n22834_ & (new_n22840_ | ~new_n22839_ | (new_n10910_ ? ~new_n20085_ : new_n22879_));
  assign new_n22834_ = new_n22835_ & (new_n22839_ | ~new_n15169_ | ~new_n7445_ | (new_n12685_ & new_n22877_));
  assign new_n22835_ = (~new_n22840_ | new_n22836_ | ~new_n22839_) & (new_n22841_ | new_n15169_ | ~new_n22876_ | new_n22839_);
  assign new_n22836_ = ~new_n22838_ & new_n22837_;
  assign new_n22837_ = new_n15166_ & new_n20048_;
  assign new_n22838_ = new_n10677_ & new_n10679_;
  assign new_n22839_ = ~new_n18290_ & new_n18321_;
  assign new_n22840_ = ~new_n7870_ & new_n16647_;
  assign new_n22841_ = ~new_n22872_ & (~new_n22863_ | ~new_n22842_ | ~new_n22874_);
  assign new_n22842_ = ~new_n22843_ & (\all_features[1875]  | \all_features[1876]  | \all_features[1877]  | \all_features[1878]  | \all_features[1879] );
  assign new_n22843_ = ~new_n22858_ & (new_n22860_ | (~new_n22861_ & (new_n22857_ | (~new_n22844_ & ~new_n22862_))));
  assign new_n22844_ = ~new_n22845_ & (new_n22847_ | (new_n22856_ & (~new_n22851_ | (~new_n22855_ & new_n22854_))));
  assign new_n22845_ = ~new_n22846_ & ~\all_features[1879] ;
  assign new_n22846_ = \all_features[1877]  & \all_features[1878]  & (\all_features[1876]  | (\all_features[1874]  & \all_features[1875]  & \all_features[1873] ));
  assign new_n22847_ = ~\all_features[1879]  & (~\all_features[1878]  | ~new_n22848_ | ~new_n22849_ | ~new_n22850_);
  assign new_n22848_ = \all_features[1872]  & \all_features[1873] ;
  assign new_n22849_ = \all_features[1876]  & \all_features[1877] ;
  assign new_n22850_ = \all_features[1874]  & \all_features[1875] ;
  assign new_n22851_ = \all_features[1879]  & (\all_features[1878]  | (\all_features[1877]  & (\all_features[1876]  | ~new_n22853_ | ~new_n22852_)));
  assign new_n22852_ = ~\all_features[1872]  & ~\all_features[1873] ;
  assign new_n22853_ = ~\all_features[1874]  & ~\all_features[1875] ;
  assign new_n22854_ = \all_features[1879]  & (\all_features[1878]  | (new_n22849_ & (\all_features[1874]  | \all_features[1875]  | \all_features[1873] )));
  assign new_n22855_ = ~\all_features[1877]  & \all_features[1878]  & \all_features[1879]  & (\all_features[1876]  ? new_n22853_ : (new_n22848_ | ~new_n22853_));
  assign new_n22856_ = \all_features[1879]  & (\all_features[1877]  | \all_features[1878]  | \all_features[1876] );
  assign new_n22857_ = ~\all_features[1879]  & (~\all_features[1878]  | (~\all_features[1876]  & ~\all_features[1877]  & ~new_n22850_));
  assign new_n22858_ = ~\all_features[1877]  & new_n22859_ & ((~\all_features[1874]  & new_n22852_) | ~\all_features[1876]  | ~\all_features[1875] );
  assign new_n22859_ = ~\all_features[1878]  & ~\all_features[1879] ;
  assign new_n22860_ = new_n22859_ & (~\all_features[1877]  | (~\all_features[1876]  & (~\all_features[1875]  | (~\all_features[1874]  & ~\all_features[1873] ))));
  assign new_n22861_ = new_n22859_ & (~\all_features[1875]  | ~new_n22849_ | (~\all_features[1874]  & ~new_n22848_));
  assign new_n22862_ = ~\all_features[1879]  & (~\all_features[1878]  | (~\all_features[1877]  & (new_n22852_ | ~\all_features[1876]  | ~new_n22850_)));
  assign new_n22863_ = new_n22871_ & (~new_n22869_ | (~new_n22864_ & new_n22870_));
  assign new_n22864_ = new_n22867_ & ((~new_n22865_ & new_n22854_ & new_n22868_) | ~new_n22856_ | ~new_n22851_);
  assign new_n22865_ = \all_features[1879]  & \all_features[1878]  & ~new_n22866_ & \all_features[1877] ;
  assign new_n22866_ = ~\all_features[1875]  & ~\all_features[1876]  & (~\all_features[1874]  | new_n22852_);
  assign new_n22867_ = ~new_n22845_ & ~new_n22847_;
  assign new_n22868_ = \all_features[1878]  & \all_features[1879]  & (\all_features[1876]  | \all_features[1877]  | new_n22848_ | ~new_n22853_);
  assign new_n22869_ = ~new_n22860_ & ~new_n22861_;
  assign new_n22870_ = ~new_n22857_ & ~new_n22862_;
  assign new_n22871_ = ~new_n22858_ & (\all_features[1875]  | \all_features[1876]  | \all_features[1877]  | \all_features[1878]  | \all_features[1879] );
  assign new_n22872_ = new_n22869_ & new_n22873_ & ~new_n22862_ & ~new_n22858_ & ~new_n22845_ & ~new_n22857_;
  assign new_n22873_ = ~new_n22847_ & (\all_features[1875]  | \all_features[1876]  | \all_features[1877]  | \all_features[1878]  | \all_features[1879] );
  assign new_n22874_ = new_n22869_ & new_n22871_ & (~new_n22870_ | ~new_n22867_ | (new_n22875_ & new_n22851_));
  assign new_n22875_ = new_n22856_ & new_n22854_ & new_n22868_;
  assign new_n22876_ = new_n13918_ & new_n13921_;
  assign new_n22877_ = new_n22878_ & new_n12682_;
  assign new_n22878_ = new_n12627_ & new_n12651_;
  assign new_n22879_ = new_n19318_ & (new_n22893_ | new_n22880_);
  assign new_n22880_ = ~new_n19327_ & ~new_n19330_ & ~new_n19320_ & ~new_n22881_ & ~new_n22887_;
  assign new_n22881_ = ~new_n19325_ & (new_n19322_ | (~new_n19333_ & (new_n19328_ | (~new_n22882_ & ~new_n19332_))));
  assign new_n22882_ = ~new_n22883_ & \all_features[4199]  & (\all_features[4198]  | \all_features[4197]  | \all_features[4196] );
  assign new_n22883_ = \all_features[4199]  & ((~new_n22886_ & ~\all_features[4197]  & \all_features[4198] ) | (~new_n22885_ & (\all_features[4198]  | (~new_n22884_ & \all_features[4197] ))));
  assign new_n22884_ = new_n19331_ & ~\all_features[4196]  & ~\all_features[4194]  & ~\all_features[4195] ;
  assign new_n22885_ = \all_features[4199]  & (\all_features[4198]  | (new_n19326_ & (\all_features[4194]  | \all_features[4195]  | \all_features[4193] )));
  assign new_n22886_ = (~\all_features[4194]  & ~\all_features[4195]  & ~\all_features[4196]  & (~\all_features[4193]  | ~\all_features[4192] )) | (\all_features[4196]  & (\all_features[4194]  | \all_features[4195] ));
  assign new_n22887_ = new_n19324_ & (new_n19333_ | new_n19322_ | (~new_n19328_ & ~new_n22888_ & ~new_n19332_));
  assign new_n22888_ = new_n22889_ & (~new_n22890_ | (~new_n22892_ & \all_features[4197]  & \all_features[4198]  & \all_features[4199] ));
  assign new_n22889_ = \all_features[4199]  & (\all_features[4198]  | (~new_n22884_ & \all_features[4197] ));
  assign new_n22890_ = \all_features[4199]  & \all_features[4198]  & ~new_n22891_ & new_n22885_;
  assign new_n22891_ = ~\all_features[4194]  & ~\all_features[4195]  & ~\all_features[4196]  & ~\all_features[4197]  & (~\all_features[4193]  | ~\all_features[4192] );
  assign new_n22892_ = ~\all_features[4195]  & ~\all_features[4196]  & (~\all_features[4194]  | new_n19331_);
  assign new_n22893_ = new_n19324_ & ~new_n19330_ & ~new_n22894_ & ~new_n19320_;
  assign new_n22894_ = ~new_n19328_ & ~new_n19322_ & ~new_n19332_ & ~new_n19333_ & (~new_n22890_ | ~new_n22889_);
  assign new_n22895_ = new_n22930_ ? ((new_n22931_ | ~new_n22897_ | ~new_n11549_) & (new_n22927_ | new_n11549_)) : new_n22896_;
  assign new_n22896_ = ~new_n8890_ & new_n7304_ & (new_n9867_ | new_n9834_);
  assign new_n22897_ = ~new_n22923_ & new_n22898_;
  assign new_n22898_ = ~new_n22899_ & ~new_n22922_;
  assign new_n22899_ = new_n22900_ & (~new_n22912_ | (new_n22909_ & new_n22920_));
  assign new_n22900_ = new_n22901_ & new_n22905_;
  assign new_n22901_ = ~new_n22902_ & (\all_features[3299]  | \all_features[3300]  | ~new_n22903_);
  assign new_n22902_ = new_n22903_ & ((~\all_features[3297]  & ~\all_features[3298]  & ~\all_features[3296] ) | ~\all_features[3300]  | ~\all_features[3299] );
  assign new_n22903_ = ~\all_features[3301]  & new_n22904_;
  assign new_n22904_ = ~\all_features[3302]  & ~\all_features[3303] ;
  assign new_n22905_ = ~new_n22906_ & ~new_n22908_;
  assign new_n22906_ = new_n22904_ & (~new_n22907_ | ~\all_features[3299]  | (~\all_features[3298]  & (~\all_features[3296]  | ~\all_features[3297] )));
  assign new_n22907_ = \all_features[3300]  & \all_features[3301] ;
  assign new_n22908_ = new_n22904_ & (~\all_features[3301]  | (~\all_features[3300]  & (~\all_features[3299]  | (~\all_features[3298]  & ~\all_features[3297] ))));
  assign new_n22909_ = \all_features[3303]  & \all_features[3302]  & ~new_n22911_ & new_n22910_;
  assign new_n22910_ = \all_features[3303]  & (\all_features[3302]  | (new_n22907_ & (\all_features[3298]  | \all_features[3299]  | \all_features[3297] )));
  assign new_n22911_ = ~\all_features[3298]  & ~\all_features[3299]  & ~\all_features[3300]  & ~\all_features[3301]  & (~\all_features[3297]  | ~\all_features[3296] );
  assign new_n22912_ = ~new_n22919_ & ~new_n22917_ & ~new_n22913_ & ~new_n22915_;
  assign new_n22913_ = ~new_n22914_ & ~\all_features[3303] ;
  assign new_n22914_ = \all_features[3301]  & \all_features[3302]  & (\all_features[3300]  | (\all_features[3298]  & \all_features[3299]  & \all_features[3297] ));
  assign new_n22915_ = ~\all_features[3303]  & (~\all_features[3299]  | ~new_n22907_ | ~new_n22916_ | ~\all_features[3298] );
  assign new_n22916_ = \all_features[3302]  & \all_features[3296]  & \all_features[3297] ;
  assign new_n22917_ = ~\all_features[3303]  & (~\all_features[3302]  | new_n22918_);
  assign new_n22918_ = ~\all_features[3301]  & (~\all_features[3299]  | ~\all_features[3300]  | ~\all_features[3298]  | (~\all_features[3297]  & ~\all_features[3296] ));
  assign new_n22919_ = ~\all_features[3303]  & (~\all_features[3302]  | (~\all_features[3301]  & ~\all_features[3300]  & (~\all_features[3299]  | ~\all_features[3298] )));
  assign new_n22920_ = \all_features[3303]  & (\all_features[3302]  | (~new_n22921_ & \all_features[3301] ));
  assign new_n22921_ = ~\all_features[3300]  & ~\all_features[3299]  & ~\all_features[3298]  & ~\all_features[3296]  & ~\all_features[3297] ;
  assign new_n22922_ = new_n22900_ & new_n22912_;
  assign new_n22923_ = new_n22901_ & (~new_n22905_ | (~new_n22924_ & ~new_n22917_ & ~new_n22919_));
  assign new_n22924_ = ~new_n22913_ & ~new_n22915_ & (~new_n22920_ | (~new_n22925_ & new_n22909_));
  assign new_n22925_ = \all_features[3303]  & \all_features[3302]  & ~new_n22926_ & \all_features[3301] ;
  assign new_n22926_ = ~\all_features[3299]  & ~\all_features[3300]  & (~\all_features[3298]  | (~\all_features[3297]  & ~\all_features[3296] ));
  assign new_n22927_ = new_n22928_ ? new_n8961_ : ~new_n15587_;
  assign new_n22928_ = ~new_n22929_ & new_n21241_;
  assign new_n22929_ = new_n21212_ & new_n21233_;
  assign new_n22930_ = new_n16337_ & (~new_n21998_ | ~new_n16338_);
  assign new_n22931_ = ~new_n22932_ & (~new_n22934_ | new_n22933_);
  assign new_n22932_ = new_n22176_ & new_n22179_;
  assign new_n22933_ = ~new_n22146_ & ~new_n22167_;
  assign new_n22934_ = ~new_n22176_ & new_n22179_;
  assign new_n22935_ = new_n15751_ ? (new_n12303_ ? new_n22936_ : new_n22938_) : new_n22942_;
  assign new_n22936_ = new_n22937_ ? ~new_n20578_ : new_n16103_;
  assign new_n22937_ = ~new_n14600_ & new_n16755_;
  assign new_n22938_ = (~new_n22939_ & new_n22941_) | (~new_n22500_ & ~new_n22941_ & (~new_n22498_ | new_n22466_));
  assign new_n22939_ = ~new_n21245_ & new_n22940_;
  assign new_n22940_ = ~new_n21233_ & ~new_n21242_;
  assign new_n22941_ = new_n22361_ & (~new_n12984_ | ~new_n22356_);
  assign new_n22942_ = new_n22386_ & (new_n19829_ | new_n13923_);
  assign new_n22943_ = new_n22944_ ? (new_n22953_ ^ new_n22991_) : (~new_n22953_ ^ new_n22991_);
  assign new_n22944_ = ~new_n22951_ & new_n22945_;
  assign new_n22945_ = (new_n22950_ | ~new_n13773_ | ~new_n22948_) & (new_n22948_ | (new_n22946_ & (~new_n20088_ | new_n22457_)));
  assign new_n22946_ = (~new_n22947_ | new_n10490_ | new_n20088_) & (new_n16571_ | ~new_n22457_ | ~new_n13921_ | ~new_n20088_);
  assign new_n22947_ = ~new_n7980_ & new_n14847_;
  assign new_n22948_ = new_n22949_ & new_n8854_;
  assign new_n22949_ = new_n8841_ & new_n8851_;
  assign new_n22950_ = (~new_n14337_ & ~new_n7327_) | (new_n14723_ & new_n7327_ & (new_n14720_ | new_n14692_));
  assign new_n22951_ = ~new_n13773_ & ~new_n10129_ & new_n22948_ & (~new_n7063_ | (~new_n7041_ & new_n22952_));
  assign new_n22952_ = ~new_n11629_ & ~new_n19049_;
  assign new_n22953_ = ~new_n22954_ & new_n22990_;
  assign new_n22954_ = ~new_n22955_ | (new_n22987_ & (new_n15671_ | ~new_n13887_ | ~new_n21430_) & (new_n22989_ | new_n21430_));
  assign new_n22955_ = ~new_n22986_ & (~new_n22982_ | ~new_n22956_);
  assign new_n22956_ = ~new_n22957_ & (\all_features[5971]  | \all_features[5972]  | \all_features[5973]  | \all_features[5974]  | \all_features[5975] );
  assign new_n22957_ = new_n22958_ & (new_n22979_ | (~new_n22977_ & (new_n22969_ | (~new_n22980_ & ~new_n22971_))));
  assign new_n22958_ = ~new_n22974_ & ~new_n22978_ & ~new_n22976_ & (new_n22979_ | new_n22977_ | new_n22959_);
  assign new_n22959_ = ~new_n22971_ & ~new_n22969_ & (~new_n22960_ | (~new_n22973_ & new_n22964_));
  assign new_n22960_ = \all_features[5975]  & (\all_features[5974]  | (~new_n22961_ & \all_features[5973] ));
  assign new_n22961_ = new_n22962_ & ~\all_features[5972]  & new_n22963_;
  assign new_n22962_ = ~\all_features[5968]  & ~\all_features[5969] ;
  assign new_n22963_ = ~\all_features[5970]  & ~\all_features[5971] ;
  assign new_n22964_ = new_n22965_ & new_n22968_ & (new_n22967_ | \all_features[5972]  | \all_features[5973]  | ~new_n22963_);
  assign new_n22965_ = \all_features[5975]  & (\all_features[5974]  | (new_n22966_ & (\all_features[5970]  | \all_features[5971]  | \all_features[5969] )));
  assign new_n22966_ = \all_features[5972]  & \all_features[5973] ;
  assign new_n22967_ = \all_features[5968]  & \all_features[5969] ;
  assign new_n22968_ = \all_features[5974]  & \all_features[5975] ;
  assign new_n22969_ = ~new_n22970_ & ~\all_features[5975] ;
  assign new_n22970_ = \all_features[5973]  & \all_features[5974]  & (\all_features[5972]  | (\all_features[5970]  & \all_features[5971]  & \all_features[5969] ));
  assign new_n22971_ = ~\all_features[5975]  & (~\all_features[5974]  | ~new_n22972_ | ~new_n22967_ | ~new_n22966_);
  assign new_n22972_ = \all_features[5970]  & \all_features[5971] ;
  assign new_n22973_ = new_n22968_ & \all_features[5973]  & ((~new_n22962_ & \all_features[5970] ) | \all_features[5972]  | \all_features[5971] );
  assign new_n22974_ = new_n22975_ & (~\all_features[5973]  | (~\all_features[5972]  & (~\all_features[5971]  | (~\all_features[5970]  & ~\all_features[5969] ))));
  assign new_n22975_ = ~\all_features[5974]  & ~\all_features[5975] ;
  assign new_n22976_ = ~\all_features[5973]  & new_n22975_ & ((~\all_features[5970]  & new_n22962_) | ~\all_features[5972]  | ~\all_features[5971] );
  assign new_n22977_ = ~\all_features[5975]  & (~\all_features[5974]  | (~\all_features[5973]  & (new_n22962_ | ~new_n22972_ | ~\all_features[5972] )));
  assign new_n22978_ = new_n22975_ & (~\all_features[5971]  | ~new_n22966_ | (~\all_features[5970]  & ~new_n22967_));
  assign new_n22979_ = ~\all_features[5975]  & (~\all_features[5974]  | (~\all_features[5972]  & ~\all_features[5973]  & ~new_n22972_));
  assign new_n22980_ = \all_features[5975]  & ((new_n22981_ & (\all_features[5974]  | \all_features[5973] )) | (~\all_features[5974]  & (\all_features[5973]  ? new_n22961_ : \all_features[5972] )));
  assign new_n22981_ = new_n22965_ & (\all_features[5973]  | ~new_n22968_ | (~new_n22967_ & ~\all_features[5972]  & new_n22963_) | (\all_features[5972]  & ~new_n22963_));
  assign new_n22982_ = new_n22985_ & ~new_n22978_ & ~new_n22983_ & ~new_n22974_;
  assign new_n22983_ = ~new_n22969_ & ~new_n22977_ & new_n22984_ & (~new_n22964_ | ~new_n22960_);
  assign new_n22984_ = ~new_n22971_ & ~new_n22979_;
  assign new_n22985_ = ~new_n22976_ & (\all_features[5971]  | \all_features[5972]  | \all_features[5973]  | \all_features[5974]  | \all_features[5975] );
  assign new_n22986_ = new_n22984_ & new_n22985_ & ~new_n22978_ & ~new_n22977_ & ~new_n22969_ & ~new_n22974_;
  assign new_n22987_ = (new_n22988_ | ~new_n15671_ | ~new_n21430_) & (new_n8030_ | new_n6591_ | new_n21430_);
  assign new_n22988_ = new_n9275_ & (new_n9249_ | ~new_n14385_);
  assign new_n22989_ = new_n8030_ ? ~new_n17936_ : ~new_n6591_;
  assign new_n22990_ = new_n22955_ & (new_n17936_ | ~new_n8030_ | new_n21430_) & (new_n15671_ | new_n13887_ | ~new_n21430_);
  assign new_n22991_ = new_n22996_ & (new_n15018_ | new_n16957_ | new_n6639_ | new_n22997_) & (new_n22992_ | ~new_n22997_);
  assign new_n22992_ = ~new_n22993_ & ((~new_n9654_ & ~new_n9686_) | new_n12798_ | new_n22995_);
  assign new_n22993_ = ~new_n19501_ & new_n12798_ & new_n11468_ & (new_n11446_ | new_n22994_);
  assign new_n22994_ = new_n15153_ & new_n15157_;
  assign new_n22995_ = new_n8320_ & new_n10775_;
  assign new_n22996_ = (~new_n22995_ | new_n12798_ | ~new_n22997_) & (new_n22998_ | ~new_n16957_ | ~new_n15751_ | new_n22997_);
  assign new_n22997_ = new_n13135_ & (~new_n13164_ | ~new_n13160_);
  assign new_n22998_ = new_n20959_ & new_n21618_;
  assign new_n22999_ = ~new_n23000_ & new_n22955_;
  assign new_n23000_ = new_n23033_ ? new_n23001_ : ((new_n20337_ | ~new_n20587_ | ~new_n23034_) & (~new_n14469_ | new_n23034_));
  assign new_n23001_ = (new_n23002_ | ~new_n23032_) & (new_n10204_ | (new_n10201_ & new_n13097_));
  assign new_n23002_ = ~new_n23003_ & ~new_n23025_;
  assign new_n23003_ = new_n23020_ & ~new_n23024_ & ~new_n23004_ & ~new_n23023_;
  assign new_n23004_ = new_n23005_ & (~new_n23018_ | ~new_n23019_ | ~new_n23015_ | ~new_n23017_);
  assign new_n23005_ = ~new_n23014_ & ~new_n23011_ & ~new_n23006_ & ~new_n23009_;
  assign new_n23006_ = ~\all_features[2623]  & (~\all_features[2622]  | (~\all_features[2621]  & (new_n23007_ | ~new_n23008_ | ~\all_features[2620] )));
  assign new_n23007_ = ~\all_features[2616]  & ~\all_features[2617] ;
  assign new_n23008_ = \all_features[2618]  & \all_features[2619] ;
  assign new_n23009_ = ~new_n23010_ & ~\all_features[2623] ;
  assign new_n23010_ = \all_features[2621]  & \all_features[2622]  & (\all_features[2620]  | (\all_features[2618]  & \all_features[2619]  & \all_features[2617] ));
  assign new_n23011_ = ~\all_features[2623]  & (~\all_features[2622]  | ~new_n23012_ | ~new_n23013_ | ~new_n23008_);
  assign new_n23012_ = \all_features[2620]  & \all_features[2621] ;
  assign new_n23013_ = \all_features[2616]  & \all_features[2617] ;
  assign new_n23014_ = ~\all_features[2623]  & (~\all_features[2622]  | (~\all_features[2620]  & ~\all_features[2621]  & ~new_n23008_));
  assign new_n23015_ = \all_features[2623]  & (\all_features[2622]  | (\all_features[2621]  & (\all_features[2620]  | ~new_n23007_ | ~new_n23016_)));
  assign new_n23016_ = ~\all_features[2618]  & ~\all_features[2619] ;
  assign new_n23017_ = \all_features[2623]  & (\all_features[2622]  | (new_n23012_ & (\all_features[2618]  | \all_features[2619]  | \all_features[2617] )));
  assign new_n23018_ = \all_features[2622]  & \all_features[2623]  & (\all_features[2620]  | \all_features[2621]  | new_n23013_ | ~new_n23016_);
  assign new_n23019_ = \all_features[2623]  & (\all_features[2621]  | \all_features[2622]  | \all_features[2620] );
  assign new_n23020_ = ~new_n23021_ & (\all_features[2619]  | \all_features[2620]  | \all_features[2621]  | \all_features[2622]  | \all_features[2623] );
  assign new_n23021_ = ~\all_features[2621]  & new_n23022_ & ((~\all_features[2618]  & new_n23007_) | ~\all_features[2620]  | ~\all_features[2619] );
  assign new_n23022_ = ~\all_features[2622]  & ~\all_features[2623] ;
  assign new_n23023_ = new_n23022_ & (~\all_features[2621]  | (~\all_features[2620]  & (~\all_features[2619]  | (~\all_features[2618]  & ~\all_features[2617] ))));
  assign new_n23024_ = new_n23022_ & (~\all_features[2619]  | ~new_n23012_ | (~\all_features[2618]  & ~new_n23013_));
  assign new_n23025_ = new_n23020_ & (~new_n23031_ | (~new_n23026_ & new_n23030_));
  assign new_n23026_ = new_n23029_ & ((~new_n23027_ & new_n23017_ & new_n23018_) | ~new_n23019_ | ~new_n23015_);
  assign new_n23027_ = \all_features[2623]  & \all_features[2622]  & ~new_n23028_ & \all_features[2621] ;
  assign new_n23028_ = ~\all_features[2619]  & ~\all_features[2620]  & (~\all_features[2618]  | new_n23007_);
  assign new_n23029_ = ~new_n23009_ & ~new_n23011_;
  assign new_n23030_ = ~new_n23006_ & ~new_n23014_;
  assign new_n23031_ = ~new_n23023_ & ~new_n23024_;
  assign new_n23032_ = new_n23031_ & new_n23030_ & new_n23020_ & new_n23029_;
  assign new_n23033_ = new_n11550_ & new_n12851_;
  assign new_n23034_ = ~new_n23035_ & ~new_n23058_;
  assign new_n23035_ = new_n23053_ & ~new_n23057_ & ~new_n23036_ & ~new_n23056_;
  assign new_n23036_ = ~new_n23051_ & ~new_n23052_ & new_n23044_ & (~new_n23049_ | ~new_n23037_);
  assign new_n23037_ = new_n23043_ & new_n23038_ & new_n23040_;
  assign new_n23038_ = \all_features[2295]  & (\all_features[2294]  | (new_n23039_ & (\all_features[2290]  | \all_features[2291]  | \all_features[2289] )));
  assign new_n23039_ = \all_features[2292]  & \all_features[2293] ;
  assign new_n23040_ = \all_features[2294]  & \all_features[2295]  & (\all_features[2292]  | \all_features[2293]  | new_n23042_ | ~new_n23041_);
  assign new_n23041_ = ~\all_features[2290]  & ~\all_features[2291] ;
  assign new_n23042_ = \all_features[2288]  & \all_features[2289] ;
  assign new_n23043_ = \all_features[2295]  & (\all_features[2293]  | \all_features[2294]  | \all_features[2292] );
  assign new_n23044_ = ~new_n23045_ & ~new_n23047_;
  assign new_n23045_ = ~new_n23046_ & ~\all_features[2295] ;
  assign new_n23046_ = \all_features[2293]  & \all_features[2294]  & (\all_features[2292]  | (\all_features[2290]  & \all_features[2291]  & \all_features[2289] ));
  assign new_n23047_ = ~\all_features[2295]  & (~\all_features[2294]  | (~\all_features[2292]  & ~\all_features[2293]  & ~new_n23048_));
  assign new_n23048_ = \all_features[2290]  & \all_features[2291] ;
  assign new_n23049_ = \all_features[2295]  & (\all_features[2294]  | (\all_features[2293]  & (\all_features[2292]  | ~new_n23050_ | ~new_n23041_)));
  assign new_n23050_ = ~\all_features[2288]  & ~\all_features[2289] ;
  assign new_n23051_ = ~\all_features[2295]  & (~\all_features[2294]  | (~\all_features[2293]  & (new_n23050_ | ~new_n23048_ | ~\all_features[2292] )));
  assign new_n23052_ = ~\all_features[2295]  & (~\all_features[2294]  | ~new_n23039_ | ~new_n23042_ | ~new_n23048_);
  assign new_n23053_ = ~new_n23054_ & (\all_features[2291]  | \all_features[2292]  | \all_features[2293]  | \all_features[2294]  | \all_features[2295] );
  assign new_n23054_ = ~\all_features[2293]  & new_n23055_ & ((~\all_features[2290]  & new_n23050_) | ~\all_features[2292]  | ~\all_features[2291] );
  assign new_n23055_ = ~\all_features[2294]  & ~\all_features[2295] ;
  assign new_n23056_ = new_n23055_ & (~\all_features[2293]  | (~\all_features[2292]  & (~\all_features[2291]  | (~\all_features[2290]  & ~\all_features[2289] ))));
  assign new_n23057_ = new_n23055_ & (~\all_features[2291]  | ~new_n23039_ | (~\all_features[2290]  & ~new_n23042_));
  assign new_n23058_ = new_n23053_ & new_n23044_ & new_n23059_ & ~new_n23051_ & ~new_n23052_;
  assign new_n23059_ = ~new_n23056_ & ~new_n23057_;
  assign new_n23060_ = new_n23066_ & (new_n21208_ | new_n23061_);
  assign new_n23061_ = (new_n23064_ | ~new_n23062_ | ~new_n16957_) & (new_n16957_ | (new_n19057_ ? new_n16762_ : ~new_n23065_));
  assign new_n23062_ = new_n7866_ & (new_n7863_ | ~new_n23063_);
  assign new_n23063_ = ~new_n7835_ & ~new_n7859_;
  assign new_n23064_ = ~new_n16482_ & new_n19432_;
  assign new_n23065_ = new_n19677_ & new_n21401_ & new_n19651_;
  assign new_n23066_ = (~new_n23069_ | new_n23068_) & (new_n23062_ | ~new_n16957_ | new_n21208_) & (new_n23067_ | ~new_n23068_ | ~new_n21208_);
  assign new_n23067_ = (new_n19717_ & new_n12338_ & new_n12753_) | (new_n9275_ & (new_n12529_ | new_n9249_) & (~new_n12338_ | ~new_n12753_));
  assign new_n23068_ = ~new_n6591_ | (~new_n6569_ & ~new_n6592_);
  assign new_n23069_ = new_n23072_ & new_n21208_ & new_n23071_ & (new_n13055_ | new_n10438_ | ~new_n23070_);
  assign new_n23070_ = ~new_n13057_ & ~new_n13041_;
  assign new_n23071_ = new_n10434_ & new_n19823_;
  assign new_n23072_ = new_n10409_ & new_n10432_;
  assign new_n23073_ = new_n23076_ & ((new_n23080_ & (new_n18633_ | new_n8097_)) | new_n18579_ | (new_n23074_ & ~new_n18633_ & ~new_n8097_));
  assign new_n23074_ = (new_n15588_ & new_n7408_) | (~new_n15904_ & ~new_n15906_ & new_n23075_ & ~new_n7408_);
  assign new_n23075_ = ~new_n15875_ & ~new_n15895_;
  assign new_n23076_ = (~new_n23077_ | new_n16762_ | new_n20168_) & (new_n23079_ | ~new_n10701_ | ~new_n18579_ | ~new_n20168_);
  assign new_n23077_ = new_n20205_ & ~new_n23078_ & new_n18579_;
  assign new_n23078_ = ~new_n20194_ & ~new_n20202_;
  assign new_n23079_ = ~new_n7991_ & (~new_n7988_ | ~new_n7980_);
  assign new_n23080_ = ~new_n19457_ & (~new_n7103_ | ~new_n23081_) & (~new_n19435_ | ~new_n20785_);
  assign new_n23081_ = new_n7128_ & new_n7131_;
  assign new_n23082_ = ~new_n23083_ & ~new_n23125_;
  assign new_n23083_ = new_n23085_ & (new_n22897_ | ~new_n23087_ | (new_n23122_ ? new_n23123_ : new_n23084_));
  assign new_n23084_ = new_n6388_ & (new_n6385_ | ~new_n6355_);
  assign new_n23085_ = new_n23086_ & (~new_n23087_ | ~new_n22897_ | (~new_n19591_ & ~new_n23121_ & new_n14351_));
  assign new_n23086_ = new_n23087_ | ((new_n23088_ | new_n12447_ | ~new_n22287_) & (new_n18459_ | new_n22287_));
  assign new_n23087_ = new_n7097_ & new_n10609_;
  assign new_n23088_ = ~new_n23089_ & new_n23117_;
  assign new_n23089_ = ~new_n23116_ & (new_n23109_ | new_n23112_ | new_n23114_ | new_n23115_ | new_n23090_);
  assign new_n23090_ = ~new_n23103_ & ~new_n23108_ & ((~new_n23091_ & new_n23100_) | new_n23107_ | new_n23105_);
  assign new_n23091_ = new_n23092_ & (new_n23098_ | ~\all_features[773]  | ~\all_features[774]  | ~\all_features[775] );
  assign new_n23092_ = \all_features[775]  & \all_features[774]  & ~new_n23093_ & new_n23096_;
  assign new_n23093_ = new_n23094_ & ~\all_features[773]  & ~new_n23095_ & ~\all_features[772] ;
  assign new_n23094_ = ~\all_features[770]  & ~\all_features[771] ;
  assign new_n23095_ = \all_features[768]  & \all_features[769] ;
  assign new_n23096_ = \all_features[775]  & (\all_features[774]  | (new_n23097_ & (\all_features[770]  | \all_features[771]  | \all_features[769] )));
  assign new_n23097_ = \all_features[772]  & \all_features[773] ;
  assign new_n23098_ = ~\all_features[771]  & ~\all_features[772]  & (~\all_features[770]  | new_n23099_);
  assign new_n23099_ = ~\all_features[768]  & ~\all_features[769] ;
  assign new_n23100_ = new_n23101_ & new_n23102_;
  assign new_n23101_ = \all_features[775]  & (\all_features[774]  | (\all_features[773]  & (\all_features[772]  | ~new_n23099_ | ~new_n23094_)));
  assign new_n23102_ = \all_features[775]  & (\all_features[773]  | \all_features[774]  | \all_features[772] );
  assign new_n23103_ = ~\all_features[775]  & (~\all_features[774]  | (~\all_features[773]  & (new_n23099_ | ~new_n23104_ | ~\all_features[772] )));
  assign new_n23104_ = \all_features[770]  & \all_features[771] ;
  assign new_n23105_ = ~new_n23106_ & ~\all_features[775] ;
  assign new_n23106_ = \all_features[773]  & \all_features[774]  & (\all_features[772]  | (\all_features[770]  & \all_features[771]  & \all_features[769] ));
  assign new_n23107_ = ~\all_features[775]  & (~\all_features[774]  | ~new_n23095_ | ~new_n23097_ | ~new_n23104_);
  assign new_n23108_ = ~\all_features[775]  & (~\all_features[774]  | (~\all_features[772]  & ~\all_features[773]  & ~new_n23104_));
  assign new_n23109_ = ~new_n23108_ & (new_n23103_ | (~new_n23105_ & (new_n23107_ | new_n23110_)));
  assign new_n23110_ = new_n23102_ & (~new_n23101_ | (~new_n23111_ & new_n23096_));
  assign new_n23111_ = ~\all_features[773]  & \all_features[774]  & \all_features[775]  & (\all_features[772]  ? new_n23094_ : (new_n23095_ | ~new_n23094_));
  assign new_n23112_ = new_n23113_ & (~\all_features[773]  | (~\all_features[772]  & (~\all_features[771]  | (~\all_features[770]  & ~\all_features[769] ))));
  assign new_n23113_ = ~\all_features[774]  & ~\all_features[775] ;
  assign new_n23114_ = new_n23113_ & (~\all_features[771]  | ~new_n23097_ | (~\all_features[770]  & ~new_n23095_));
  assign new_n23115_ = ~\all_features[773]  & new_n23113_ & ((~\all_features[770]  & new_n23099_) | ~\all_features[772]  | ~\all_features[771] );
  assign new_n23116_ = ~\all_features[775]  & ~\all_features[774]  & ~\all_features[773]  & ~\all_features[771]  & ~\all_features[772] ;
  assign new_n23117_ = new_n23112_ | ~new_n23119_ | ((new_n23105_ | ~new_n23120_) & (new_n23118_ | new_n23114_));
  assign new_n23118_ = ~new_n23103_ & ~new_n23105_ & ~new_n23107_ & ~new_n23108_ & (~new_n23100_ | ~new_n23092_);
  assign new_n23119_ = ~new_n23115_ & ~new_n23116_;
  assign new_n23120_ = ~new_n23114_ & ~new_n23108_ & ~new_n23103_ & ~new_n23107_;
  assign new_n23121_ = ~new_n6883_ & (~new_n6880_ | ~new_n6869_);
  assign new_n23122_ = ~new_n10682_ & (~new_n13924_ | new_n13932_);
  assign new_n23123_ = new_n6770_ & new_n23124_;
  assign new_n23124_ = ~new_n6799_ & ~new_n6801_;
  assign new_n23125_ = new_n18459_ & ~new_n23087_ & ~new_n22287_;
  assign new_n23126_ = new_n23127_ ? (new_n23143_ ^ new_n23154_) : (~new_n23143_ ^ new_n23154_);
  assign new_n23127_ = ~new_n23128_ & new_n23141_;
  assign new_n23128_ = new_n23129_ & (new_n16263_ | (~new_n20971_ & new_n7408_ & new_n23064_) | (new_n23138_ & ~new_n23064_));
  assign new_n23129_ = ~new_n16263_ | ((new_n23130_ | (new_n23131_ & (new_n23137_ | new_n23135_))) & (new_n23136_ | ~new_n23131_ | ~new_n23135_));
  assign new_n23130_ = ~new_n23131_ & ~new_n23133_ & (new_n17444_ | (new_n17416_ & new_n17437_ & new_n17446_));
  assign new_n23131_ = new_n23132_ & new_n12398_;
  assign new_n23132_ = new_n12376_ & new_n12404_;
  assign new_n23133_ = new_n23134_ & ~new_n17353_ & ~new_n22438_;
  assign new_n23134_ = ~new_n17330_ & ~new_n17357_;
  assign new_n23135_ = new_n18102_ & new_n11884_;
  assign new_n23136_ = new_n10871_ & (new_n10868_ | ~new_n10839_);
  assign new_n23137_ = ~new_n7221_ & (~new_n7218_ | ~new_n7194_);
  assign new_n23138_ = new_n23139_ ? new_n23140_ : ~new_n22546_;
  assign new_n23139_ = ~new_n8188_ & (~new_n8166_ | ~new_n8191_);
  assign new_n23140_ = ~new_n17886_ & ~new_n17888_;
  assign new_n23141_ = new_n16263_ ? new_n23142_ : ((new_n20971_ | ~new_n7408_ | ~new_n23064_) & (~new_n23138_ | new_n23064_));
  assign new_n23142_ = ~new_n23130_ & (~new_n23131_ | ~new_n23135_ | ~new_n23136_);
  assign new_n23143_ = ~new_n23151_ & new_n23144_;
  assign new_n23144_ = new_n23145_ & (~new_n22897_ | ~new_n14388_ | (new_n21641_ ? new_n23150_ : ~new_n23149_));
  assign new_n23145_ = (new_n14388_ | new_n23146_ | ~new_n22897_) & (new_n6701_ | new_n22036_ | ~new_n23148_ | new_n22897_);
  assign new_n23146_ = new_n13038_ & new_n23133_ & new_n23147_;
  assign new_n23147_ = new_n13015_ & new_n14339_;
  assign new_n23148_ = new_n20342_ & ~new_n20371_ & ~new_n20406_;
  assign new_n23149_ = new_n22633_ & (new_n22611_ | ~new_n22634_);
  assign new_n23150_ = ~new_n14091_ & new_n17804_;
  assign new_n23151_ = ~new_n22897_ & ((~new_n23152_ & new_n6701_) | (~new_n23148_ & ~new_n12305_ & new_n21685_ & ~new_n6701_));
  assign new_n23152_ = (~new_n19547_ | new_n19280_) & (~new_n9234_ | (~new_n9211_ & ~new_n23153_));
  assign new_n23153_ = new_n9237_ & new_n9241_;
  assign new_n23154_ = new_n23157_ & (new_n23161_ ? ~new_n23163_ : (new_n10936_ | new_n23155_));
  assign new_n23155_ = new_n21615_ ? (~new_n14845_ | (~new_n23156_ & ~new_n14843_)) : new_n22386_;
  assign new_n23156_ = new_n14814_ & new_n14834_;
  assign new_n23157_ = ~new_n10936_ | ((new_n23159_ | new_n23158_ | ~new_n23160_) & (new_n8590_ | ~new_n19147_ | new_n23160_));
  assign new_n23158_ = new_n9867_ & ~new_n15531_ & new_n15914_;
  assign new_n23159_ = new_n12598_ & ~new_n8357_ & new_n15531_;
  assign new_n23160_ = new_n13503_ & (new_n13506_ | new_n13480_);
  assign new_n23161_ = new_n22872_ & (new_n22874_ | ~new_n23162_);
  assign new_n23162_ = ~new_n22842_ & ~new_n22863_;
  assign new_n23163_ = new_n23164_ & (~new_n13369_ | new_n13392_);
  assign new_n23164_ = ~new_n13391_ & ~new_n10936_ & (new_n13921_ | (new_n13909_ & new_n13918_));
  assign new_n23165_ = ~new_n23166_ & new_n23176_;
  assign new_n23166_ = new_n23171_ & (~new_n10773_ | ((~new_n15588_ | ~new_n23175_ | new_n18579_) & (new_n23167_ | ~new_n18579_)));
  assign new_n23167_ = new_n23168_ ? ~new_n23169_ : new_n20171_;
  assign new_n23168_ = new_n8097_ & (new_n8094_ | new_n8061_);
  assign new_n23169_ = new_n23170_ & new_n13838_;
  assign new_n23170_ = new_n13830_ & new_n13840_;
  assign new_n23171_ = new_n10773_ | (new_n10701_ ? new_n23172_ : new_n23173_);
  assign new_n23172_ = new_n17675_ ? ~new_n13523_ : ~new_n22461_;
  assign new_n23173_ = ~new_n13516_ & new_n23174_;
  assign new_n23174_ = new_n23063_ & new_n12756_;
  assign new_n23175_ = ~new_n18941_ & new_n22702_;
  assign new_n23176_ = new_n23177_ & (~new_n10773_ | ((new_n23180_ | ~new_n18579_) & (new_n23175_ | ~new_n15588_ | new_n18579_)));
  assign new_n23177_ = (new_n18579_ | ~new_n23178_ | ~new_n10773_) & (new_n10773_ | (new_n10701_ ? ~new_n23172_ : ~new_n23173_));
  assign new_n23178_ = ~new_n15588_ & new_n23179_;
  assign new_n23179_ = ~new_n9093_ & ~new_n9097_;
  assign new_n23180_ = new_n23168_ ? new_n23169_ : ~new_n20171_;
  assign new_n23181_ = ~new_n23191_ & (new_n23192_ | (new_n23182_ & (new_n23189_ | ~new_n23133_ | ~new_n23195_)));
  assign new_n23182_ = new_n23133_ ? (~new_n23189_ | (new_n16228_ & new_n23190_)) : new_n23183_;
  assign new_n23183_ = new_n15549_ ? new_n23188_ : ~new_n23184_;
  assign new_n23184_ = new_n19604_ & (new_n19626_ | (~new_n23185_ & ~new_n19624_));
  assign new_n23185_ = ~new_n19629_ & (new_n19628_ | (~new_n19622_ & (new_n19608_ | (~new_n19620_ & ~new_n23186_))));
  assign new_n23186_ = ~new_n19619_ & (~new_n19618_ | (new_n19617_ & (~new_n19612_ | (~new_n23187_ & new_n19614_))));
  assign new_n23187_ = \all_features[5742]  & \all_features[5743]  & (\all_features[5741]  | (~new_n19615_ & \all_features[5740] ));
  assign new_n23188_ = new_n15675_ & new_n17849_;
  assign new_n23189_ = new_n12980_ & (new_n12978_ | ~new_n14045_);
  assign new_n23190_ = new_n8772_ & new_n8768_;
  assign new_n23191_ = ~new_n14350_ & new_n23192_ & (new_n23194_ ? ~new_n11575_ : ~new_n12152_);
  assign new_n23192_ = new_n23193_ & new_n10024_;
  assign new_n23193_ = new_n10002_ & new_n10032_;
  assign new_n23194_ = ~new_n12187_ & (~new_n12185_ | ~new_n12175_);
  assign new_n23195_ = new_n10607_ & (new_n10604_ | ~new_n23196_);
  assign new_n23196_ = ~new_n10575_ & ~new_n10596_;
  assign new_n23197_ = new_n23198_ & (new_n15152_ | new_n23241_ | new_n15786_);
  assign new_n23198_ = ~new_n23216_ & (new_n23218_ ? ~new_n23219_ : (~new_n23199_ | (~new_n23221_ & new_n23239_)));
  assign new_n23199_ = new_n16362_ & ~new_n23200_ & new_n15786_;
  assign new_n23200_ = new_n23201_ & ~new_n23215_ & ~new_n23214_ & ~new_n23211_ & ~new_n23213_;
  assign new_n23201_ = ~new_n23210_ & ~new_n23209_ & ~new_n23202_ & ~new_n23205_;
  assign new_n23202_ = ~\all_features[1975]  & (~\all_features[1974]  | (~\all_features[1973]  & (new_n23204_ | ~\all_features[1972]  | ~new_n23203_)));
  assign new_n23203_ = \all_features[1970]  & \all_features[1971] ;
  assign new_n23204_ = ~\all_features[1968]  & ~\all_features[1969] ;
  assign new_n23205_ = new_n23206_ & (~\all_features[1971]  | ~new_n23208_ | (~\all_features[1970]  & ~new_n23207_));
  assign new_n23206_ = ~\all_features[1974]  & ~\all_features[1975] ;
  assign new_n23207_ = \all_features[1968]  & \all_features[1969] ;
  assign new_n23208_ = \all_features[1972]  & \all_features[1973] ;
  assign new_n23209_ = ~\all_features[1973]  & new_n23206_ & ((~\all_features[1970]  & new_n23204_) | ~\all_features[1972]  | ~\all_features[1971] );
  assign new_n23210_ = ~\all_features[1975]  & (~\all_features[1974]  | (~\all_features[1972]  & ~\all_features[1973]  & ~new_n23203_));
  assign new_n23211_ = ~new_n23212_ & ~\all_features[1975] ;
  assign new_n23212_ = \all_features[1973]  & \all_features[1974]  & (\all_features[1972]  | (\all_features[1970]  & \all_features[1971]  & \all_features[1969] ));
  assign new_n23213_ = new_n23206_ & (~\all_features[1973]  | (~\all_features[1972]  & (~\all_features[1971]  | (~\all_features[1970]  & ~\all_features[1969] ))));
  assign new_n23214_ = ~\all_features[1975]  & (~\all_features[1974]  | ~new_n23207_ | ~new_n23208_ | ~new_n23203_);
  assign new_n23215_ = ~\all_features[1975]  & ~\all_features[1974]  & ~\all_features[1973]  & ~\all_features[1971]  & ~\all_features[1972] ;
  assign new_n23216_ = new_n15152_ & new_n23217_ & ~new_n19717_ & ~new_n15786_;
  assign new_n23217_ = ~new_n22467_ & new_n22546_;
  assign new_n23218_ = new_n14294_ & (~new_n14325_ | ~new_n14321_);
  assign new_n23219_ = ~new_n8161_ & new_n23220_ & new_n15786_ & (new_n21357_ | new_n21387_);
  assign new_n23220_ = ~new_n8134_ & ~new_n8159_;
  assign new_n23221_ = ~new_n23222_ & (new_n23215_ | (~new_n23209_ & (new_n23213_ | new_n23235_)));
  assign new_n23222_ = new_n23233_ & (~new_n23234_ | (new_n23231_ & (~new_n23232_ | new_n23223_)));
  assign new_n23223_ = new_n23230_ & ~new_n23226_ & new_n23224_;
  assign new_n23224_ = \all_features[1975]  & (\all_features[1974]  | new_n23225_);
  assign new_n23225_ = \all_features[1973]  & (\all_features[1970]  | \all_features[1971]  | \all_features[1972]  | ~new_n23204_);
  assign new_n23226_ = ~new_n23228_ & new_n23227_ & \all_features[1974]  & \all_features[1975]  & (~\all_features[1973]  | new_n23229_);
  assign new_n23227_ = \all_features[1975]  & (\all_features[1974]  | (new_n23208_ & (\all_features[1970]  | \all_features[1971]  | \all_features[1969] )));
  assign new_n23228_ = ~\all_features[1973]  & ~\all_features[1972]  & ~\all_features[1971]  & ~new_n23207_ & ~\all_features[1970] ;
  assign new_n23229_ = ~\all_features[1971]  & ~\all_features[1972]  & (~\all_features[1970]  | new_n23204_);
  assign new_n23230_ = \all_features[1975]  & (\all_features[1973]  | \all_features[1974]  | \all_features[1972] );
  assign new_n23231_ = ~new_n23202_ & ~new_n23210_;
  assign new_n23232_ = ~new_n23211_ & ~new_n23214_;
  assign new_n23233_ = ~new_n23209_ & ~new_n23215_;
  assign new_n23234_ = ~new_n23213_ & ~new_n23205_;
  assign new_n23235_ = ~new_n23205_ & (new_n23210_ | (~new_n23202_ & (new_n23211_ | (~new_n23214_ & ~new_n23236_))));
  assign new_n23236_ = new_n23230_ & (~new_n23224_ | (new_n23227_ & (new_n23238_ | ~new_n23237_)));
  assign new_n23237_ = \all_features[1975]  & ~new_n23228_ & \all_features[1974] ;
  assign new_n23238_ = \all_features[1974]  & \all_features[1975]  & (\all_features[1973]  | (\all_features[1972]  & (\all_features[1971]  | \all_features[1970] )));
  assign new_n23239_ = new_n23233_ & new_n23234_ & (~new_n23232_ | ~new_n23231_ | (new_n23240_ & new_n23224_));
  assign new_n23240_ = new_n23230_ & new_n23237_ & new_n23227_;
  assign new_n23241_ = (~new_n21769_ & new_n19231_) ? new_n13349_ : ~new_n23242_;
  assign new_n23242_ = ~new_n23271_ & (~new_n23264_ | ~new_n23243_ | ~new_n23273_);
  assign new_n23243_ = ~new_n23244_ & (\all_features[1539]  | \all_features[1540]  | \all_features[1541]  | \all_features[1542]  | \all_features[1543] );
  assign new_n23244_ = ~new_n23260_ & (new_n23258_ | (~new_n23262_ & (new_n23263_ | (~new_n23261_ & ~new_n23245_))));
  assign new_n23245_ = ~new_n23246_ & (new_n23248_ | (new_n23257_ & (~new_n23252_ | (~new_n23256_ & new_n23255_))));
  assign new_n23246_ = ~new_n23247_ & ~\all_features[1543] ;
  assign new_n23247_ = \all_features[1541]  & \all_features[1542]  & (\all_features[1540]  | (\all_features[1538]  & \all_features[1539]  & \all_features[1537] ));
  assign new_n23248_ = ~\all_features[1543]  & (~\all_features[1542]  | ~new_n23249_ | ~new_n23250_ | ~new_n23251_);
  assign new_n23249_ = \all_features[1538]  & \all_features[1539] ;
  assign new_n23250_ = \all_features[1536]  & \all_features[1537] ;
  assign new_n23251_ = \all_features[1540]  & \all_features[1541] ;
  assign new_n23252_ = \all_features[1543]  & (\all_features[1542]  | (\all_features[1541]  & (\all_features[1540]  | ~new_n23254_ | ~new_n23253_)));
  assign new_n23253_ = ~\all_features[1536]  & ~\all_features[1537] ;
  assign new_n23254_ = ~\all_features[1538]  & ~\all_features[1539] ;
  assign new_n23255_ = \all_features[1543]  & (\all_features[1542]  | (new_n23251_ & (\all_features[1538]  | \all_features[1539]  | \all_features[1537] )));
  assign new_n23256_ = ~\all_features[1541]  & \all_features[1542]  & \all_features[1543]  & (\all_features[1540]  ? new_n23254_ : (new_n23250_ | ~new_n23254_));
  assign new_n23257_ = \all_features[1543]  & (\all_features[1541]  | \all_features[1542]  | \all_features[1540] );
  assign new_n23258_ = new_n23259_ & (~\all_features[1541]  | (~\all_features[1540]  & (~\all_features[1539]  | (~\all_features[1538]  & ~\all_features[1537] ))));
  assign new_n23259_ = ~\all_features[1542]  & ~\all_features[1543] ;
  assign new_n23260_ = ~\all_features[1541]  & new_n23259_ & ((~\all_features[1538]  & new_n23253_) | ~\all_features[1540]  | ~\all_features[1539] );
  assign new_n23261_ = ~\all_features[1543]  & (~\all_features[1542]  | (~\all_features[1541]  & (new_n23253_ | ~new_n23249_ | ~\all_features[1540] )));
  assign new_n23262_ = new_n23259_ & (~\all_features[1539]  | ~new_n23251_ | (~\all_features[1538]  & ~new_n23250_));
  assign new_n23263_ = ~\all_features[1543]  & (~\all_features[1542]  | (~\all_features[1540]  & ~\all_features[1541]  & ~new_n23249_));
  assign new_n23264_ = new_n23269_ & (~new_n23270_ | (~new_n23265_ & ~new_n23261_ & ~new_n23263_));
  assign new_n23265_ = ~new_n23246_ & ~new_n23248_ & (~new_n23257_ | ~new_n23252_ | new_n23266_);
  assign new_n23266_ = new_n23255_ & new_n23267_ & (new_n23268_ | ~\all_features[1541]  | ~\all_features[1542]  | ~\all_features[1543] );
  assign new_n23267_ = \all_features[1542]  & \all_features[1543]  & (\all_features[1540]  | \all_features[1541]  | new_n23250_ | ~new_n23254_);
  assign new_n23268_ = ~\all_features[1539]  & ~\all_features[1540]  & (~\all_features[1538]  | new_n23253_);
  assign new_n23269_ = ~new_n23260_ & (\all_features[1539]  | \all_features[1540]  | \all_features[1541]  | \all_features[1542]  | \all_features[1543] );
  assign new_n23270_ = ~new_n23258_ & ~new_n23262_;
  assign new_n23271_ = new_n23272_ & new_n23269_ & ~new_n23262_ & ~new_n23261_ & ~new_n23246_ & ~new_n23258_;
  assign new_n23272_ = ~new_n23248_ & ~new_n23263_;
  assign new_n23273_ = new_n23269_ & new_n23270_ & (new_n23274_ | new_n23246_ | new_n23261_ | ~new_n23272_);
  assign new_n23274_ = new_n23257_ & new_n23267_ & new_n23252_ & new_n23255_;
  assign new_n23275_ = ~new_n23321_ & new_n23276_;
  assign new_n23276_ = new_n23277_ & (new_n23318_ | ~new_n23320_) & (~new_n11615_ | ~new_n23316_);
  assign new_n23277_ = ~new_n23280_ & (~new_n23315_ | ~new_n23278_) & (~new_n22051_ | ~new_n23314_);
  assign new_n23278_ = new_n23279_ & ~new_n23133_ & new_n19157_;
  assign new_n23279_ = ~new_n23193_ & ~new_n10024_;
  assign new_n23280_ = new_n23279_ & (new_n23133_ ? new_n23281_ : ~new_n19157_);
  assign new_n23281_ = ~new_n23313_ & ~new_n23282_ & ((~new_n23283_ & ~new_n23308_) | new_n23310_ | ~new_n23304_);
  assign new_n23282_ = ~new_n6495_ & new_n16852_;
  assign new_n23283_ = ~new_n23297_ & (new_n23299_ | (~new_n23300_ & (new_n23301_ | (~new_n23284_ & ~new_n23302_))));
  assign new_n23284_ = ~new_n23291_ & (~new_n23295_ | (new_n23285_ & (~new_n23294_ | (~new_n23296_ & new_n23288_))));
  assign new_n23285_ = \all_features[3399]  & (\all_features[3398]  | new_n23286_);
  assign new_n23286_ = \all_features[3397]  & (\all_features[3394]  | \all_features[3395]  | \all_features[3396]  | ~new_n23287_);
  assign new_n23287_ = ~\all_features[3392]  & ~\all_features[3393] ;
  assign new_n23288_ = \all_features[3399]  & ~new_n23289_ & \all_features[3398] ;
  assign new_n23289_ = ~\all_features[3397]  & ~\all_features[3396]  & ~\all_features[3395]  & ~new_n23290_ & ~\all_features[3394] ;
  assign new_n23290_ = \all_features[3392]  & \all_features[3393] ;
  assign new_n23291_ = ~\all_features[3399]  & (~\all_features[3398]  | ~new_n23290_ | ~new_n23292_ | ~new_n23293_);
  assign new_n23292_ = \all_features[3396]  & \all_features[3397] ;
  assign new_n23293_ = \all_features[3394]  & \all_features[3395] ;
  assign new_n23294_ = \all_features[3399]  & (\all_features[3398]  | (new_n23292_ & (\all_features[3394]  | \all_features[3395]  | \all_features[3393] )));
  assign new_n23295_ = \all_features[3399]  & (\all_features[3397]  | \all_features[3398]  | \all_features[3396] );
  assign new_n23296_ = \all_features[3398]  & \all_features[3399]  & (\all_features[3397]  | (\all_features[3396]  & (\all_features[3395]  | \all_features[3394] )));
  assign new_n23297_ = new_n23298_ & (~\all_features[3397]  | (~\all_features[3396]  & (~\all_features[3395]  | (~\all_features[3394]  & ~\all_features[3393] ))));
  assign new_n23298_ = ~\all_features[3398]  & ~\all_features[3399] ;
  assign new_n23299_ = new_n23298_ & (~\all_features[3395]  | ~new_n23292_ | (~\all_features[3394]  & ~new_n23290_));
  assign new_n23300_ = ~\all_features[3399]  & (~\all_features[3398]  | (~\all_features[3396]  & ~\all_features[3397]  & ~new_n23293_));
  assign new_n23301_ = ~\all_features[3399]  & (~\all_features[3398]  | (~\all_features[3397]  & (new_n23287_ | ~new_n23293_ | ~\all_features[3396] )));
  assign new_n23302_ = ~new_n23303_ & ~\all_features[3399] ;
  assign new_n23303_ = \all_features[3397]  & \all_features[3398]  & (\all_features[3396]  | (\all_features[3394]  & \all_features[3395]  & \all_features[3393] ));
  assign new_n23304_ = ~new_n23301_ & new_n23306_ & ((new_n23285_ & new_n23305_) | new_n23302_ | ~new_n23309_);
  assign new_n23305_ = new_n23295_ & new_n23288_ & new_n23294_;
  assign new_n23306_ = new_n23307_ & ~new_n23300_ & ~new_n23308_ & ~new_n23297_;
  assign new_n23307_ = ~new_n23299_ & (\all_features[3395]  | \all_features[3396]  | \all_features[3397]  | \all_features[3398]  | \all_features[3399] );
  assign new_n23308_ = ~\all_features[3397]  & new_n23298_ & ((~\all_features[3394]  & new_n23287_) | ~\all_features[3396]  | ~\all_features[3395] );
  assign new_n23309_ = ~new_n23300_ & ~new_n23291_;
  assign new_n23310_ = ~new_n23291_ & ~new_n23302_ & (~new_n23295_ | new_n23311_ | ~new_n23285_);
  assign new_n23311_ = ~new_n23289_ & new_n23294_ & \all_features[3398]  & \all_features[3399]  & (~\all_features[3397]  | new_n23312_);
  assign new_n23312_ = ~\all_features[3395]  & ~\all_features[3396]  & (~\all_features[3394]  | new_n23287_);
  assign new_n23313_ = new_n23309_ & new_n23307_ & ~new_n23302_ & ~new_n23301_ & ~new_n23308_ & ~new_n23297_;
  assign new_n23314_ = new_n23282_ & new_n23133_ & new_n23279_;
  assign new_n23315_ = ~new_n8059_ & (~new_n8056_ | ~new_n9644_);
  assign new_n23316_ = ~new_n22609_ & new_n23317_;
  assign new_n23317_ = ~new_n18385_ & ~new_n23279_;
  assign new_n23318_ = new_n23319_ ? new_n11060_ : new_n13887_;
  assign new_n23319_ = new_n12850_ & new_n17631_;
  assign new_n23320_ = ~new_n23279_ & new_n18385_;
  assign new_n23321_ = new_n23323_ & new_n23322_ & (new_n23315_ | ~new_n23278_);
  assign new_n23322_ = (~new_n23320_ | ~new_n23318_) & (new_n11615_ | ~new_n23316_);
  assign new_n23323_ = (~new_n23314_ | new_n22051_) & (~new_n23317_ | ~new_n22609_ | ~new_n23324_);
  assign new_n23324_ = new_n12375_ & new_n12731_;
  assign new_n23325_ = new_n23326_ & (new_n14278_ | ~new_n23334_ | ~new_n23342_ | ~new_n8927_);
  assign new_n23326_ = ~new_n23327_ & new_n23332_ & (~new_n23339_ | (new_n23341_ & new_n22602_) | (new_n23340_ & ~new_n22602_));
  assign new_n23327_ = new_n23328_ & (new_n6603_ ? (~new_n13242_ | (~new_n18110_ & ~new_n13238_)) : ~new_n23331_);
  assign new_n23328_ = ~new_n18420_ & ~new_n23329_;
  assign new_n23329_ = new_n23330_ & ~new_n23271_ & ~new_n23273_;
  assign new_n23330_ = ~new_n23243_ & ~new_n23264_;
  assign new_n23331_ = new_n22691_ & new_n22554_;
  assign new_n23332_ = (new_n15022_ | ~new_n14278_ | ~new_n23334_) & (~new_n23333_ | (new_n23337_ & new_n16102_));
  assign new_n23333_ = ~new_n18420_ & new_n23329_;
  assign new_n23334_ = ~new_n23335_ & new_n18420_;
  assign new_n23335_ = ~new_n23336_ & ~new_n17961_;
  assign new_n23336_ = new_n17939_ & new_n17964_;
  assign new_n23337_ = new_n18795_ & new_n23338_;
  assign new_n23338_ = new_n6950_ & new_n6953_;
  assign new_n23339_ = new_n18420_ & new_n23335_;
  assign new_n23340_ = new_n22423_ & (new_n22420_ | ~new_n22390_);
  assign new_n23341_ = new_n9129_ & (new_n9131_ | new_n9122_);
  assign new_n23342_ = ~new_n23344_ & new_n23343_ & (~new_n23334_ | (~new_n15022_ & new_n14278_) | (new_n8927_ & ~new_n14278_));
  assign new_n23343_ = (~new_n23333_ | ~new_n16102_ | ~new_n23337_) & (new_n6603_ | ~new_n23331_ | ~new_n23328_);
  assign new_n23344_ = new_n23339_ & (new_n22602_ ? new_n23341_ : new_n23340_);
  assign \o[29]  = new_n23346_ ? (new_n23347_ ^ new_n23348_) : (~new_n23347_ ^ new_n23348_);
  assign new_n23346_ = (new_n23275_ & new_n23325_) | (~new_n22265_ & (new_n23275_ | new_n23325_));
  assign new_n23347_ = (new_n23181_ & new_n23197_) | (~new_n22266_ & (new_n23181_ | new_n23197_));
  assign new_n23348_ = new_n23349_ ? (~new_n23350_ ^ new_n23387_) : (new_n23350_ ^ new_n23387_);
  assign new_n23349_ = (~new_n23126_ & new_n23165_) | (~new_n22267_ & (~new_n23126_ | new_n23165_));
  assign new_n23350_ = new_n23351_ ? (new_n23352_ ^ new_n23384_) : (~new_n23352_ ^ new_n23384_);
  assign new_n23351_ = (~new_n22830_ & new_n23082_) | (~new_n22268_ & (~new_n22830_ | new_n23082_));
  assign new_n23352_ = new_n23353_ ? (new_n23363_ ^ new_n23364_) : (~new_n23363_ ^ new_n23364_);
  assign new_n23353_ = new_n23354_ ? (~new_n23355_ ^ new_n23362_) : (new_n23355_ ^ new_n23362_);
  assign new_n23354_ = (new_n22434_ & new_n22463_) | (~new_n22270_ & (new_n22434_ | new_n22463_));
  assign new_n23355_ = new_n23356_ ? (~new_n23360_ ^ new_n23361_) : (new_n23360_ ^ new_n23361_);
  assign new_n23356_ = new_n23357_ ? (new_n23358_ ^ new_n23359_) : (~new_n23358_ ^ new_n23359_);
  assign new_n23357_ = new_n22351_ & new_n22375_;
  assign new_n23358_ = new_n22378_ & new_n22430_;
  assign new_n23359_ = ~new_n23125_ & new_n23083_;
  assign new_n23360_ = (new_n22953_ & new_n22991_) | (new_n22944_ & (new_n22953_ | new_n22991_));
  assign new_n23361_ = new_n22954_ & new_n22990_;
  assign new_n23362_ = (~new_n22943_ & new_n22999_) | (~new_n22832_ & (~new_n22943_ | new_n22999_));
  assign new_n23363_ = (~new_n22535_ & new_n22792_) | (~new_n22269_ & (~new_n22535_ | new_n22792_));
  assign new_n23364_ = new_n23365_ ? (new_n23372_ ^ new_n23373_) : (~new_n23372_ ^ new_n23373_);
  assign new_n23365_ = new_n23366_ ? (~new_n23367_ ^ new_n23371_) : (new_n23367_ ^ new_n23371_);
  assign new_n23366_ = (new_n22350_ & new_n22377_) | (new_n22271_ & (new_n22350_ | new_n22377_));
  assign new_n23367_ = new_n23368_ ? (new_n23369_ ^ new_n23370_) : (~new_n23369_ ^ new_n23370_);
  assign new_n23368_ = new_n22272_ & new_n22348_;
  assign new_n23369_ = new_n23128_ & new_n23141_;
  assign new_n23370_ = new_n23166_ & new_n23176_;
  assign new_n23371_ = (new_n22704_ & new_n22769_) | (new_n22650_ & (new_n22704_ | new_n22769_));
  assign new_n23372_ = (~new_n22649_ & new_n22781_) | (~new_n22536_ & (~new_n22649_ | new_n22781_));
  assign new_n23373_ = new_n23374_ ? (~new_n23375_ ^ new_n23379_) : (new_n23375_ ^ new_n23379_);
  assign new_n23374_ = ~new_n22537_ & ~new_n22598_;
  assign new_n23375_ = new_n23376_ ? (new_n23377_ ^ new_n23378_) : (~new_n23377_ ^ new_n23378_);
  assign new_n23376_ = new_n23276_ & new_n23321_;
  assign new_n23377_ = new_n22651_ & new_n22699_;
  assign new_n23378_ = new_n22599_ & new_n22646_;
  assign new_n23379_ = new_n23380_ ^ new_n23383_;
  assign new_n23380_ = new_n22595_ & ~new_n23382_ & new_n23381_;
  assign new_n23381_ = new_n22539_ & (new_n10910_ | ~new_n22541_ | ~new_n22562_);
  assign new_n23382_ = ~new_n22547_ & ~new_n22551_;
  assign new_n23383_ = new_n23326_ & new_n23342_;
  assign new_n23384_ = ~new_n23385_ ^ new_n23386_;
  assign new_n23385_ = (new_n23060_ & new_n23073_) | (~new_n22831_ & (new_n23060_ | new_n23073_));
  assign new_n23386_ = (new_n22895_ & new_n22935_) | (new_n22833_ & (new_n22895_ | new_n22935_));
  assign new_n23387_ = (new_n23143_ & new_n23154_) | (new_n23127_ & (new_n23143_ | new_n23154_));
  assign \o[30]  = ~new_n23389_ ^ new_n23390_;
  assign new_n23389_ = (~new_n23348_ & new_n23347_) | (new_n23346_ & (~new_n23348_ | new_n23347_));
  assign new_n23390_ = new_n23391_ ^ new_n23392_;
  assign new_n23391_ = (~new_n23350_ & new_n23387_) | (new_n23349_ & (~new_n23350_ | new_n23387_));
  assign new_n23392_ = new_n23393_ ? (~new_n23394_ ^ new_n23411_) : (new_n23394_ ^ new_n23411_);
  assign new_n23393_ = (~new_n23352_ & ~new_n23384_) | (new_n23351_ & (~new_n23352_ | ~new_n23384_));
  assign new_n23394_ = new_n23395_ ? (~new_n23396_ ^ new_n23410_) : (new_n23396_ ^ new_n23410_);
  assign new_n23395_ = (~new_n23364_ & new_n23363_) | (~new_n23353_ & (~new_n23364_ | new_n23363_));
  assign new_n23396_ = new_n23397_ ? (new_n23401_ ^ new_n23402_) : (~new_n23401_ ^ new_n23402_);
  assign new_n23397_ = new_n23398_ ? (new_n23399_ ^ new_n23400_) : (~new_n23399_ ^ new_n23400_);
  assign new_n23398_ = (~new_n23367_ & new_n23371_) | (new_n23366_ & (~new_n23367_ | new_n23371_));
  assign new_n23399_ = (new_n23360_ & new_n23361_) | (~new_n23356_ & (new_n23360_ | new_n23361_));
  assign new_n23400_ = (new_n23358_ & new_n23359_) | (new_n23357_ & (new_n23358_ | new_n23359_));
  assign new_n23401_ = (~new_n23373_ & new_n23372_) | (~new_n23365_ & (~new_n23373_ | new_n23372_));
  assign new_n23402_ = new_n23403_ ? (new_n23406_ ^ new_n23407_) : (~new_n23406_ ^ new_n23407_);
  assign new_n23403_ = ~new_n23404_ ^ new_n23405_;
  assign new_n23404_ = (new_n23369_ & new_n23370_) | (new_n23368_ & (new_n23369_ | new_n23370_));
  assign new_n23405_ = (new_n23377_ & new_n23378_) | (new_n23376_ & (new_n23377_ | new_n23378_));
  assign new_n23406_ = (~new_n23375_ & ~new_n23379_) | (~new_n23374_ & (~new_n23375_ | ~new_n23379_));
  assign new_n23407_ = new_n23408_ ^ new_n23409_;
  assign new_n23408_ = ~new_n23380_ & ~new_n23383_;
  assign new_n23409_ = new_n22595_ & new_n23381_ & new_n23382_;
  assign new_n23410_ = (~new_n23355_ & new_n23362_) | (new_n23354_ & (~new_n23355_ | new_n23362_));
  assign new_n23411_ = new_n23385_ & new_n23386_;
  assign \o[31]  = ((new_n23413_ | new_n23414_) & (new_n23415_ ^ new_n23416_)) | (~new_n23413_ & ~new_n23414_ & (~new_n23415_ ^ new_n23416_));
  assign new_n23413_ = ~new_n23390_ & new_n23389_;
  assign new_n23414_ = ~new_n23392_ & new_n23391_;
  assign new_n23415_ = (~new_n23394_ & new_n23411_) | (new_n23393_ & (~new_n23394_ | new_n23411_));
  assign new_n23416_ = ~new_n23417_ ^ new_n23418_;
  assign new_n23417_ = (~new_n23396_ & new_n23410_) | (new_n23395_ & (~new_n23396_ | new_n23410_));
  assign new_n23418_ = new_n23419_ ? (new_n23420_ ^ new_n23424_) : (~new_n23420_ ^ new_n23424_);
  assign new_n23419_ = (~new_n23402_ & new_n23401_) | (~new_n23397_ & (~new_n23402_ | new_n23401_));
  assign new_n23420_ = new_n23421_ ? (new_n23422_ ^ new_n23423_) : (~new_n23422_ ^ new_n23423_);
  assign new_n23421_ = (~new_n23407_ & new_n23406_) | (~new_n23403_ & (~new_n23407_ | new_n23406_));
  assign new_n23422_ = new_n23404_ & new_n23405_;
  assign new_n23423_ = ~new_n23408_ & new_n23409_;
  assign new_n23424_ = (new_n23399_ & new_n23400_) | (new_n23398_ & (new_n23399_ | new_n23400_));
  assign \o[32]  = ~new_n23426_ ^ new_n23427_;
  assign new_n23426_ = (new_n23415_ | (~new_n23416_ & (new_n23414_ | new_n23413_))) & (new_n23414_ | new_n23413_ | ~new_n23416_);
  assign new_n23427_ = new_n23428_ ^ new_n23429_;
  assign new_n23428_ = new_n23417_ & new_n23418_;
  assign new_n23429_ = ~new_n23430_ ^ new_n23431_;
  assign new_n23430_ = (~new_n23420_ & new_n23424_) | (new_n23419_ & (~new_n23420_ | new_n23424_));
  assign new_n23431_ = (new_n23422_ & new_n23423_) | (new_n23421_ & (new_n23422_ | new_n23423_));
  assign \o[33]  = (~new_n23435_ & (new_n23433_ | new_n23434_)) | (~new_n23433_ & ~new_n23434_ & new_n23435_);
  assign new_n23433_ = ~new_n23427_ & new_n23426_;
  assign new_n23434_ = ~new_n23429_ & new_n23428_;
  assign new_n23435_ = new_n23430_ & new_n23431_;
  assign \o[34]  = new_n23435_ & (new_n23434_ | new_n23433_);
  assign \o[35]  = new_n23438_ ^ new_n24559_;
  assign new_n23438_ = new_n23439_ ? (~new_n24366_ ^ new_n24542_) : (new_n24366_ ^ new_n24542_);
  assign new_n23439_ = new_n23440_ ? (new_n24124_ ^ new_n24353_) : (~new_n24124_ ^ new_n24353_);
  assign new_n23440_ = new_n23441_ ? (new_n23940_ ^ new_n24114_) : (~new_n23940_ ^ new_n24114_);
  assign new_n23441_ = new_n23442_ ? (new_n23773_ ^ new_n23931_) : (~new_n23773_ ^ new_n23931_);
  assign new_n23442_ = new_n23443_ ? (new_n23601_ ^ new_n23659_) : (~new_n23601_ ^ new_n23659_);
  assign new_n23443_ = ~new_n23444_ & new_n23599_;
  assign new_n23444_ = new_n23445_ & (~new_n23548_ | ~new_n23550_ | ~new_n23554_ | ~new_n23480_);
  assign new_n23445_ = ~new_n23446_ & new_n23481_ & (~new_n23480_ | (new_n23550_ & new_n23548_) | (~new_n23552_ & ~new_n23548_));
  assign new_n23446_ = new_n23447_ & new_n23450_;
  assign new_n23447_ = ~new_n20087_ & new_n23448_;
  assign new_n23448_ = ~new_n23449_ & new_n18750_;
  assign new_n23449_ = ~new_n9065_ & new_n23179_;
  assign new_n23450_ = ~new_n23451_ & new_n23475_;
  assign new_n23451_ = new_n23467_ & (~new_n23470_ | (~new_n23452_ & ~new_n23473_ & ~new_n23474_));
  assign new_n23452_ = ~new_n23461_ & ~new_n23463_ & (~new_n23466_ | ~new_n23465_ | new_n23453_);
  assign new_n23453_ = new_n23454_ & new_n23456_ & (new_n23459_ | ~\all_features[2645]  | ~\all_features[2646]  | ~\all_features[2647] );
  assign new_n23454_ = \all_features[2647]  & (\all_features[2646]  | (new_n23455_ & (\all_features[2642]  | \all_features[2643]  | \all_features[2641] )));
  assign new_n23455_ = \all_features[2644]  & \all_features[2645] ;
  assign new_n23456_ = \all_features[2646]  & \all_features[2647]  & (\all_features[2644]  | \all_features[2645]  | new_n23457_ | ~new_n23458_);
  assign new_n23457_ = \all_features[2640]  & \all_features[2641] ;
  assign new_n23458_ = ~\all_features[2642]  & ~\all_features[2643] ;
  assign new_n23459_ = ~\all_features[2643]  & ~\all_features[2644]  & (~\all_features[2642]  | new_n23460_);
  assign new_n23460_ = ~\all_features[2640]  & ~\all_features[2641] ;
  assign new_n23461_ = ~new_n23462_ & ~\all_features[2647] ;
  assign new_n23462_ = \all_features[2645]  & \all_features[2646]  & (\all_features[2644]  | (\all_features[2642]  & \all_features[2643]  & \all_features[2641] ));
  assign new_n23463_ = ~\all_features[2647]  & (~\all_features[2646]  | ~new_n23464_ | ~new_n23457_ | ~new_n23455_);
  assign new_n23464_ = \all_features[2642]  & \all_features[2643] ;
  assign new_n23465_ = \all_features[2647]  & (\all_features[2646]  | (\all_features[2645]  & (\all_features[2644]  | ~new_n23458_ | ~new_n23460_)));
  assign new_n23466_ = \all_features[2647]  & (\all_features[2645]  | \all_features[2646]  | \all_features[2644] );
  assign new_n23467_ = ~new_n23468_ & (\all_features[2643]  | \all_features[2644]  | \all_features[2645]  | \all_features[2646]  | \all_features[2647] );
  assign new_n23468_ = ~\all_features[2645]  & new_n23469_ & ((~\all_features[2642]  & new_n23460_) | ~\all_features[2644]  | ~\all_features[2643] );
  assign new_n23469_ = ~\all_features[2646]  & ~\all_features[2647] ;
  assign new_n23470_ = ~new_n23471_ & ~new_n23472_;
  assign new_n23471_ = new_n23469_ & (~\all_features[2645]  | (~\all_features[2644]  & (~\all_features[2643]  | (~\all_features[2642]  & ~\all_features[2641] ))));
  assign new_n23472_ = new_n23469_ & (~\all_features[2643]  | ~new_n23455_ | (~\all_features[2642]  & ~new_n23457_));
  assign new_n23473_ = ~\all_features[2647]  & (~\all_features[2646]  | (~\all_features[2645]  & (new_n23460_ | ~new_n23464_ | ~\all_features[2644] )));
  assign new_n23474_ = ~\all_features[2647]  & (~\all_features[2646]  | (~\all_features[2644]  & ~\all_features[2645]  & ~new_n23464_));
  assign new_n23475_ = ~new_n23476_ & ~new_n23478_;
  assign new_n23476_ = new_n23477_ & new_n23467_ & ~new_n23472_ & ~new_n23473_ & ~new_n23461_ & ~new_n23471_;
  assign new_n23477_ = ~new_n23463_ & ~new_n23474_;
  assign new_n23478_ = new_n23467_ & new_n23470_ & (new_n23479_ | new_n23461_ | new_n23473_ | ~new_n23477_);
  assign new_n23479_ = new_n23466_ & new_n23456_ & new_n23465_ & new_n23454_;
  assign new_n23480_ = ~new_n23449_ & ~new_n18750_;
  assign new_n23481_ = ~new_n23449_ | ~new_n23515_ | (new_n23482_ ? ~new_n14162_ : new_n14435_);
  assign new_n23482_ = ~new_n23483_ & new_n23510_;
  assign new_n23483_ = ~new_n23509_ & (~new_n23502_ | (~new_n23507_ & (new_n23500_ | new_n23508_ | ~new_n23484_)));
  assign new_n23484_ = ~new_n23496_ & ~new_n23494_ & ((~new_n23491_ & new_n23485_) | ~new_n23499_ | ~new_n23498_);
  assign new_n23485_ = \all_features[2223]  & \all_features[2222]  & ~new_n23488_ & new_n23486_;
  assign new_n23486_ = \all_features[2223]  & (\all_features[2222]  | (new_n23487_ & (\all_features[2218]  | \all_features[2219]  | \all_features[2217] )));
  assign new_n23487_ = \all_features[2220]  & \all_features[2221] ;
  assign new_n23488_ = new_n23490_ & ~\all_features[2221]  & ~new_n23489_ & ~\all_features[2220] ;
  assign new_n23489_ = \all_features[2216]  & \all_features[2217] ;
  assign new_n23490_ = ~\all_features[2218]  & ~\all_features[2219] ;
  assign new_n23491_ = \all_features[2223]  & \all_features[2222]  & ~new_n23492_ & \all_features[2221] ;
  assign new_n23492_ = ~\all_features[2219]  & ~\all_features[2220]  & (~\all_features[2218]  | new_n23493_);
  assign new_n23493_ = ~\all_features[2216]  & ~\all_features[2217] ;
  assign new_n23494_ = ~new_n23495_ & ~\all_features[2223] ;
  assign new_n23495_ = \all_features[2221]  & \all_features[2222]  & (\all_features[2220]  | (\all_features[2218]  & \all_features[2219]  & \all_features[2217] ));
  assign new_n23496_ = ~\all_features[2223]  & (~\all_features[2222]  | ~new_n23497_ | ~new_n23489_ | ~new_n23487_);
  assign new_n23497_ = \all_features[2218]  & \all_features[2219] ;
  assign new_n23498_ = \all_features[2223]  & (\all_features[2222]  | (\all_features[2221]  & (\all_features[2220]  | ~new_n23490_ | ~new_n23493_)));
  assign new_n23499_ = \all_features[2223]  & (\all_features[2221]  | \all_features[2222]  | \all_features[2220] );
  assign new_n23500_ = ~new_n23494_ & (new_n23496_ | (new_n23499_ & (~new_n23498_ | (~new_n23501_ & new_n23486_))));
  assign new_n23501_ = ~\all_features[2221]  & \all_features[2222]  & \all_features[2223]  & (\all_features[2220]  ? new_n23490_ : (new_n23489_ | ~new_n23490_));
  assign new_n23502_ = ~new_n23506_ & ~new_n23503_ & ~new_n23505_;
  assign new_n23503_ = new_n23504_ & (~\all_features[2221]  | (~\all_features[2220]  & (~\all_features[2219]  | (~\all_features[2218]  & ~\all_features[2217] ))));
  assign new_n23504_ = ~\all_features[2222]  & ~\all_features[2223] ;
  assign new_n23505_ = ~\all_features[2221]  & new_n23504_ & ((~\all_features[2218]  & new_n23493_) | ~\all_features[2220]  | ~\all_features[2219] );
  assign new_n23506_ = new_n23504_ & (~\all_features[2219]  | ~new_n23487_ | (~\all_features[2218]  & ~new_n23489_));
  assign new_n23507_ = ~\all_features[2223]  & (~\all_features[2222]  | (~\all_features[2220]  & ~\all_features[2221]  & ~new_n23497_));
  assign new_n23508_ = ~\all_features[2223]  & (~\all_features[2222]  | (~\all_features[2221]  & (new_n23493_ | ~\all_features[2220]  | ~new_n23497_)));
  assign new_n23509_ = ~\all_features[2223]  & ~\all_features[2222]  & ~\all_features[2221]  & ~\all_features[2219]  & ~\all_features[2220] ;
  assign new_n23510_ = new_n23503_ | ~new_n23513_ | ((new_n23494_ | ~new_n23514_) & (new_n23511_ | new_n23506_));
  assign new_n23511_ = new_n23512_ & (~new_n23485_ | ~new_n23498_ | ~new_n23499_);
  assign new_n23512_ = ~new_n23496_ & ~new_n23494_ & ~new_n23507_ & ~new_n23508_;
  assign new_n23513_ = ~new_n23505_ & ~new_n23509_;
  assign new_n23514_ = ~new_n23506_ & ~new_n23496_ & ~new_n23507_ & ~new_n23508_;
  assign new_n23515_ = ~new_n23516_ & new_n23543_;
  assign new_n23516_ = ~new_n23542_ & (~new_n23535_ | (~new_n23540_ & (new_n23533_ | new_n23541_ | ~new_n23517_)));
  assign new_n23517_ = ~new_n23529_ & ~new_n23527_ & ((~new_n23524_ & new_n23518_) | ~new_n23532_ | ~new_n23531_);
  assign new_n23518_ = \all_features[1311]  & \all_features[1310]  & ~new_n23521_ & new_n23519_;
  assign new_n23519_ = \all_features[1311]  & (\all_features[1310]  | (new_n23520_ & (\all_features[1306]  | \all_features[1307]  | \all_features[1305] )));
  assign new_n23520_ = \all_features[1308]  & \all_features[1309] ;
  assign new_n23521_ = new_n23523_ & ~\all_features[1309]  & ~new_n23522_ & ~\all_features[1308] ;
  assign new_n23522_ = \all_features[1304]  & \all_features[1305] ;
  assign new_n23523_ = ~\all_features[1306]  & ~\all_features[1307] ;
  assign new_n23524_ = \all_features[1311]  & \all_features[1310]  & ~new_n23525_ & \all_features[1309] ;
  assign new_n23525_ = ~\all_features[1307]  & ~\all_features[1308]  & (~\all_features[1306]  | new_n23526_);
  assign new_n23526_ = ~\all_features[1304]  & ~\all_features[1305] ;
  assign new_n23527_ = ~new_n23528_ & ~\all_features[1311] ;
  assign new_n23528_ = \all_features[1309]  & \all_features[1310]  & (\all_features[1308]  | (\all_features[1306]  & \all_features[1307]  & \all_features[1305] ));
  assign new_n23529_ = ~\all_features[1311]  & (~\all_features[1310]  | ~new_n23530_ | ~new_n23522_ | ~new_n23520_);
  assign new_n23530_ = \all_features[1306]  & \all_features[1307] ;
  assign new_n23531_ = \all_features[1311]  & (\all_features[1310]  | (\all_features[1309]  & (\all_features[1308]  | ~new_n23523_ | ~new_n23526_)));
  assign new_n23532_ = \all_features[1311]  & (\all_features[1309]  | \all_features[1310]  | \all_features[1308] );
  assign new_n23533_ = ~new_n23527_ & (new_n23529_ | (new_n23532_ & (~new_n23531_ | (~new_n23534_ & new_n23519_))));
  assign new_n23534_ = ~\all_features[1309]  & \all_features[1310]  & \all_features[1311]  & (\all_features[1308]  ? new_n23523_ : (new_n23522_ | ~new_n23523_));
  assign new_n23535_ = ~new_n23539_ & ~new_n23536_ & ~new_n23538_;
  assign new_n23536_ = new_n23537_ & (~\all_features[1309]  | (~\all_features[1308]  & (~\all_features[1307]  | (~\all_features[1306]  & ~\all_features[1305] ))));
  assign new_n23537_ = ~\all_features[1310]  & ~\all_features[1311] ;
  assign new_n23538_ = ~\all_features[1309]  & new_n23537_ & ((~\all_features[1306]  & new_n23526_) | ~\all_features[1308]  | ~\all_features[1307] );
  assign new_n23539_ = new_n23537_ & (~\all_features[1307]  | ~new_n23520_ | (~\all_features[1306]  & ~new_n23522_));
  assign new_n23540_ = ~\all_features[1311]  & (~\all_features[1310]  | (~\all_features[1308]  & ~\all_features[1309]  & ~new_n23530_));
  assign new_n23541_ = ~\all_features[1311]  & (~\all_features[1310]  | (~\all_features[1309]  & (new_n23526_ | ~\all_features[1308]  | ~new_n23530_)));
  assign new_n23542_ = ~\all_features[1311]  & ~\all_features[1310]  & ~\all_features[1309]  & ~\all_features[1307]  & ~\all_features[1308] ;
  assign new_n23543_ = new_n23536_ | ~new_n23546_ | ((new_n23527_ | ~new_n23547_) & (new_n23544_ | new_n23539_));
  assign new_n23544_ = new_n23545_ & (~new_n23518_ | ~new_n23531_ | ~new_n23532_);
  assign new_n23545_ = ~new_n23529_ & ~new_n23527_ & ~new_n23540_ & ~new_n23541_;
  assign new_n23546_ = ~new_n23538_ & ~new_n23542_;
  assign new_n23547_ = ~new_n23539_ & ~new_n23529_ & ~new_n23540_ & ~new_n23541_;
  assign new_n23548_ = new_n18961_ & new_n23549_;
  assign new_n23549_ = ~new_n20443_ & ~new_n20447_;
  assign new_n23550_ = ~new_n15497_ & new_n23551_;
  assign new_n23551_ = new_n15528_ & new_n15530_;
  assign new_n23552_ = new_n23551_ & new_n23553_;
  assign new_n23553_ = new_n15498_ & new_n15518_;
  assign new_n23554_ = ~new_n23555_ & (~new_n23448_ | ~new_n18786_ | ~new_n20087_);
  assign new_n23555_ = ~new_n23515_ & new_n23449_ & (new_n23556_ ? ~new_n23598_ : new_n23592_);
  assign new_n23556_ = new_n23557_ & new_n23583_;
  assign new_n23557_ = ~new_n23558_ & ~new_n23581_;
  assign new_n23558_ = new_n23578_ & ~new_n23559_ & new_n23575_;
  assign new_n23559_ = ~new_n23574_ & ~new_n23573_ & ~new_n23571_ & ~new_n23560_ & ~new_n23563_;
  assign new_n23560_ = ~\all_features[2183]  & (~\all_features[2182]  | new_n23561_);
  assign new_n23561_ = ~\all_features[2181]  & (new_n23562_ | ~\all_features[2179]  | ~\all_features[2180]  | ~\all_features[2178] );
  assign new_n23562_ = ~\all_features[2176]  & ~\all_features[2177] ;
  assign new_n23563_ = new_n23570_ & new_n23569_ & new_n23564_ & new_n23566_;
  assign new_n23564_ = \all_features[2183]  & (\all_features[2182]  | (new_n23565_ & (\all_features[2178]  | \all_features[2179]  | \all_features[2177] )));
  assign new_n23565_ = \all_features[2180]  & \all_features[2181] ;
  assign new_n23566_ = \all_features[2182]  & \all_features[2183]  & (\all_features[2180]  | \all_features[2181]  | new_n23568_ | ~new_n23567_);
  assign new_n23567_ = ~\all_features[2178]  & ~\all_features[2179] ;
  assign new_n23568_ = \all_features[2176]  & \all_features[2177] ;
  assign new_n23569_ = \all_features[2183]  & (\all_features[2182]  | (\all_features[2181]  & (\all_features[2180]  | ~new_n23567_ | ~new_n23562_)));
  assign new_n23570_ = \all_features[2183]  & (\all_features[2181]  | \all_features[2182]  | \all_features[2180] );
  assign new_n23571_ = ~new_n23572_ & ~\all_features[2183] ;
  assign new_n23572_ = \all_features[2181]  & \all_features[2182]  & (\all_features[2180]  | (\all_features[2178]  & \all_features[2179]  & \all_features[2177] ));
  assign new_n23573_ = ~\all_features[2183]  & (~new_n23568_ | ~\all_features[2178]  | ~\all_features[2179]  | ~\all_features[2182]  | ~new_n23565_);
  assign new_n23574_ = ~\all_features[2183]  & (~\all_features[2182]  | (~\all_features[2181]  & ~\all_features[2180]  & (~\all_features[2179]  | ~\all_features[2178] )));
  assign new_n23575_ = ~new_n23576_ & (\all_features[2179]  | \all_features[2180]  | \all_features[2181]  | \all_features[2182]  | \all_features[2183] );
  assign new_n23576_ = ~\all_features[2181]  & new_n23577_ & ((~\all_features[2178]  & new_n23562_) | ~\all_features[2180]  | ~\all_features[2179] );
  assign new_n23577_ = ~\all_features[2182]  & ~\all_features[2183] ;
  assign new_n23578_ = ~new_n23579_ & ~new_n23580_;
  assign new_n23579_ = new_n23577_ & (~\all_features[2181]  | (~\all_features[2180]  & (~\all_features[2179]  | (~\all_features[2178]  & ~\all_features[2177] ))));
  assign new_n23580_ = new_n23577_ & (~\all_features[2179]  | ~new_n23565_ | (~new_n23568_ & ~\all_features[2178] ));
  assign new_n23581_ = new_n23575_ & new_n23582_ & ~new_n23571_ & ~new_n23579_;
  assign new_n23582_ = ~new_n23574_ & ~new_n23580_ & ~new_n23560_ & ~new_n23573_;
  assign new_n23583_ = ~new_n23584_ & ~new_n23588_;
  assign new_n23584_ = new_n23575_ & (~new_n23578_ | (~new_n23560_ & ~new_n23585_ & ~new_n23574_));
  assign new_n23585_ = ~new_n23573_ & ~new_n23571_ & (~new_n23570_ | ~new_n23569_ | new_n23586_);
  assign new_n23586_ = new_n23564_ & new_n23566_ & (new_n23587_ | ~\all_features[2181]  | ~\all_features[2182]  | ~\all_features[2183] );
  assign new_n23587_ = ~\all_features[2179]  & ~\all_features[2180]  & (~\all_features[2178]  | new_n23562_);
  assign new_n23588_ = ~new_n23589_ & (\all_features[2179]  | \all_features[2180]  | \all_features[2181]  | \all_features[2182]  | \all_features[2183] );
  assign new_n23589_ = ~new_n23576_ & (new_n23579_ | (~new_n23580_ & (new_n23574_ | (~new_n23560_ & ~new_n23590_))));
  assign new_n23590_ = ~new_n23571_ & (new_n23573_ | (new_n23570_ & (~new_n23569_ | (~new_n23591_ & new_n23564_))));
  assign new_n23591_ = ~\all_features[2181]  & \all_features[2182]  & \all_features[2183]  & (\all_features[2180]  ? new_n23567_ : (new_n23568_ | ~new_n23567_));
  assign new_n23592_ = new_n23593_ & ~new_n23003_ & ~new_n23032_;
  assign new_n23593_ = ~new_n23025_ & ~new_n23594_;
  assign new_n23594_ = ~new_n23595_ & (\all_features[2619]  | \all_features[2620]  | \all_features[2621]  | \all_features[2622]  | \all_features[2623] );
  assign new_n23595_ = ~new_n23021_ & (new_n23023_ | (~new_n23024_ & (new_n23014_ | (~new_n23006_ & ~new_n23596_))));
  assign new_n23596_ = ~new_n23009_ & (new_n23011_ | (new_n23019_ & (~new_n23015_ | (~new_n23597_ & new_n23017_))));
  assign new_n23597_ = ~\all_features[2621]  & \all_features[2622]  & \all_features[2623]  & (\all_features[2620]  ? new_n23016_ : (new_n23013_ | ~new_n23016_));
  assign new_n23598_ = new_n6702_ & new_n18812_;
  assign new_n23599_ = new_n23600_ & (new_n23450_ | ~new_n23447_) & (new_n23548_ | new_n23552_ | ~new_n23480_);
  assign new_n23600_ = ~new_n23449_ | ((new_n14162_ | ~new_n23482_ | ~new_n23515_) & (new_n23556_ | new_n23592_ | new_n23515_));
  assign new_n23601_ = new_n23602_ & (new_n23655_ | (new_n23656_ & new_n23658_));
  assign new_n23602_ = new_n23647_ & new_n23603_ & new_n23641_;
  assign new_n23603_ = (new_n23605_ | ~new_n14162_ | ~new_n23640_ | ~new_n7556_) & (new_n23604_ | new_n6354_ | new_n7556_);
  assign new_n23604_ = new_n6389_ & (new_n23239_ | new_n23200_ | ~new_n23221_);
  assign new_n23605_ = ~new_n23636_ & new_n23606_;
  assign new_n23606_ = ~new_n23632_ & new_n23607_;
  assign new_n23607_ = ~new_n23608_ & ~new_n23630_;
  assign new_n23608_ = new_n23625_ & ~new_n23629_ & ~new_n23609_ & ~new_n23628_;
  assign new_n23609_ = new_n23610_ & (~new_n23623_ | ~new_n23624_ | ~new_n23620_ | ~new_n23622_);
  assign new_n23610_ = ~new_n23617_ & ~new_n23615_ & ~new_n23611_ & ~new_n23613_;
  assign new_n23611_ = ~\all_features[2415]  & (~\all_features[2414]  | (~\all_features[2412]  & ~\all_features[2413]  & ~new_n23612_));
  assign new_n23612_ = \all_features[2410]  & \all_features[2411] ;
  assign new_n23613_ = ~\all_features[2415]  & (~\all_features[2414]  | (~\all_features[2413]  & (new_n23614_ | ~new_n23612_ | ~\all_features[2412] )));
  assign new_n23614_ = ~\all_features[2408]  & ~\all_features[2409] ;
  assign new_n23615_ = ~new_n23616_ & ~\all_features[2415] ;
  assign new_n23616_ = \all_features[2413]  & \all_features[2414]  & (\all_features[2412]  | (\all_features[2410]  & \all_features[2411]  & \all_features[2409] ));
  assign new_n23617_ = ~\all_features[2415]  & (~\all_features[2414]  | ~new_n23618_ | ~new_n23619_ | ~new_n23612_);
  assign new_n23618_ = \all_features[2408]  & \all_features[2409] ;
  assign new_n23619_ = \all_features[2412]  & \all_features[2413] ;
  assign new_n23620_ = \all_features[2415]  & (\all_features[2414]  | (\all_features[2413]  & (\all_features[2412]  | ~new_n23621_ | ~new_n23614_)));
  assign new_n23621_ = ~\all_features[2410]  & ~\all_features[2411] ;
  assign new_n23622_ = \all_features[2415]  & (\all_features[2414]  | (new_n23619_ & (\all_features[2410]  | \all_features[2411]  | \all_features[2409] )));
  assign new_n23623_ = \all_features[2414]  & \all_features[2415]  & (\all_features[2412]  | \all_features[2413]  | new_n23618_ | ~new_n23621_);
  assign new_n23624_ = \all_features[2415]  & (\all_features[2413]  | \all_features[2414]  | \all_features[2412] );
  assign new_n23625_ = ~new_n23626_ & (\all_features[2411]  | \all_features[2412]  | \all_features[2413]  | \all_features[2414]  | \all_features[2415] );
  assign new_n23626_ = ~\all_features[2413]  & new_n23627_ & ((~\all_features[2410]  & new_n23614_) | ~\all_features[2412]  | ~\all_features[2411] );
  assign new_n23627_ = ~\all_features[2414]  & ~\all_features[2415] ;
  assign new_n23628_ = new_n23627_ & (~\all_features[2413]  | (~\all_features[2412]  & (~\all_features[2411]  | (~\all_features[2410]  & ~\all_features[2409] ))));
  assign new_n23629_ = new_n23627_ & (~\all_features[2411]  | ~new_n23619_ | (~\all_features[2410]  & ~new_n23618_));
  assign new_n23630_ = new_n23631_ & new_n23625_ & ~new_n23628_ & ~new_n23615_;
  assign new_n23631_ = ~new_n23617_ & ~new_n23613_ & ~new_n23629_ & ~new_n23611_;
  assign new_n23632_ = new_n23625_ & (new_n23629_ | new_n23628_ | (~new_n23633_ & ~new_n23611_ & ~new_n23613_));
  assign new_n23633_ = ~new_n23615_ & ~new_n23617_ & (~new_n23624_ | ~new_n23620_ | new_n23634_);
  assign new_n23634_ = new_n23622_ & new_n23623_ & (new_n23635_ | ~\all_features[2413]  | ~\all_features[2414]  | ~\all_features[2415] );
  assign new_n23635_ = ~\all_features[2411]  & ~\all_features[2412]  & (~\all_features[2410]  | new_n23614_);
  assign new_n23636_ = ~new_n23637_ & (\all_features[2411]  | \all_features[2412]  | \all_features[2413]  | \all_features[2414]  | \all_features[2415] );
  assign new_n23637_ = ~new_n23626_ & (new_n23628_ | (~new_n23629_ & (new_n23611_ | (~new_n23638_ & ~new_n23613_))));
  assign new_n23638_ = ~new_n23615_ & (new_n23617_ | (new_n23624_ & (~new_n23620_ | (~new_n23639_ & new_n23622_))));
  assign new_n23639_ = ~\all_features[2413]  & \all_features[2414]  & \all_features[2415]  & (\all_features[2412]  ? new_n23621_ : (new_n23618_ | ~new_n23621_));
  assign new_n23640_ = ~new_n12721_ & new_n20169_;
  assign new_n23641_ = (~new_n6354_ | new_n7226_ | new_n7556_) & (new_n23640_ | ~new_n14162_ | ~new_n23642_ | ~new_n7556_);
  assign new_n23642_ = new_n22372_ & (new_n13335_ | (~new_n13343_ & (new_n13339_ | new_n23643_)));
  assign new_n23643_ = ~new_n13337_ & (new_n13342_ | (~new_n13345_ & (new_n13340_ | (~new_n13331_ & ~new_n23644_))));
  assign new_n23644_ = ~new_n23645_ & \all_features[1735]  & (\all_features[1734]  | \all_features[1733]  | \all_features[1732] );
  assign new_n23645_ = \all_features[1735]  & ((~new_n23646_ & ~\all_features[1733]  & \all_features[1734] ) | (~new_n21581_ & (\all_features[1734]  | (~new_n21576_ & \all_features[1733] ))));
  assign new_n23646_ = (\all_features[1732]  & ~new_n21577_) | (~new_n13332_ & ~\all_features[1732]  & new_n21577_);
  assign new_n23647_ = (new_n7556_ | ~new_n7226_ | ~new_n6354_ | ~new_n23654_) & (new_n16026_ | ~new_n23648_);
  assign new_n23648_ = new_n23649_ & ~new_n14162_ & new_n7556_;
  assign new_n23649_ = new_n19350_ & (new_n19374_ | (~new_n19372_ & (new_n19376_ | new_n23650_)));
  assign new_n23650_ = ~new_n19375_ & (new_n19368_ | (~new_n19369_ & (new_n19364_ | (~new_n19366_ & ~new_n23651_))));
  assign new_n23651_ = ~new_n23652_ & \all_features[2215]  & (\all_features[2214]  | \all_features[2213]  | \all_features[2212] );
  assign new_n23652_ = \all_features[2215]  & ((~new_n23653_ & ~\all_features[2213]  & \all_features[2214] ) | (~new_n19359_ & (\all_features[2214]  | (~new_n19353_ & \all_features[2213] ))));
  assign new_n23653_ = (\all_features[2212]  & ~new_n19355_) | (~new_n19362_ & ~\all_features[2212]  & new_n19355_);
  assign new_n23654_ = new_n8225_ & (new_n8202_ | ~new_n12191_);
  assign new_n23655_ = new_n23648_ & new_n16026_;
  assign new_n23656_ = new_n23657_ & (new_n7556_ | ((new_n23654_ | ~new_n7226_ | ~new_n6354_) & (~new_n23604_ | new_n6354_)));
  assign new_n23657_ = ~new_n7556_ | ((new_n23640_ | new_n23642_ | ~new_n14162_) & (new_n23123_ | new_n23649_ | new_n14162_));
  assign new_n23658_ = new_n7556_ & new_n23123_ & ~new_n14162_ & ~new_n23649_;
  assign new_n23659_ = ~new_n23772_ & new_n23660_;
  assign new_n23660_ = new_n23661_ & (new_n23770_ | new_n23649_ | new_n12082_) & (~new_n14690_ | new_n23699_ | ~new_n12082_);
  assign new_n23661_ = (~new_n23664_ | ~new_n23663_) & (~new_n23662_ | (new_n6533_ ? new_n18121_ : ~new_n23665_));
  assign new_n23662_ = ~new_n12082_ & new_n23649_;
  assign new_n23663_ = ~new_n14690_ & new_n12082_;
  assign new_n23664_ = ~new_n16102_ & ~new_n11338_;
  assign new_n23665_ = new_n23666_ & (new_n23689_ | (~new_n23696_ & ~new_n23687_));
  assign new_n23666_ = ~new_n23685_ & (~new_n23686_ | (~new_n23667_ & ~new_n23692_ & ~new_n23691_ & new_n23693_));
  assign new_n23667_ = ~new_n23679_ & ~new_n23681_ & (new_n23684_ | new_n23682_ | new_n23668_);
  assign new_n23668_ = new_n23678_ & ~new_n23672_ & new_n23669_;
  assign new_n23669_ = \all_features[1759]  & (\all_features[1758]  | new_n23670_);
  assign new_n23670_ = \all_features[1757]  & (\all_features[1754]  | \all_features[1755]  | \all_features[1756]  | ~new_n23671_);
  assign new_n23671_ = ~\all_features[1752]  & ~\all_features[1753] ;
  assign new_n23672_ = ~new_n23675_ & new_n23673_ & \all_features[1758]  & \all_features[1759]  & (~\all_features[1757]  | new_n23677_);
  assign new_n23673_ = \all_features[1759]  & (\all_features[1758]  | (new_n23674_ & (\all_features[1754]  | \all_features[1755]  | \all_features[1753] )));
  assign new_n23674_ = \all_features[1756]  & \all_features[1757] ;
  assign new_n23675_ = ~\all_features[1757]  & ~\all_features[1756]  & ~\all_features[1755]  & ~new_n23676_ & ~\all_features[1754] ;
  assign new_n23676_ = \all_features[1752]  & \all_features[1753] ;
  assign new_n23677_ = ~\all_features[1755]  & ~\all_features[1756]  & (~\all_features[1754]  | new_n23671_);
  assign new_n23678_ = \all_features[1759]  & (\all_features[1757]  | \all_features[1758]  | \all_features[1756] );
  assign new_n23679_ = ~\all_features[1759]  & (~\all_features[1758]  | (~\all_features[1756]  & ~\all_features[1757]  & ~new_n23680_));
  assign new_n23680_ = \all_features[1754]  & \all_features[1755] ;
  assign new_n23681_ = ~\all_features[1759]  & (~\all_features[1758]  | (~\all_features[1757]  & (new_n23671_ | ~new_n23680_ | ~\all_features[1756] )));
  assign new_n23682_ = ~new_n23683_ & ~\all_features[1759] ;
  assign new_n23683_ = \all_features[1757]  & \all_features[1758]  & (\all_features[1756]  | (\all_features[1754]  & \all_features[1755]  & \all_features[1753] ));
  assign new_n23684_ = ~\all_features[1759]  & (~\all_features[1758]  | ~new_n23676_ | ~new_n23674_ | ~new_n23680_);
  assign new_n23685_ = new_n23690_ & new_n23686_ & ~new_n23692_ & ~new_n23682_;
  assign new_n23686_ = ~new_n23687_ & ~new_n23689_;
  assign new_n23687_ = ~\all_features[1757]  & new_n23688_ & ((~\all_features[1754]  & new_n23671_) | ~\all_features[1756]  | ~\all_features[1755] );
  assign new_n23688_ = ~\all_features[1758]  & ~\all_features[1759] ;
  assign new_n23689_ = ~\all_features[1759]  & ~\all_features[1758]  & ~\all_features[1757]  & ~\all_features[1755]  & ~\all_features[1756] ;
  assign new_n23690_ = ~new_n23684_ & ~new_n23681_ & ~new_n23691_ & ~new_n23679_;
  assign new_n23691_ = new_n23688_ & (~\all_features[1755]  | ~new_n23674_ | (~\all_features[1754]  & ~new_n23676_));
  assign new_n23692_ = new_n23688_ & (~\all_features[1757]  | (~\all_features[1756]  & (~\all_features[1755]  | (~\all_features[1754]  & ~\all_features[1753] ))));
  assign new_n23693_ = new_n23695_ & (~new_n23673_ | ~new_n23678_ | ~new_n23694_ | ~new_n23669_);
  assign new_n23694_ = \all_features[1759]  & ~new_n23675_ & \all_features[1758] ;
  assign new_n23695_ = ~new_n23684_ & ~new_n23682_ & ~new_n23679_ & ~new_n23681_;
  assign new_n23696_ = ~new_n23692_ & (new_n23691_ | (~new_n23679_ & (new_n23681_ | (~new_n23697_ & ~new_n23682_))));
  assign new_n23697_ = ~new_n23684_ & (~new_n23678_ | (new_n23669_ & (~new_n23673_ | (~new_n23698_ & new_n23694_))));
  assign new_n23698_ = \all_features[1758]  & \all_features[1759]  & (\all_features[1757]  | (\all_features[1756]  & (\all_features[1755]  | \all_features[1754] )));
  assign new_n23699_ = new_n23735_ ? ~new_n23700_ : new_n23592_;
  assign new_n23700_ = new_n23701_ & (new_n23726_ | (~new_n23732_ & ~new_n23725_));
  assign new_n23701_ = new_n23702_ & (~new_n23724_ | (~new_n23728_ & ~new_n23727_ & ~new_n23722_));
  assign new_n23702_ = new_n23727_ | ~new_n23724_ | ((new_n23718_ | ~new_n23721_) & (new_n23703_ | new_n23722_));
  assign new_n23703_ = ~new_n23718_ & ~new_n23720_ & new_n23711_ & (~new_n23715_ | ~new_n23704_);
  assign new_n23704_ = new_n23710_ & new_n23705_ & new_n23708_;
  assign new_n23705_ = \all_features[2439]  & ~new_n23706_ & \all_features[2438] ;
  assign new_n23706_ = ~\all_features[2437]  & ~\all_features[2436]  & ~\all_features[2435]  & ~new_n23707_ & ~\all_features[2434] ;
  assign new_n23707_ = \all_features[2432]  & \all_features[2433] ;
  assign new_n23708_ = \all_features[2439]  & (\all_features[2438]  | (new_n23709_ & (\all_features[2434]  | \all_features[2435]  | \all_features[2433] )));
  assign new_n23709_ = \all_features[2436]  & \all_features[2437] ;
  assign new_n23710_ = \all_features[2439]  & (\all_features[2437]  | \all_features[2438]  | \all_features[2436] );
  assign new_n23711_ = ~new_n23712_ & ~new_n23714_;
  assign new_n23712_ = ~\all_features[2439]  & (~\all_features[2438]  | ~new_n23713_ | ~new_n23707_ | ~new_n23709_);
  assign new_n23713_ = \all_features[2434]  & \all_features[2435] ;
  assign new_n23714_ = ~\all_features[2439]  & (~\all_features[2438]  | (~\all_features[2436]  & ~\all_features[2437]  & ~new_n23713_));
  assign new_n23715_ = \all_features[2439]  & (\all_features[2438]  | new_n23716_);
  assign new_n23716_ = \all_features[2437]  & (\all_features[2434]  | \all_features[2435]  | \all_features[2436]  | ~new_n23717_);
  assign new_n23717_ = ~\all_features[2432]  & ~\all_features[2433] ;
  assign new_n23718_ = ~new_n23719_ & ~\all_features[2439] ;
  assign new_n23719_ = \all_features[2437]  & \all_features[2438]  & (\all_features[2436]  | (\all_features[2434]  & \all_features[2435]  & \all_features[2433] ));
  assign new_n23720_ = ~\all_features[2439]  & (~\all_features[2438]  | (~\all_features[2437]  & (new_n23717_ | ~new_n23713_ | ~\all_features[2436] )));
  assign new_n23721_ = new_n23711_ & ~new_n23720_ & ~new_n23722_;
  assign new_n23722_ = new_n23723_ & (~\all_features[2435]  | ~new_n23709_ | (~\all_features[2434]  & ~new_n23707_));
  assign new_n23723_ = ~\all_features[2438]  & ~\all_features[2439] ;
  assign new_n23724_ = ~new_n23725_ & ~new_n23726_;
  assign new_n23725_ = ~\all_features[2437]  & new_n23723_ & ((~\all_features[2434]  & new_n23717_) | ~\all_features[2436]  | ~\all_features[2435] );
  assign new_n23726_ = ~\all_features[2439]  & ~\all_features[2438]  & ~\all_features[2437]  & ~\all_features[2435]  & ~\all_features[2436] ;
  assign new_n23727_ = new_n23723_ & (~\all_features[2437]  | (~\all_features[2436]  & (~\all_features[2435]  | (~\all_features[2434]  & ~\all_features[2433] ))));
  assign new_n23728_ = ~new_n23720_ & ~new_n23714_ & (new_n23712_ | new_n23718_ | new_n23729_);
  assign new_n23729_ = new_n23710_ & ~new_n23730_ & new_n23715_;
  assign new_n23730_ = ~new_n23706_ & new_n23708_ & \all_features[2438]  & \all_features[2439]  & (~\all_features[2437]  | new_n23731_);
  assign new_n23731_ = ~\all_features[2435]  & ~\all_features[2436]  & (~\all_features[2434]  | new_n23717_);
  assign new_n23732_ = ~new_n23727_ & (new_n23722_ | (~new_n23714_ & (new_n23720_ | (~new_n23718_ & ~new_n23733_))));
  assign new_n23733_ = ~new_n23712_ & (~new_n23710_ | (new_n23715_ & (~new_n23708_ | (~new_n23734_ & new_n23705_))));
  assign new_n23734_ = \all_features[2438]  & \all_features[2439]  & (\all_features[2437]  | (\all_features[2436]  & (\all_features[2435]  | \all_features[2434] )));
  assign new_n23735_ = new_n23736_ & new_n23765_;
  assign new_n23736_ = ~new_n23737_ & ~new_n23761_;
  assign new_n23737_ = new_n23758_ & (~new_n23752_ | (~new_n23738_ & ~new_n23756_ & ~new_n23760_));
  assign new_n23738_ = ~new_n23749_ & ~new_n23748_ & (~new_n23751_ | ~new_n23747_ | new_n23739_);
  assign new_n23739_ = new_n23740_ & new_n23742_ & (new_n23745_ | ~\all_features[1741]  | ~\all_features[1742]  | ~\all_features[1743] );
  assign new_n23740_ = \all_features[1743]  & (\all_features[1742]  | (new_n23741_ & (\all_features[1738]  | \all_features[1739]  | \all_features[1737] )));
  assign new_n23741_ = \all_features[1740]  & \all_features[1741] ;
  assign new_n23742_ = \all_features[1742]  & \all_features[1743]  & (\all_features[1740]  | \all_features[1741]  | new_n23743_ | ~new_n23744_);
  assign new_n23743_ = \all_features[1736]  & \all_features[1737] ;
  assign new_n23744_ = ~\all_features[1738]  & ~\all_features[1739] ;
  assign new_n23745_ = ~\all_features[1739]  & ~\all_features[1740]  & (~\all_features[1738]  | new_n23746_);
  assign new_n23746_ = ~\all_features[1736]  & ~\all_features[1737] ;
  assign new_n23747_ = \all_features[1743]  & (\all_features[1742]  | (\all_features[1741]  & (\all_features[1740]  | ~new_n23746_ | ~new_n23744_)));
  assign new_n23748_ = ~\all_features[1743]  & (~new_n23741_ | ~\all_features[1738]  | ~\all_features[1739]  | ~\all_features[1742]  | ~new_n23743_);
  assign new_n23749_ = ~new_n23750_ & ~\all_features[1743] ;
  assign new_n23750_ = \all_features[1741]  & \all_features[1742]  & (\all_features[1740]  | (\all_features[1738]  & \all_features[1739]  & \all_features[1737] ));
  assign new_n23751_ = \all_features[1743]  & (\all_features[1741]  | \all_features[1742]  | \all_features[1740] );
  assign new_n23752_ = ~new_n23753_ & ~new_n23755_;
  assign new_n23753_ = new_n23754_ & (~\all_features[1739]  | ~new_n23741_ | (~\all_features[1738]  & ~new_n23743_));
  assign new_n23754_ = ~\all_features[1742]  & ~\all_features[1743] ;
  assign new_n23755_ = new_n23754_ & (~\all_features[1741]  | (~\all_features[1740]  & (~\all_features[1739]  | (~\all_features[1738]  & ~\all_features[1737] ))));
  assign new_n23756_ = ~\all_features[1743]  & (~\all_features[1742]  | new_n23757_);
  assign new_n23757_ = ~\all_features[1741]  & (new_n23746_ | ~\all_features[1739]  | ~\all_features[1740]  | ~\all_features[1738] );
  assign new_n23758_ = ~new_n23759_ & (\all_features[1739]  | \all_features[1740]  | \all_features[1741]  | \all_features[1742]  | \all_features[1743] );
  assign new_n23759_ = ~\all_features[1741]  & new_n23754_ & ((~\all_features[1738]  & new_n23746_) | ~\all_features[1740]  | ~\all_features[1739] );
  assign new_n23760_ = ~\all_features[1743]  & (~\all_features[1742]  | (~\all_features[1741]  & ~\all_features[1740]  & (~\all_features[1739]  | ~\all_features[1738] )));
  assign new_n23761_ = ~new_n23762_ & (\all_features[1739]  | \all_features[1740]  | \all_features[1741]  | \all_features[1742]  | \all_features[1743] );
  assign new_n23762_ = ~new_n23759_ & (new_n23755_ | (~new_n23753_ & (new_n23760_ | (~new_n23756_ & ~new_n23763_))));
  assign new_n23763_ = ~new_n23749_ & (new_n23748_ | (new_n23751_ & (~new_n23747_ | (~new_n23764_ & new_n23740_))));
  assign new_n23764_ = ~\all_features[1741]  & \all_features[1742]  & \all_features[1743]  & (\all_features[1740]  ? new_n23744_ : (new_n23743_ | ~new_n23744_));
  assign new_n23765_ = ~new_n23766_ & ~new_n23769_;
  assign new_n23766_ = new_n23752_ & new_n23758_ & (new_n23756_ | new_n23767_ | new_n23748_ | ~new_n23768_);
  assign new_n23767_ = new_n23751_ & new_n23747_ & new_n23740_ & new_n23742_;
  assign new_n23768_ = ~new_n23749_ & ~new_n23760_;
  assign new_n23769_ = new_n23752_ & new_n23768_ & new_n23758_ & ~new_n23756_ & ~new_n23748_;
  assign new_n23770_ = new_n12849_ ? new_n23771_ : new_n14290_;
  assign new_n23771_ = ~new_n20098_ & new_n19237_;
  assign new_n23772_ = (~new_n23663_ | new_n23664_) & (~new_n23662_ | (new_n6533_ ? ~new_n18121_ : new_n23665_));
  assign new_n23773_ = new_n23774_ ? (new_n23828_ ^ new_n23883_) : (~new_n23828_ ^ new_n23883_);
  assign new_n23774_ = ~new_n23775_ & new_n23824_;
  assign new_n23775_ = ~new_n23783_ & new_n23776_ & (~new_n23820_ | (new_n23823_ & new_n12264_) | (~new_n23822_ & ~new_n12264_));
  assign new_n23776_ = ~new_n10000_ | ((~new_n23777_ | ~new_n23779_) & (new_n23782_ | ~new_n23780_ | new_n23779_));
  assign new_n23777_ = new_n23778_ & ~new_n20156_ & ~new_n17176_;
  assign new_n23778_ = new_n12048_ & new_n12081_;
  assign new_n23779_ = ~new_n22458_ & new_n15477_;
  assign new_n23780_ = ~new_n10562_ & new_n23781_;
  assign new_n23781_ = ~new_n10540_ & ~new_n10569_;
  assign new_n23782_ = ~new_n20662_ & ~new_n20693_;
  assign new_n23783_ = new_n10000_ & ((~new_n23778_ & new_n23784_ & new_n23779_) | (new_n15867_ & new_n23782_ & ~new_n23779_));
  assign new_n23784_ = ~new_n23785_ & new_n23814_;
  assign new_n23785_ = ~new_n23786_ & ~new_n23810_;
  assign new_n23786_ = new_n23801_ & (~new_n23806_ | (~new_n23804_ & ~new_n23787_ & ~new_n23809_));
  assign new_n23787_ = ~new_n23799_ & ~new_n23797_ & (~new_n23800_ | ~new_n23796_ | new_n23788_);
  assign new_n23788_ = new_n23789_ & new_n23791_ & (new_n23794_ | ~\all_features[5493]  | ~\all_features[5494]  | ~\all_features[5495] );
  assign new_n23789_ = \all_features[5495]  & (\all_features[5494]  | (new_n23790_ & (\all_features[5490]  | \all_features[5491]  | \all_features[5489] )));
  assign new_n23790_ = \all_features[5492]  & \all_features[5493] ;
  assign new_n23791_ = \all_features[5494]  & \all_features[5495]  & (\all_features[5492]  | \all_features[5493]  | new_n23793_ | ~new_n23792_);
  assign new_n23792_ = ~\all_features[5490]  & ~\all_features[5491] ;
  assign new_n23793_ = \all_features[5488]  & \all_features[5489] ;
  assign new_n23794_ = ~\all_features[5491]  & ~\all_features[5492]  & (~\all_features[5490]  | new_n23795_);
  assign new_n23795_ = ~\all_features[5488]  & ~\all_features[5489] ;
  assign new_n23796_ = \all_features[5495]  & (\all_features[5494]  | (\all_features[5493]  & (\all_features[5492]  | ~new_n23792_ | ~new_n23795_)));
  assign new_n23797_ = ~new_n23798_ & ~\all_features[5495] ;
  assign new_n23798_ = \all_features[5493]  & \all_features[5494]  & (\all_features[5492]  | (\all_features[5490]  & \all_features[5491]  & \all_features[5489] ));
  assign new_n23799_ = ~\all_features[5495]  & (~new_n23793_ | ~\all_features[5490]  | ~\all_features[5491]  | ~\all_features[5494]  | ~new_n23790_);
  assign new_n23800_ = \all_features[5495]  & (\all_features[5493]  | \all_features[5494]  | \all_features[5492] );
  assign new_n23801_ = ~new_n23802_ & (\all_features[5491]  | \all_features[5492]  | \all_features[5493]  | \all_features[5494]  | \all_features[5495] );
  assign new_n23802_ = ~\all_features[5493]  & new_n23803_ & ((~\all_features[5490]  & new_n23795_) | ~\all_features[5492]  | ~\all_features[5491] );
  assign new_n23803_ = ~\all_features[5494]  & ~\all_features[5495] ;
  assign new_n23804_ = ~\all_features[5495]  & (~\all_features[5494]  | new_n23805_);
  assign new_n23805_ = ~\all_features[5493]  & (new_n23795_ | ~\all_features[5491]  | ~\all_features[5492]  | ~\all_features[5490] );
  assign new_n23806_ = ~new_n23807_ & ~new_n23808_;
  assign new_n23807_ = new_n23803_ & (~\all_features[5493]  | (~\all_features[5492]  & (~\all_features[5491]  | (~\all_features[5490]  & ~\all_features[5489] ))));
  assign new_n23808_ = new_n23803_ & (~\all_features[5491]  | ~new_n23790_ | (~new_n23793_ & ~\all_features[5490] ));
  assign new_n23809_ = ~\all_features[5495]  & (~\all_features[5494]  | (~\all_features[5493]  & ~\all_features[5492]  & (~\all_features[5491]  | ~\all_features[5490] )));
  assign new_n23810_ = ~new_n23811_ & (\all_features[5491]  | \all_features[5492]  | \all_features[5493]  | \all_features[5494]  | \all_features[5495] );
  assign new_n23811_ = ~new_n23802_ & (new_n23807_ | (~new_n23808_ & (new_n23809_ | (~new_n23804_ & ~new_n23812_))));
  assign new_n23812_ = ~new_n23797_ & (new_n23799_ | (new_n23800_ & (~new_n23796_ | (~new_n23813_ & new_n23789_))));
  assign new_n23813_ = ~\all_features[5493]  & \all_features[5494]  & \all_features[5495]  & (\all_features[5492]  ? new_n23792_ : (new_n23793_ | ~new_n23792_));
  assign new_n23814_ = new_n23815_ & new_n23818_;
  assign new_n23815_ = new_n23806_ & ~new_n23816_ & new_n23801_;
  assign new_n23816_ = ~new_n23809_ & ~new_n23799_ & ~new_n23797_ & ~new_n23804_ & ~new_n23817_;
  assign new_n23817_ = new_n23800_ & new_n23796_ & new_n23789_ & new_n23791_;
  assign new_n23818_ = new_n23801_ & new_n23819_ & ~new_n23797_ & ~new_n23807_;
  assign new_n23819_ = ~new_n23809_ & ~new_n23808_ & ~new_n23804_ & ~new_n23799_;
  assign new_n23820_ = ~new_n10000_ & new_n23821_;
  assign new_n23821_ = ~new_n8704_ & new_n21530_;
  assign new_n23822_ = ~new_n15916_ & new_n11094_;
  assign new_n23823_ = new_n23558_ & new_n23581_;
  assign new_n23824_ = ~new_n23825_ & new_n23826_ & (new_n23822_ | new_n12264_ | ~new_n23820_);
  assign new_n23825_ = ~new_n23777_ & new_n10000_ & new_n23779_ & (~new_n23784_ | new_n23778_);
  assign new_n23826_ = (new_n23779_ | new_n23827_ | ~new_n10000_) & (new_n23821_ | new_n10000_ | (~new_n18324_ & ~new_n23702_));
  assign new_n23827_ = new_n23782_ ? new_n15867_ : new_n23780_;
  assign new_n23828_ = ~new_n23829_ & new_n23881_;
  assign new_n23829_ = new_n23875_ & new_n23830_ & (new_n23880_ | new_n23878_ | ~new_n23877_);
  assign new_n23830_ = (new_n23868_ | ~new_n23831_) & (~new_n14046_ | ~new_n23832_ | new_n23869_ | new_n14211_);
  assign new_n23831_ = ~new_n23867_ & ~new_n23832_ & ~new_n22998_;
  assign new_n23832_ = ~new_n23863_ & new_n23833_;
  assign new_n23833_ = ~new_n23859_ & new_n23834_;
  assign new_n23834_ = ~new_n23835_ & ~new_n23857_;
  assign new_n23835_ = new_n23852_ & ~new_n23856_ & ~new_n23836_ & ~new_n23855_;
  assign new_n23836_ = new_n23837_ & (~new_n23850_ | ~new_n23851_ | ~new_n23847_ | ~new_n23849_);
  assign new_n23837_ = ~new_n23844_ & ~new_n23842_ & ~new_n23838_ & ~new_n23840_;
  assign new_n23838_ = ~\all_features[831]  & (~\all_features[830]  | (~\all_features[828]  & ~\all_features[829]  & ~new_n23839_));
  assign new_n23839_ = \all_features[826]  & \all_features[827] ;
  assign new_n23840_ = ~\all_features[831]  & (~\all_features[830]  | (~\all_features[829]  & (new_n23841_ | ~new_n23839_ | ~\all_features[828] )));
  assign new_n23841_ = ~\all_features[824]  & ~\all_features[825] ;
  assign new_n23842_ = ~new_n23843_ & ~\all_features[831] ;
  assign new_n23843_ = \all_features[829]  & \all_features[830]  & (\all_features[828]  | (\all_features[826]  & \all_features[827]  & \all_features[825] ));
  assign new_n23844_ = ~\all_features[831]  & (~\all_features[830]  | ~new_n23845_ | ~new_n23846_ | ~new_n23839_);
  assign new_n23845_ = \all_features[824]  & \all_features[825] ;
  assign new_n23846_ = \all_features[828]  & \all_features[829] ;
  assign new_n23847_ = \all_features[831]  & (\all_features[830]  | (\all_features[829]  & (\all_features[828]  | ~new_n23848_ | ~new_n23841_)));
  assign new_n23848_ = ~\all_features[826]  & ~\all_features[827] ;
  assign new_n23849_ = \all_features[831]  & (\all_features[830]  | (new_n23846_ & (\all_features[826]  | \all_features[827]  | \all_features[825] )));
  assign new_n23850_ = \all_features[830]  & \all_features[831]  & (\all_features[828]  | \all_features[829]  | new_n23845_ | ~new_n23848_);
  assign new_n23851_ = \all_features[831]  & (\all_features[829]  | \all_features[830]  | \all_features[828] );
  assign new_n23852_ = ~new_n23853_ & (\all_features[827]  | \all_features[828]  | \all_features[829]  | \all_features[830]  | \all_features[831] );
  assign new_n23853_ = ~\all_features[829]  & new_n23854_ & ((~\all_features[826]  & new_n23841_) | ~\all_features[828]  | ~\all_features[827] );
  assign new_n23854_ = ~\all_features[830]  & ~\all_features[831] ;
  assign new_n23855_ = new_n23854_ & (~\all_features[829]  | (~\all_features[828]  & (~\all_features[827]  | (~\all_features[826]  & ~\all_features[825] ))));
  assign new_n23856_ = new_n23854_ & (~\all_features[827]  | ~new_n23846_ | (~\all_features[826]  & ~new_n23845_));
  assign new_n23857_ = new_n23858_ & new_n23852_ & ~new_n23855_ & ~new_n23842_;
  assign new_n23858_ = ~new_n23844_ & ~new_n23840_ & ~new_n23856_ & ~new_n23838_;
  assign new_n23859_ = new_n23852_ & (new_n23856_ | new_n23855_ | (~new_n23860_ & ~new_n23838_ & ~new_n23840_));
  assign new_n23860_ = ~new_n23842_ & ~new_n23844_ & (~new_n23851_ | ~new_n23847_ | new_n23861_);
  assign new_n23861_ = new_n23849_ & new_n23850_ & (new_n23862_ | ~\all_features[829]  | ~\all_features[830]  | ~\all_features[831] );
  assign new_n23862_ = ~\all_features[827]  & ~\all_features[828]  & (~\all_features[826]  | new_n23841_);
  assign new_n23863_ = ~new_n23864_ & (\all_features[827]  | \all_features[828]  | \all_features[829]  | \all_features[830]  | \all_features[831] );
  assign new_n23864_ = ~new_n23853_ & (new_n23855_ | (~new_n23856_ & (new_n23838_ | (~new_n23865_ & ~new_n23840_))));
  assign new_n23865_ = ~new_n23842_ & (new_n23844_ | (new_n23851_ & (~new_n23847_ | (~new_n23866_ & new_n23849_))));
  assign new_n23866_ = ~\all_features[829]  & \all_features[830]  & \all_features[831]  & (\all_features[828]  ? new_n23848_ : (new_n23845_ | ~new_n23848_));
  assign new_n23867_ = ~new_n21882_ & new_n21855_;
  assign new_n23868_ = ~new_n12257_ & (~new_n12254_ | ~new_n12793_);
  assign new_n23869_ = new_n23870_ & ~new_n22080_ & ~new_n22083_;
  assign new_n23870_ = ~new_n22053_ & (new_n22068_ | (~new_n22066_ & (new_n22071_ | (~new_n22070_ & ~new_n23871_))));
  assign new_n23871_ = ~new_n22073_ & (new_n22075_ | (~new_n22078_ & (new_n22077_ | (~new_n23872_ & new_n23874_))));
  assign new_n23872_ = \all_features[5231]  & ((~new_n23873_ & ~\all_features[5229]  & \all_features[5230] ) | (~new_n22060_ & (\all_features[5230]  | (~new_n22056_ & \all_features[5229] ))));
  assign new_n23873_ = (\all_features[5228]  & ~new_n22058_) | (~new_n22063_ & ~\all_features[5228]  & new_n22058_);
  assign new_n23874_ = \all_features[5231]  & (\all_features[5229]  | \all_features[5230]  | \all_features[5228] );
  assign new_n23875_ = (new_n23867_ | ~new_n22998_ | new_n23832_) & (~new_n23832_ | (new_n14046_ ? ~new_n14211_ : new_n23876_));
  assign new_n23876_ = ~new_n10271_ & ~new_n16855_ & new_n9579_ & (~new_n10273_ | ~new_n10249_);
  assign new_n23877_ = ~new_n23832_ & new_n23867_;
  assign new_n23878_ = new_n16355_ & new_n23879_;
  assign new_n23879_ = ~new_n9993_ & ~new_n9995_;
  assign new_n23880_ = ~new_n15756_ & new_n10976_;
  assign new_n23881_ = new_n23882_ & (~new_n23832_ | ((new_n14211_ | ~new_n23869_ | ~new_n14046_) & (~new_n23876_ | new_n14046_)));
  assign new_n23882_ = (~new_n23868_ | ~new_n23831_) & (~new_n23877_ | (new_n23880_ ? new_n20973_ : ~new_n23878_));
  assign new_n23883_ = ~new_n23928_ & new_n23884_;
  assign new_n23884_ = new_n23923_ & (new_n10775_ | ~new_n23920_) & (new_n21767_ | new_n23885_);
  assign new_n23885_ = (new_n23886_ | ~new_n23919_) & (new_n12727_ | ~new_n21692_ | new_n23919_);
  assign new_n23886_ = (new_n23887_ & (~new_n23911_ | ~new_n23915_)) ? ~new_n23700_ : new_n15030_;
  assign new_n23887_ = new_n23910_ | ~new_n23908_ | ((new_n23899_ | new_n23897_) & (new_n23905_ | ~new_n23888_));
  assign new_n23888_ = new_n23889_ & ~new_n23895_ & ~new_n23897_;
  assign new_n23889_ = ~new_n23890_ & ~new_n23894_;
  assign new_n23890_ = ~\all_features[1527]  & (~\all_features[1526]  | ~new_n23891_ | ~new_n23892_ | ~new_n23893_);
  assign new_n23891_ = \all_features[1522]  & \all_features[1523] ;
  assign new_n23892_ = \all_features[1520]  & \all_features[1521] ;
  assign new_n23893_ = \all_features[1524]  & \all_features[1525] ;
  assign new_n23894_ = ~\all_features[1527]  & (~\all_features[1526]  | (~\all_features[1524]  & ~\all_features[1525]  & ~new_n23891_));
  assign new_n23895_ = ~\all_features[1527]  & (~\all_features[1526]  | (~\all_features[1525]  & (new_n23896_ | ~new_n23891_ | ~\all_features[1524] )));
  assign new_n23896_ = ~\all_features[1520]  & ~\all_features[1521] ;
  assign new_n23897_ = new_n23898_ & (~\all_features[1523]  | ~new_n23893_ | (~\all_features[1522]  & ~new_n23892_));
  assign new_n23898_ = ~\all_features[1526]  & ~\all_features[1527] ;
  assign new_n23899_ = ~new_n23905_ & ~new_n23895_ & new_n23889_ & (~new_n23907_ | ~new_n23900_);
  assign new_n23900_ = new_n23904_ & new_n23901_ & new_n23902_;
  assign new_n23901_ = \all_features[1527]  & (\all_features[1526]  | (new_n23893_ & (\all_features[1522]  | \all_features[1523]  | \all_features[1521] )));
  assign new_n23902_ = \all_features[1526]  & \all_features[1527]  & (\all_features[1524]  | \all_features[1525]  | new_n23892_ | ~new_n23903_);
  assign new_n23903_ = ~\all_features[1522]  & ~\all_features[1523] ;
  assign new_n23904_ = \all_features[1527]  & (\all_features[1525]  | \all_features[1526]  | \all_features[1524] );
  assign new_n23905_ = ~new_n23906_ & ~\all_features[1527] ;
  assign new_n23906_ = \all_features[1525]  & \all_features[1526]  & (\all_features[1524]  | (\all_features[1522]  & \all_features[1523]  & \all_features[1521] ));
  assign new_n23907_ = \all_features[1527]  & (\all_features[1526]  | (\all_features[1525]  & (\all_features[1524]  | ~new_n23903_ | ~new_n23896_)));
  assign new_n23908_ = ~new_n23909_ & (\all_features[1523]  | \all_features[1524]  | \all_features[1525]  | \all_features[1526]  | \all_features[1527] );
  assign new_n23909_ = ~\all_features[1525]  & new_n23898_ & ((~\all_features[1522]  & new_n23896_) | ~\all_features[1524]  | ~\all_features[1523] );
  assign new_n23910_ = new_n23898_ & (~\all_features[1525]  | (~\all_features[1524]  & (~\all_features[1523]  | (~\all_features[1522]  & ~\all_features[1521] ))));
  assign new_n23911_ = new_n23908_ & (new_n23897_ | new_n23910_ | (~new_n23912_ & ~new_n23895_ & ~new_n23894_));
  assign new_n23912_ = ~new_n23905_ & ~new_n23890_ & (~new_n23904_ | ~new_n23907_ | new_n23913_);
  assign new_n23913_ = new_n23901_ & new_n23902_ & (new_n23914_ | ~\all_features[1525]  | ~\all_features[1526]  | ~\all_features[1527] );
  assign new_n23914_ = ~\all_features[1523]  & ~\all_features[1524]  & (~\all_features[1522]  | new_n23896_);
  assign new_n23915_ = ~new_n23916_ & (\all_features[1523]  | \all_features[1524]  | \all_features[1525]  | \all_features[1526]  | \all_features[1527] );
  assign new_n23916_ = ~new_n23909_ & (new_n23910_ | (~new_n23897_ & (new_n23894_ | (~new_n23895_ & ~new_n23917_))));
  assign new_n23917_ = ~new_n23905_ & (new_n23890_ | (new_n23904_ & (~new_n23907_ | (~new_n23918_ & new_n23901_))));
  assign new_n23918_ = ~\all_features[1525]  & \all_features[1526]  & \all_features[1527]  & (\all_features[1524]  ? new_n23903_ : (new_n23892_ | ~new_n23903_));
  assign new_n23919_ = new_n23140_ & ~new_n17857_ & ~new_n17877_;
  assign new_n23920_ = new_n21767_ & ~new_n23921_ & ~new_n23922_;
  assign new_n23921_ = ~new_n7993_ & ~new_n8028_;
  assign new_n23922_ = new_n23196_ & new_n12152_;
  assign new_n23923_ = (~new_n23925_ | new_n23927_) & (~new_n23924_ | (new_n18120_ ? new_n15917_ : ~new_n23926_));
  assign new_n23924_ = new_n21767_ & new_n23922_;
  assign new_n23925_ = ~new_n23919_ & ~new_n21692_ & ~new_n21767_;
  assign new_n23926_ = ~new_n20684_ & new_n23782_;
  assign new_n23927_ = new_n13014_ & new_n17844_;
  assign new_n23928_ = ~new_n23929_ & new_n23930_ & (~new_n10775_ | ~new_n23920_);
  assign new_n23929_ = new_n21767_ & ((new_n23921_ & ~new_n23922_) | (~new_n23926_ & ~new_n18120_ & new_n23922_));
  assign new_n23930_ = (~new_n23924_ | ~new_n15917_ | ~new_n18120_) & (~new_n23927_ | ~new_n23925_);
  assign new_n23931_ = new_n23932_ & new_n23938_;
  assign new_n23932_ = new_n23933_ & (new_n23934_ | ~new_n23936_ | (new_n20405_ ? new_n23937_ : ~new_n20117_));
  assign new_n23933_ = (new_n23935_ | new_n23936_) & (~new_n23934_ | ~new_n23936_ | (new_n10947_ ? new_n12732_ : ~new_n7902_));
  assign new_n23934_ = new_n10379_ & new_n8391_;
  assign new_n23935_ = new_n17392_ & new_n17414_;
  assign new_n23936_ = ~\all_features[1103]  & (~\all_features[1102]  | (~\all_features[1101]  & (~\all_features[1100]  | ~\all_features[1099] )));
  assign new_n23937_ = new_n15664_ & new_n15660_ & new_n15632_ & new_n15656_;
  assign new_n23938_ = ~new_n23936_ | (new_n23934_ ? new_n23939_ : (new_n20405_ ? ~new_n23937_ : new_n20117_));
  assign new_n23939_ = new_n10947_ ? ~new_n12732_ : new_n7902_;
  assign new_n23940_ = new_n23941_ ? (~new_n23931_ ^ new_n24036_) : (new_n23931_ ^ new_n24036_);
  assign new_n23941_ = new_n23942_ ? (new_n23958_ ^ new_n24003_) : (~new_n23958_ ^ new_n24003_);
  assign new_n23942_ = ~new_n23943_ & new_n23956_;
  assign new_n23943_ = new_n23944_ & (~new_n23832_ | ~new_n23954_ | ~new_n20923_);
  assign new_n23944_ = ~new_n23945_ & (new_n23832_ | ~new_n23953_ | (new_n15672_ ? new_n11668_ : new_n12908_));
  assign new_n23945_ = new_n23832_ & ~new_n20923_ & ~new_n23946_;
  assign new_n23946_ = new_n23947_ & new_n14495_ & (~new_n23948_ | (new_n22501_ & new_n23949_));
  assign new_n23947_ = new_n14471_ & new_n14493_;
  assign new_n23948_ = ~new_n22528_ & ~new_n22530_;
  assign new_n23949_ = ~new_n22521_ & (new_n22519_ | new_n23950_);
  assign new_n23950_ = ~new_n22523_ & (new_n22524_ | (~new_n22526_ & (new_n22527_ | (~new_n23951_ & ~new_n22504_))));
  assign new_n23951_ = ~new_n22506_ & (~new_n22517_ | (new_n22516_ & (~new_n22513_ | (~new_n23952_ & new_n22514_))));
  assign new_n23952_ = \all_features[2422]  & \all_features[2423]  & (\all_features[2421]  | (~new_n22515_ & \all_features[2420] ));
  assign new_n23953_ = ~new_n10761_ & (~new_n10767_ | ~new_n10739_);
  assign new_n23954_ = new_n11060_ & (~new_n12354_ | (~new_n23955_ & ~new_n14164_));
  assign new_n23955_ = new_n14173_ & new_n14177_;
  assign new_n23956_ = new_n23832_ ? (new_n20923_ ? new_n23954_ : ~new_n23946_) : new_n23957_;
  assign new_n23957_ = new_n23953_ & (new_n15672_ | ~new_n12908_);
  assign new_n23958_ = ~new_n23959_ & new_n23999_;
  assign new_n23959_ = new_n23960_ & (new_n23963_ | (~new_n23970_ & (new_n19342_ | ~new_n13846_ | ~new_n23971_)));
  assign new_n23960_ = ~new_n23961_ & (~new_n23963_ | (~new_n23965_ & new_n21207_) | (~new_n23967_ & ~new_n23969_ & ~new_n21207_));
  assign new_n23961_ = new_n23962_ & new_n11905_;
  assign new_n23962_ = ~new_n23963_ & ~new_n13846_ & ~new_n19342_;
  assign new_n23963_ = new_n22645_ & new_n23964_;
  assign new_n23964_ = ~new_n15763_ & ~new_n15786_;
  assign new_n23965_ = ~new_n23966_ & (~new_n11699_ | (~new_n11675_ & new_n13203_));
  assign new_n23966_ = new_n12398_ & (new_n12376_ | ~new_n12731_);
  assign new_n23967_ = ~new_n11857_ & new_n23968_;
  assign new_n23968_ = ~new_n11846_ & ~new_n11854_;
  assign new_n23969_ = new_n15082_ & new_n15050_ & new_n15079_;
  assign new_n23970_ = ~new_n14119_ & new_n16757_ & new_n19342_ & (~new_n14122_ | new_n14090_);
  assign new_n23971_ = new_n23998_ | (~new_n23990_ & new_n23972_);
  assign new_n23972_ = new_n23990_ & (new_n23994_ | (~new_n23995_ & new_n23973_ & (new_n23982_ | new_n23988_)));
  assign new_n23973_ = ~new_n23982_ & ~new_n23984_ & (~new_n23987_ | ~new_n23986_ | new_n23974_);
  assign new_n23974_ = new_n23975_ & ~new_n23980_ & new_n23977_;
  assign new_n23975_ = \all_features[3855]  & (\all_features[3854]  | (new_n23976_ & (\all_features[3850]  | \all_features[3851]  | \all_features[3849] )));
  assign new_n23976_ = \all_features[3852]  & \all_features[3853] ;
  assign new_n23977_ = new_n23979_ & (\all_features[3852]  | \all_features[3853]  | ~new_n23978_ | (\all_features[3849]  & \all_features[3848] ));
  assign new_n23978_ = ~\all_features[3850]  & ~\all_features[3851] ;
  assign new_n23979_ = \all_features[3854]  & \all_features[3855] ;
  assign new_n23980_ = new_n23979_ & \all_features[3853]  & ((~new_n23981_ & \all_features[3850] ) | \all_features[3852]  | \all_features[3851] );
  assign new_n23981_ = ~\all_features[3848]  & ~\all_features[3849] ;
  assign new_n23982_ = ~new_n23983_ & ~\all_features[3855] ;
  assign new_n23983_ = \all_features[3853]  & \all_features[3854]  & (\all_features[3852]  | (\all_features[3850]  & \all_features[3851]  & \all_features[3849] ));
  assign new_n23984_ = ~\all_features[3855]  & (~new_n23976_ | ~\all_features[3848]  | ~\all_features[3849]  | ~\all_features[3854]  | ~new_n23985_);
  assign new_n23985_ = \all_features[3850]  & \all_features[3851] ;
  assign new_n23986_ = \all_features[3855]  & (\all_features[3854]  | (\all_features[3853]  & (\all_features[3852]  | ~new_n23978_ | ~new_n23981_)));
  assign new_n23987_ = \all_features[3855]  & (\all_features[3853]  | \all_features[3854]  | \all_features[3852] );
  assign new_n23988_ = ~new_n23984_ & (~new_n23987_ | (new_n23986_ & (~new_n23975_ | (~new_n23989_ & new_n23977_))));
  assign new_n23989_ = new_n23979_ & (\all_features[3853]  | (~new_n23978_ & \all_features[3852] ));
  assign new_n23990_ = \all_features[3854]  | \all_features[3855]  | (~new_n23993_ & new_n23991_ & \all_features[3853] );
  assign new_n23991_ = new_n23976_ & \all_features[3851]  & (\all_features[3850]  | (\all_features[3848]  & \all_features[3849] ));
  assign new_n23993_ = ~\all_features[3852]  & (~\all_features[3851]  | (~\all_features[3850]  & ~\all_features[3849] ));
  assign new_n23994_ = ~\all_features[3855]  & (~\all_features[3854]  | (~\all_features[3852]  & ~\all_features[3853]  & ~new_n23985_));
  assign new_n23995_ = ~\all_features[3855]  & (~\all_features[3854]  | (~\all_features[3853]  & (new_n23981_ | ~\all_features[3852]  | ~new_n23985_)));
  assign new_n23998_ = ~\all_features[3855]  & ~\all_features[3854]  & ~\all_features[3853]  & ~\all_features[3851]  & ~\all_features[3852] ;
  assign new_n23999_ = new_n24000_ & (new_n11905_ | ~new_n23962_);
  assign new_n24000_ = (new_n16757_ | new_n24002_ | ~new_n19342_ | new_n23963_) & (~new_n23966_ | ~new_n24001_ | ~new_n23963_);
  assign new_n24001_ = new_n21207_ & (new_n10478_ | ~new_n19150_);
  assign new_n24002_ = new_n9314_ & new_n9340_;
  assign new_n24003_ = new_n24004_ & new_n24024_;
  assign new_n24004_ = new_n24023_ | (new_n23963_ ? (new_n24005_ ? new_n9313_ : ~new_n14290_) : new_n24006_);
  assign new_n24005_ = new_n10206_ & new_n10240_;
  assign new_n24006_ = (~new_n24019_ & new_n24009_ & new_n24007_) | (new_n24008_ & new_n7188_ & ~new_n24007_);
  assign new_n24007_ = new_n10207_ & ~new_n10238_ & ~new_n10240_;
  assign new_n24008_ = new_n7164_ & new_n7192_;
  assign new_n24009_ = ~new_n24010_ & ~new_n20852_;
  assign new_n24010_ = new_n24018_ & ~new_n24011_ & new_n24017_;
  assign new_n24011_ = ~new_n20862_ & ~new_n20865_ & ~new_n20854_ & ~new_n20861_ & (~new_n24014_ | ~new_n24012_);
  assign new_n24012_ = \all_features[3527]  & (\all_features[3526]  | (~new_n24013_ & \all_features[3525] ));
  assign new_n24013_ = new_n20856_ & ~\all_features[3524]  & ~\all_features[3522]  & ~\all_features[3523] ;
  assign new_n24014_ = \all_features[3527]  & \all_features[3526]  & ~new_n24016_ & new_n24015_;
  assign new_n24015_ = \all_features[3527]  & (\all_features[3526]  | (new_n20859_ & (\all_features[3522]  | \all_features[3523]  | \all_features[3521] )));
  assign new_n24016_ = ~\all_features[3522]  & ~\all_features[3523]  & ~\all_features[3524]  & ~\all_features[3525]  & (~\all_features[3521]  | ~\all_features[3520] );
  assign new_n24017_ = ~new_n20860_ & ~new_n20866_;
  assign new_n24018_ = ~new_n20864_ & ~new_n20857_;
  assign new_n24019_ = new_n24017_ & (~new_n24018_ | (~new_n24020_ & ~new_n20854_ & ~new_n20861_));
  assign new_n24020_ = ~new_n20862_ & ~new_n20865_ & (~new_n24012_ | (~new_n24021_ & new_n24014_));
  assign new_n24021_ = \all_features[3527]  & \all_features[3526]  & ~new_n24022_ & \all_features[3525] ;
  assign new_n24022_ = ~\all_features[3523]  & ~\all_features[3524]  & (~\all_features[3522]  | new_n20856_);
  assign new_n24023_ = new_n12529_ & new_n19829_;
  assign new_n24024_ = ~new_n24023_ | (new_n24034_ ? (new_n23122_ ? new_n22531_ : new_n17214_) : new_n24025_);
  assign new_n24025_ = (~new_n22922_ & (new_n24026_ | ~new_n22899_)) ? ~new_n24033_ : new_n17933_;
  assign new_n24026_ = ~new_n24027_ & ~new_n22923_;
  assign new_n24027_ = ~new_n24028_ & (\all_features[3299]  | \all_features[3300]  | ~new_n22903_);
  assign new_n24028_ = ~new_n22902_ & (new_n22908_ | (~new_n22906_ & (new_n22919_ | new_n24029_)));
  assign new_n24029_ = ~new_n22917_ & (new_n22913_ | (~new_n22915_ & (~new_n24032_ | new_n24030_)));
  assign new_n24030_ = \all_features[3303]  & ((~new_n24031_ & ~\all_features[3301]  & \all_features[3302] ) | (~new_n22910_ & (\all_features[3302]  | (~new_n22921_ & \all_features[3301] ))));
  assign new_n24031_ = (~\all_features[3298]  & ~\all_features[3299]  & ~\all_features[3300]  & (~\all_features[3297]  | ~\all_features[3296] )) | (\all_features[3300]  & (\all_features[3298]  | \all_features[3299] ));
  assign new_n24032_ = \all_features[3303]  & (\all_features[3301]  | \all_features[3302]  | \all_features[3300] );
  assign new_n24033_ = ~new_n23584_ & new_n23557_;
  assign new_n24034_ = ~new_n22423_ & (~new_n22420_ | ~new_n24035_);
  assign new_n24035_ = new_n22391_ & new_n22415_;
  assign new_n24036_ = ~new_n24113_ & new_n24037_;
  assign new_n24037_ = new_n24076_ ? ~new_n24038_ : ((new_n22386_ & ~new_n24077_) | (new_n23557_ & new_n24112_ & new_n24077_));
  assign new_n24038_ = new_n24041_ & ~new_n24039_ & new_n21615_;
  assign new_n24039_ = new_n24040_ & new_n11369_;
  assign new_n24040_ = new_n20308_ & new_n11365_;
  assign new_n24041_ = ~new_n24072_ & new_n24042_;
  assign new_n24042_ = ~new_n24043_ & new_n24067_;
  assign new_n24043_ = new_n24059_ & (~new_n24062_ | (~new_n24044_ & ~new_n24065_ & ~new_n24066_));
  assign new_n24044_ = ~new_n24053_ & ~new_n24055_ & (~new_n24058_ | ~new_n24057_ | new_n24045_);
  assign new_n24045_ = new_n24046_ & new_n24048_ & (new_n24051_ | ~\all_features[1277]  | ~\all_features[1278]  | ~\all_features[1279] );
  assign new_n24046_ = \all_features[1279]  & (\all_features[1278]  | (new_n24047_ & (\all_features[1274]  | \all_features[1275]  | \all_features[1273] )));
  assign new_n24047_ = \all_features[1276]  & \all_features[1277] ;
  assign new_n24048_ = \all_features[1278]  & \all_features[1279]  & (\all_features[1276]  | \all_features[1277]  | new_n24049_ | ~new_n24050_);
  assign new_n24049_ = \all_features[1272]  & \all_features[1273] ;
  assign new_n24050_ = ~\all_features[1274]  & ~\all_features[1275] ;
  assign new_n24051_ = ~\all_features[1275]  & ~\all_features[1276]  & (~\all_features[1274]  | new_n24052_);
  assign new_n24052_ = ~\all_features[1272]  & ~\all_features[1273] ;
  assign new_n24053_ = ~new_n24054_ & ~\all_features[1279] ;
  assign new_n24054_ = \all_features[1277]  & \all_features[1278]  & (\all_features[1276]  | (\all_features[1274]  & \all_features[1275]  & \all_features[1273] ));
  assign new_n24055_ = ~\all_features[1279]  & (~\all_features[1278]  | ~new_n24056_ | ~new_n24049_ | ~new_n24047_);
  assign new_n24056_ = \all_features[1274]  & \all_features[1275] ;
  assign new_n24057_ = \all_features[1279]  & (\all_features[1278]  | (\all_features[1277]  & (\all_features[1276]  | ~new_n24050_ | ~new_n24052_)));
  assign new_n24058_ = \all_features[1279]  & (\all_features[1277]  | \all_features[1278]  | \all_features[1276] );
  assign new_n24059_ = ~new_n24060_ & (\all_features[1275]  | \all_features[1276]  | \all_features[1277]  | \all_features[1278]  | \all_features[1279] );
  assign new_n24060_ = ~\all_features[1277]  & new_n24061_ & ((~\all_features[1274]  & new_n24052_) | ~\all_features[1276]  | ~\all_features[1275] );
  assign new_n24061_ = ~\all_features[1278]  & ~\all_features[1279] ;
  assign new_n24062_ = ~new_n24063_ & ~new_n24064_;
  assign new_n24063_ = new_n24061_ & (~\all_features[1277]  | (~\all_features[1276]  & (~\all_features[1275]  | (~\all_features[1274]  & ~\all_features[1273] ))));
  assign new_n24064_ = new_n24061_ & (~\all_features[1275]  | ~new_n24047_ | (~\all_features[1274]  & ~new_n24049_));
  assign new_n24065_ = ~\all_features[1279]  & (~\all_features[1278]  | (~\all_features[1277]  & (new_n24052_ | ~new_n24056_ | ~\all_features[1276] )));
  assign new_n24066_ = ~\all_features[1279]  & (~\all_features[1278]  | (~\all_features[1276]  & ~\all_features[1277]  & ~new_n24056_));
  assign new_n24067_ = ~new_n24068_ & ~new_n24070_;
  assign new_n24068_ = new_n24069_ & new_n24059_ & ~new_n24064_ & ~new_n24065_ & ~new_n24053_ & ~new_n24063_;
  assign new_n24069_ = ~new_n24055_ & ~new_n24066_;
  assign new_n24070_ = new_n24059_ & new_n24062_ & (new_n24071_ | new_n24053_ | new_n24065_ | ~new_n24069_);
  assign new_n24071_ = new_n24058_ & new_n24048_ & new_n24057_ & new_n24046_;
  assign new_n24072_ = ~new_n24073_ & (\all_features[1275]  | \all_features[1276]  | \all_features[1277]  | \all_features[1278]  | \all_features[1279] );
  assign new_n24073_ = ~new_n24060_ & (new_n24063_ | (~new_n24064_ & (new_n24066_ | (~new_n24065_ & ~new_n24074_))));
  assign new_n24074_ = ~new_n24053_ & (new_n24055_ | (new_n24058_ & (~new_n24057_ | (~new_n24075_ & new_n24046_))));
  assign new_n24075_ = ~\all_features[1277]  & \all_features[1278]  & \all_features[1279]  & (\all_features[1276]  ? new_n24050_ : (new_n24049_ | ~new_n24050_));
  assign new_n24076_ = ~new_n9606_ & (~new_n9584_ | ~new_n10526_);
  assign new_n24077_ = ~new_n24110_ & ~new_n24099_ & ~new_n24107_ & (new_n24105_ | (~new_n24104_ & ~new_n24078_));
  assign new_n24078_ = ~new_n24092_ & (new_n24094_ | (~new_n24095_ & (new_n24096_ | (~new_n24079_ & ~new_n24097_))));
  assign new_n24079_ = ~new_n24086_ & (~new_n24090_ | (new_n24080_ & (~new_n24089_ | (~new_n24091_ & new_n24083_))));
  assign new_n24080_ = \all_features[2663]  & (\all_features[2662]  | new_n24081_);
  assign new_n24081_ = \all_features[2661]  & (\all_features[2658]  | \all_features[2659]  | \all_features[2660]  | ~new_n24082_);
  assign new_n24082_ = ~\all_features[2656]  & ~\all_features[2657] ;
  assign new_n24083_ = \all_features[2663]  & ~new_n24084_ & \all_features[2662] ;
  assign new_n24084_ = ~\all_features[2661]  & ~\all_features[2660]  & ~\all_features[2659]  & ~new_n24085_ & ~\all_features[2658] ;
  assign new_n24085_ = \all_features[2656]  & \all_features[2657] ;
  assign new_n24086_ = ~\all_features[2663]  & (~\all_features[2662]  | ~new_n24085_ | ~new_n24087_ | ~new_n24088_);
  assign new_n24087_ = \all_features[2660]  & \all_features[2661] ;
  assign new_n24088_ = \all_features[2658]  & \all_features[2659] ;
  assign new_n24089_ = \all_features[2663]  & (\all_features[2662]  | (new_n24087_ & (\all_features[2658]  | \all_features[2659]  | \all_features[2657] )));
  assign new_n24090_ = \all_features[2663]  & (\all_features[2661]  | \all_features[2662]  | \all_features[2660] );
  assign new_n24091_ = \all_features[2662]  & \all_features[2663]  & (\all_features[2661]  | (\all_features[2660]  & (\all_features[2659]  | \all_features[2658] )));
  assign new_n24092_ = new_n24093_ & (~\all_features[2661]  | (~\all_features[2660]  & (~\all_features[2659]  | (~\all_features[2658]  & ~\all_features[2657] ))));
  assign new_n24093_ = ~\all_features[2662]  & ~\all_features[2663] ;
  assign new_n24094_ = new_n24093_ & (~\all_features[2659]  | ~new_n24087_ | (~\all_features[2658]  & ~new_n24085_));
  assign new_n24095_ = ~\all_features[2663]  & (~\all_features[2662]  | (~\all_features[2660]  & ~\all_features[2661]  & ~new_n24088_));
  assign new_n24096_ = ~\all_features[2663]  & (~\all_features[2662]  | (~\all_features[2661]  & (new_n24082_ | ~new_n24088_ | ~\all_features[2660] )));
  assign new_n24097_ = ~new_n24098_ & ~\all_features[2663] ;
  assign new_n24098_ = \all_features[2661]  & \all_features[2662]  & (\all_features[2660]  | (\all_features[2658]  & \all_features[2659]  & \all_features[2657] ));
  assign new_n24099_ = new_n24103_ & (~new_n24106_ | (~new_n24100_ & ~new_n24095_ & ~new_n24096_));
  assign new_n24100_ = ~new_n24086_ & ~new_n24097_ & (~new_n24090_ | new_n24101_ | ~new_n24080_);
  assign new_n24101_ = ~new_n24084_ & new_n24089_ & \all_features[2662]  & \all_features[2663]  & (~\all_features[2661]  | new_n24102_);
  assign new_n24102_ = ~\all_features[2659]  & ~\all_features[2660]  & (~\all_features[2658]  | new_n24082_);
  assign new_n24103_ = ~new_n24104_ & ~new_n24105_;
  assign new_n24104_ = ~\all_features[2661]  & new_n24093_ & ((~\all_features[2658]  & new_n24082_) | ~\all_features[2660]  | ~\all_features[2659] );
  assign new_n24105_ = ~\all_features[2663]  & ~\all_features[2662]  & ~\all_features[2661]  & ~\all_features[2659]  & ~\all_features[2660] ;
  assign new_n24106_ = ~new_n24092_ & ~new_n24094_;
  assign new_n24107_ = new_n24106_ & ~new_n24108_ & new_n24103_;
  assign new_n24108_ = new_n24109_ & (~new_n24089_ | ~new_n24090_ | ~new_n24083_ | ~new_n24080_);
  assign new_n24109_ = ~new_n24086_ & ~new_n24097_ & ~new_n24095_ & ~new_n24096_;
  assign new_n24110_ = new_n24111_ & new_n24103_ & ~new_n24092_ & ~new_n24097_;
  assign new_n24111_ = ~new_n24086_ & ~new_n24096_ & ~new_n24094_ & ~new_n24095_;
  assign new_n24112_ = new_n11820_ & new_n11823_;
  assign new_n24113_ = ~new_n21615_ & new_n24076_ & new_n16567_ & (new_n23476_ | (new_n23451_ & new_n23478_));
  assign new_n24114_ = (new_n24120_ & new_n24076_ & (new_n21615_ | ~new_n24122_)) | (new_n24115_ & ~new_n24123_ & ~new_n24076_);
  assign new_n24115_ = (new_n24116_ | new_n24117_ | ~new_n12117_) & (new_n12117_ | (new_n7443_ ? new_n23557_ : new_n24119_));
  assign new_n24116_ = ~new_n10761_ & (~new_n10739_ | new_n10762_);
  assign new_n24117_ = new_n17589_ & new_n24118_;
  assign new_n24118_ = ~new_n17619_ & ~new_n17621_;
  assign new_n24119_ = new_n21108_ & new_n21106_ & new_n21078_ & new_n21102_;
  assign new_n24120_ = (~new_n24121_ | new_n21615_ | (~new_n15409_ & new_n16103_)) & (~new_n23139_ | new_n19089_ | ~new_n21615_);
  assign new_n24121_ = new_n9726_ & (~new_n9755_ | ~new_n9751_);
  assign new_n24122_ = ~new_n24121_ & ~new_n19238_;
  assign new_n24123_ = new_n20436_ & new_n20408_ & new_n12117_ & new_n24117_;
  assign new_n24124_ = new_n24125_ ? (~new_n24328_ ^ new_n24349_) : (new_n24328_ ^ new_n24349_);
  assign new_n24125_ = new_n24126_ ? (new_n24195_ ^ new_n24253_) : (~new_n24195_ ^ new_n24253_);
  assign new_n24126_ = new_n24127_ ? (new_n24149_ ^ new_n24175_) : (~new_n24149_ ^ new_n24175_);
  assign new_n24127_ = ~new_n24128_ & new_n24146_;
  assign new_n24128_ = new_n24129_ & new_n24140_ & (~new_n24142_ | (~new_n24143_ & new_n24077_) | (~new_n24145_ & ~new_n24077_));
  assign new_n24129_ = (~new_n24135_ | ~new_n24133_) & (~new_n24130_ | (new_n24132_ ? ~new_n24134_ : new_n16658_));
  assign new_n24130_ = ~new_n24005_ & new_n24131_;
  assign new_n24131_ = ~new_n13805_ & new_n6885_;
  assign new_n24132_ = new_n22898_ & new_n24026_;
  assign new_n24133_ = new_n14336_ & ~new_n21692_ & ~new_n24131_;
  assign new_n24134_ = ~new_n15032_ & new_n10702_;
  assign new_n24135_ = new_n9544_ & (~new_n9518_ | (~new_n9543_ & (new_n9542_ | new_n24136_)));
  assign new_n24136_ = ~new_n9540_ & (new_n9538_ | (~new_n9521_ & (new_n9523_ | (~new_n24137_ & ~new_n9533_))));
  assign new_n24137_ = ~new_n9535_ & (~\all_features[3999]  | new_n24138_ | (~\all_features[3996]  & ~\all_features[3997]  & ~\all_features[3998] ));
  assign new_n24138_ = \all_features[3999]  & ((~new_n24139_ & ~\all_features[3997]  & \all_features[3998] ) | (~new_n9530_ & (\all_features[3998]  | (~new_n9526_ & \all_features[3997] ))));
  assign new_n24139_ = (~\all_features[3994]  & ~\all_features[3995]  & ~\all_features[3996]  & (~\all_features[3993]  | ~\all_features[3992] )) | (\all_features[3996]  & (\all_features[3994]  | \all_features[3995] ));
  assign new_n24140_ = (~new_n24141_ | new_n24131_) & (~new_n24005_ | ~new_n24131_ | (new_n9313_ ? new_n24119_ : ~new_n19125_));
  assign new_n24141_ = new_n14336_ & new_n21692_;
  assign new_n24142_ = ~new_n14336_ & ~new_n24131_;
  assign new_n24143_ = ~new_n20924_ & new_n24144_;
  assign new_n24144_ = ~new_n20954_ & ~new_n20956_;
  assign new_n24145_ = new_n15143_ & (~new_n15139_ | ~new_n15115_);
  assign new_n24146_ = ~new_n24148_ & new_n24147_ & (~new_n24142_ | (new_n24143_ & new_n24077_) | (new_n24145_ & ~new_n24077_));
  assign new_n24147_ = (~new_n24133_ | new_n24135_) & (~new_n24130_ | (new_n24132_ ? new_n24134_ : ~new_n16658_));
  assign new_n24148_ = new_n24131_ & new_n24005_ & ~new_n9313_ & ~new_n19125_;
  assign new_n24149_ = ~new_n24150_ & new_n24172_;
  assign new_n24150_ = new_n24151_ & (~new_n24171_ | (new_n19548_ & new_n24170_) | (~new_n22998_ & ~new_n24170_));
  assign new_n24151_ = new_n24152_ & (~new_n24162_ | (~new_n24163_ & new_n21605_) | (~new_n24164_ & ~new_n21605_));
  assign new_n24152_ = ~new_n24155_ & ~new_n24159_ & (~new_n24160_ | (~new_n24153_ & ~new_n20158_) | (~new_n21571_ & new_n20158_));
  assign new_n24153_ = ~new_n24154_ & ~new_n12791_;
  assign new_n24154_ = ~new_n18894_ & new_n12762_;
  assign new_n24155_ = ~new_n8985_ & new_n17937_ & new_n24156_ & new_n24157_ & (~new_n8963_ | new_n24158_);
  assign new_n24156_ = ~new_n8232_ & ~new_n8264_;
  assign new_n24157_ = new_n16446_ & (new_n16448_ | (new_n16442_ & new_n16418_));
  assign new_n24158_ = ~new_n8987_ & ~new_n11624_;
  assign new_n24159_ = new_n17937_ & ~new_n24157_ & new_n24156_;
  assign new_n24160_ = ~new_n24156_ & ~new_n24161_;
  assign new_n24161_ = new_n12376_ & new_n12398_;
  assign new_n24162_ = ~new_n17937_ & new_n24156_;
  assign new_n24163_ = new_n19677_ & (new_n19651_ | new_n21401_);
  assign new_n24164_ = ~new_n18288_ & (~new_n24165_ | ~new_n18259_);
  assign new_n24165_ = (new_n24166_ | (new_n18284_ & (~\all_features[4819]  | ~\all_features[4820]  | (~\all_features[4818]  & new_n18264_)))) & (~new_n18284_ | \all_features[4819]  | \all_features[4820] );
  assign new_n24166_ = ~new_n18273_ & (new_n18272_ | (~new_n18276_ & (new_n18278_ | (~new_n24167_ & ~new_n18281_))));
  assign new_n24167_ = ~new_n18280_ & (~\all_features[4823]  | new_n24168_ | (~\all_features[4820]  & ~\all_features[4821]  & ~\all_features[4822] ));
  assign new_n24168_ = \all_features[4823]  & ((~new_n24169_ & ~\all_features[4821]  & \all_features[4822] ) | (~new_n18266_ & (\all_features[4822]  | (~new_n18263_ & \all_features[4821] ))));
  assign new_n24169_ = (\all_features[4820]  & (\all_features[4818]  | \all_features[4819] )) | (~new_n18269_ & ~\all_features[4818]  & ~\all_features[4819]  & ~\all_features[4820] );
  assign new_n24170_ = new_n21703_ & new_n11201_;
  assign new_n24171_ = ~new_n24156_ & new_n24161_;
  assign new_n24172_ = new_n24173_ & (~new_n24171_ | (~new_n19548_ & new_n24170_) | (new_n22998_ & ~new_n24170_));
  assign new_n24173_ = ~new_n24174_ & (~new_n24160_ | (new_n24153_ & ~new_n20158_) | (new_n21571_ & new_n20158_));
  assign new_n24174_ = new_n24162_ & (new_n21605_ ? ~new_n24163_ : ~new_n24164_);
  assign new_n24175_ = new_n24183_ & ~new_n24176_ & ~new_n24194_;
  assign new_n24176_ = new_n24181_ & ((~new_n24177_ & ~new_n14469_) | (~new_n19500_ & new_n24182_ & new_n14469_));
  assign new_n24177_ = (new_n24180_ & new_n10682_) ? new_n24178_ : ~new_n8697_;
  assign new_n24178_ = new_n16105_ & new_n24179_;
  assign new_n24179_ = new_n15860_ & new_n15862_;
  assign new_n24180_ = new_n13924_ & new_n13933_;
  assign new_n24181_ = new_n21570_ & new_n22929_;
  assign new_n24182_ = ~new_n6495_ & (~new_n6491_ | ~new_n6461_);
  assign new_n24183_ = (new_n24184_ | new_n24185_ | new_n24181_) & (new_n24182_ | ~new_n14469_ | ~new_n24181_);
  assign new_n24184_ = (~new_n7443_ & ~new_n18045_) | (new_n16101_ & new_n18045_ & (new_n16098_ | new_n16065_));
  assign new_n24185_ = new_n12537_ & (~new_n24190_ | ~new_n24186_);
  assign new_n24186_ = new_n12540_ & (new_n12545_ | new_n12544_ | (~new_n12549_ & ~new_n12554_ & ~new_n24187_));
  assign new_n24187_ = ~new_n12553_ & ~new_n12551_ & (~new_n12559_ | ~new_n12555_ | new_n24188_);
  assign new_n24188_ = new_n12557_ & new_n12558_ & (new_n24189_ | ~\all_features[3533]  | ~\all_features[3534]  | ~\all_features[3535] );
  assign new_n24189_ = ~\all_features[3531]  & ~\all_features[3532]  & (~\all_features[3530]  | new_n12542_);
  assign new_n24190_ = ~new_n24191_ & (\all_features[3531]  | \all_features[3532]  | \all_features[3533]  | \all_features[3534]  | \all_features[3535] );
  assign new_n24191_ = ~new_n12541_ & (new_n12544_ | (~new_n12545_ & (new_n12554_ | (~new_n12549_ & ~new_n24192_))));
  assign new_n24192_ = ~new_n12551_ & (new_n12553_ | (new_n12559_ & (~new_n12555_ | (~new_n24193_ & new_n12557_))));
  assign new_n24193_ = ~\all_features[3533]  & \all_features[3534]  & \all_features[3535]  & (\all_features[3532]  ? new_n12556_ : (new_n12547_ | ~new_n12556_));
  assign new_n24194_ = ~new_n24181_ & new_n24185_ & ((~new_n22997_ & ~new_n23971_) | (new_n23551_ & new_n15518_ & new_n23971_));
  assign new_n24195_ = new_n24196_ ? (new_n24211_ ^ new_n24212_) : (~new_n24211_ ^ new_n24212_);
  assign new_n24196_ = new_n24205_ ? ((new_n24202_ | ~new_n24204_) & (new_n14336_ | new_n10681_ | new_n24204_)) : ~new_n24197_;
  assign new_n24197_ = new_n24200_ ? new_n24198_ : (new_n7803_ ? ~new_n24199_ : ~new_n24201_);
  assign new_n24198_ = ~new_n13405_ & (new_n15745_ | ~new_n22790_);
  assign new_n24199_ = ~new_n6627_ & (~new_n6605_ | new_n6629_);
  assign new_n24200_ = new_n14154_ & (new_n14156_ | ~new_n14784_);
  assign new_n24201_ = new_n9482_ & new_n9460_ & new_n12842_;
  assign new_n24202_ = new_n24203_ ? ~new_n23605_ : ~new_n15713_;
  assign new_n24203_ = ~new_n21352_ & new_n11160_;
  assign new_n24204_ = ~new_n7736_ & (~new_n7733_ | ~new_n7722_);
  assign new_n24205_ = ~new_n15265_ & ~new_n24206_ & ~new_n21626_ & ~new_n21636_;
  assign new_n24206_ = ~new_n15267_ & (new_n15277_ | (~new_n15274_ & (new_n15272_ | (~new_n15269_ & ~new_n24207_))));
  assign new_n24207_ = ~new_n15280_ & (new_n15275_ | (~new_n15279_ & (~new_n24210_ | new_n24208_)));
  assign new_n24208_ = \all_features[1047]  & ((~new_n24209_ & ~\all_features[1045]  & \all_features[1046] ) | (~new_n21633_ & (\all_features[1046]  | (~new_n21629_ & \all_features[1045] ))));
  assign new_n24209_ = (~\all_features[1042]  & ~\all_features[1043]  & ~\all_features[1044]  & (~\all_features[1041]  | ~\all_features[1040] )) | (\all_features[1044]  & (\all_features[1042]  | \all_features[1043] ));
  assign new_n24210_ = \all_features[1047]  & (\all_features[1045]  | \all_features[1046]  | \all_features[1044] );
  assign new_n24211_ = ~new_n23938_ & new_n23932_;
  assign new_n24212_ = ~new_n24213_ & new_n24251_;
  assign new_n24213_ = ~new_n24214_ & (new_n20870_ | new_n12791_ | ~new_n24250_);
  assign new_n24214_ = new_n24216_ & (new_n24249_ ? new_n24248_ : new_n24215_);
  assign new_n24215_ = new_n24154_ & new_n12791_;
  assign new_n24216_ = ~new_n20048_ & ~new_n24217_;
  assign new_n24217_ = ~new_n24218_ & new_n24240_ & (new_n24247_ | new_n24223_ | new_n24225_ | ~new_n24245_);
  assign new_n24218_ = ~new_n24233_ & (new_n24235_ | (~new_n24237_ & (new_n24238_ | (~new_n24219_ & ~new_n24239_))));
  assign new_n24219_ = ~new_n24223_ & (new_n24225_ | (new_n24232_ & (~new_n24220_ | (~new_n24229_ & new_n24231_))));
  assign new_n24220_ = \all_features[4903]  & (\all_features[4902]  | new_n24221_);
  assign new_n24221_ = \all_features[4901]  & (\all_features[4898]  | \all_features[4899]  | \all_features[4900]  | ~new_n24222_);
  assign new_n24222_ = ~\all_features[4896]  & ~\all_features[4897] ;
  assign new_n24223_ = ~new_n24224_ & ~\all_features[4903] ;
  assign new_n24224_ = \all_features[4901]  & \all_features[4902]  & (\all_features[4900]  | (\all_features[4898]  & \all_features[4899]  & \all_features[4897] ));
  assign new_n24225_ = ~\all_features[4903]  & (~\all_features[4902]  | ~new_n24226_ | ~new_n24227_ | ~new_n24228_);
  assign new_n24226_ = \all_features[4896]  & \all_features[4897] ;
  assign new_n24227_ = \all_features[4900]  & \all_features[4901] ;
  assign new_n24228_ = \all_features[4898]  & \all_features[4899] ;
  assign new_n24229_ = ~\all_features[4901]  & new_n24230_ & ((~\all_features[4900]  & (new_n24226_ | \all_features[4898]  | \all_features[4899] )) | (~\all_features[4898]  & ~\all_features[4899]  & \all_features[4900] ));
  assign new_n24230_ = \all_features[4902]  & \all_features[4903] ;
  assign new_n24231_ = \all_features[4903]  & (\all_features[4902]  | (new_n24227_ & (\all_features[4898]  | \all_features[4899]  | \all_features[4897] )));
  assign new_n24232_ = \all_features[4903]  & (\all_features[4901]  | \all_features[4902]  | \all_features[4900] );
  assign new_n24233_ = new_n24234_ & ((~\all_features[4898]  & new_n24222_) | ~\all_features[4900]  | ~\all_features[4899] );
  assign new_n24234_ = ~\all_features[4903]  & ~\all_features[4901]  & ~\all_features[4902] ;
  assign new_n24235_ = ~\all_features[4903]  & ~new_n24236_ & ~\all_features[4902] ;
  assign new_n24236_ = \all_features[4901]  & (\all_features[4900]  | (\all_features[4899]  & (\all_features[4898]  | \all_features[4897] )));
  assign new_n24237_ = ~\all_features[4902]  & ~\all_features[4903]  & (~\all_features[4899]  | ~new_n24227_ | (~\all_features[4898]  & ~new_n24226_));
  assign new_n24238_ = ~\all_features[4903]  & (~\all_features[4902]  | (~\all_features[4900]  & ~\all_features[4901]  & ~new_n24228_));
  assign new_n24239_ = ~\all_features[4903]  & (~\all_features[4902]  | (~\all_features[4901]  & (new_n24222_ | ~new_n24228_ | ~\all_features[4900] )));
  assign new_n24240_ = ~new_n24235_ & ~new_n24223_ & new_n24246_ & new_n24245_ & (new_n24225_ | new_n24241_);
  assign new_n24241_ = new_n24232_ & ~new_n24242_ & new_n24220_;
  assign new_n24242_ = new_n24231_ & new_n24243_ & (~\all_features[4901]  | ~new_n24230_ | new_n24244_);
  assign new_n24243_ = new_n24230_ & (new_n24226_ | \all_features[4898]  | \all_features[4899]  | \all_features[4900]  | \all_features[4901] );
  assign new_n24244_ = ~\all_features[4899]  & ~\all_features[4900]  & (~\all_features[4898]  | new_n24222_);
  assign new_n24245_ = ~new_n24238_ & ~new_n24239_;
  assign new_n24246_ = ~new_n24233_ & ~new_n24237_ & ~new_n24225_ & (\all_features[4900]  | \all_features[4899]  | ~new_n24234_);
  assign new_n24247_ = new_n24232_ & new_n24231_ & new_n24220_ & new_n24243_;
  assign new_n24248_ = new_n7550_ & (new_n7547_ | ~new_n7517_);
  assign new_n24249_ = new_n8031_ & new_n9649_;
  assign new_n24250_ = ~new_n24217_ & new_n20048_;
  assign new_n24251_ = ~new_n24252_ & (~new_n24216_ | (new_n24215_ & ~new_n24249_) | (new_n24248_ & new_n24249_));
  assign new_n24252_ = new_n24250_ & (new_n12791_ | new_n20870_);
  assign new_n24253_ = new_n24254_ & new_n24326_;
  assign new_n24254_ = new_n24255_ & (~new_n24258_ | new_n24257_) & (new_n16410_ | new_n24292_ | ~new_n24008_ | ~new_n24257_);
  assign new_n24255_ = ~new_n24257_ | ((~new_n16410_ | ~new_n24256_ | ~new_n24008_) & (new_n19197_ | ~new_n23065_ | new_n24008_));
  assign new_n24256_ = ~new_n8666_ & new_n11167_;
  assign new_n24257_ = ~new_n20533_ & ~new_n20531_ & ~new_n20519_;
  assign new_n24258_ = new_n24259_ ? (~new_n24288_ & (~new_n24260_ | ~new_n24281_ | ~new_n24290_)) : ~new_n13391_;
  assign new_n24259_ = new_n10271_ & ~new_n10272_ & new_n10249_;
  assign new_n24260_ = ~new_n24261_ & (\all_features[1403]  | \all_features[1404]  | \all_features[1405]  | \all_features[1406]  | \all_features[1407] );
  assign new_n24261_ = ~new_n24277_ & (new_n24275_ | (~new_n24279_ & (new_n24280_ | (~new_n24278_ & ~new_n24262_))));
  assign new_n24262_ = ~new_n24263_ & (new_n24265_ | (new_n24274_ & (~new_n24269_ | (~new_n24273_ & new_n24272_))));
  assign new_n24263_ = ~new_n24264_ & ~\all_features[1407] ;
  assign new_n24264_ = \all_features[1405]  & \all_features[1406]  & (\all_features[1404]  | (\all_features[1402]  & \all_features[1403]  & \all_features[1401] ));
  assign new_n24265_ = ~\all_features[1407]  & (~\all_features[1406]  | ~new_n24266_ | ~new_n24267_ | ~new_n24268_);
  assign new_n24266_ = \all_features[1402]  & \all_features[1403] ;
  assign new_n24267_ = \all_features[1400]  & \all_features[1401] ;
  assign new_n24268_ = \all_features[1404]  & \all_features[1405] ;
  assign new_n24269_ = \all_features[1407]  & (\all_features[1406]  | (\all_features[1405]  & (\all_features[1404]  | ~new_n24271_ | ~new_n24270_)));
  assign new_n24270_ = ~\all_features[1400]  & ~\all_features[1401] ;
  assign new_n24271_ = ~\all_features[1402]  & ~\all_features[1403] ;
  assign new_n24272_ = \all_features[1407]  & (\all_features[1406]  | (new_n24268_ & (\all_features[1402]  | \all_features[1403]  | \all_features[1401] )));
  assign new_n24273_ = ~\all_features[1405]  & \all_features[1406]  & \all_features[1407]  & (\all_features[1404]  ? new_n24271_ : (new_n24267_ | ~new_n24271_));
  assign new_n24274_ = \all_features[1407]  & (\all_features[1405]  | \all_features[1406]  | \all_features[1404] );
  assign new_n24275_ = new_n24276_ & (~\all_features[1405]  | (~\all_features[1404]  & (~\all_features[1403]  | (~\all_features[1402]  & ~\all_features[1401] ))));
  assign new_n24276_ = ~\all_features[1406]  & ~\all_features[1407] ;
  assign new_n24277_ = ~\all_features[1405]  & new_n24276_ & ((~\all_features[1402]  & new_n24270_) | ~\all_features[1404]  | ~\all_features[1403] );
  assign new_n24278_ = ~\all_features[1407]  & (~\all_features[1406]  | (~\all_features[1405]  & (new_n24270_ | ~new_n24266_ | ~\all_features[1404] )));
  assign new_n24279_ = new_n24276_ & (~\all_features[1403]  | ~new_n24268_ | (~\all_features[1402]  & ~new_n24267_));
  assign new_n24280_ = ~\all_features[1407]  & (~\all_features[1406]  | (~\all_features[1404]  & ~\all_features[1405]  & ~new_n24266_));
  assign new_n24281_ = new_n24286_ & (~new_n24287_ | (~new_n24282_ & ~new_n24278_ & ~new_n24280_));
  assign new_n24282_ = ~new_n24263_ & ~new_n24265_ & (~new_n24274_ | ~new_n24269_ | new_n24283_);
  assign new_n24283_ = new_n24272_ & new_n24284_ & (new_n24285_ | ~\all_features[1405]  | ~\all_features[1406]  | ~\all_features[1407] );
  assign new_n24284_ = \all_features[1406]  & \all_features[1407]  & (\all_features[1404]  | \all_features[1405]  | new_n24267_ | ~new_n24271_);
  assign new_n24285_ = ~\all_features[1403]  & ~\all_features[1404]  & (~\all_features[1402]  | new_n24270_);
  assign new_n24286_ = ~new_n24277_ & (\all_features[1403]  | \all_features[1404]  | \all_features[1405]  | \all_features[1406]  | \all_features[1407] );
  assign new_n24287_ = ~new_n24275_ & ~new_n24279_;
  assign new_n24288_ = new_n24289_ & new_n24286_ & ~new_n24279_ & ~new_n24278_ & ~new_n24263_ & ~new_n24275_;
  assign new_n24289_ = ~new_n24265_ & ~new_n24280_;
  assign new_n24290_ = new_n24286_ & new_n24287_ & (new_n24291_ | new_n24263_ | new_n24278_ | ~new_n24289_);
  assign new_n24291_ = new_n24274_ & new_n24284_ & new_n24269_ & new_n24272_;
  assign new_n24292_ = new_n24324_ & new_n24322_ & new_n24293_ & new_n24315_;
  assign new_n24293_ = ~new_n24314_ & (new_n24309_ | (~new_n24311_ & (new_n24312_ | (~new_n24294_ & ~new_n24313_))));
  assign new_n24294_ = ~new_n24301_ & (new_n24304_ | (~new_n24306_ & (~new_n24308_ | (~new_n24295_ & new_n24307_))));
  assign new_n24295_ = new_n24296_ & (\all_features[2517]  | ~new_n24300_ | (~new_n24298_ & ~\all_features[2516]  & new_n24299_) | (\all_features[2516]  & ~new_n24299_));
  assign new_n24296_ = \all_features[2519]  & (\all_features[2518]  | (new_n24297_ & (\all_features[2514]  | \all_features[2515]  | \all_features[2513] )));
  assign new_n24297_ = \all_features[2516]  & \all_features[2517] ;
  assign new_n24298_ = \all_features[2512]  & \all_features[2513] ;
  assign new_n24299_ = ~\all_features[2514]  & ~\all_features[2515] ;
  assign new_n24300_ = \all_features[2518]  & \all_features[2519] ;
  assign new_n24301_ = ~\all_features[2519]  & (~\all_features[2518]  | (~\all_features[2517]  & (new_n24302_ | ~new_n24303_ | ~\all_features[2516] )));
  assign new_n24302_ = ~\all_features[2512]  & ~\all_features[2513] ;
  assign new_n24303_ = \all_features[2514]  & \all_features[2515] ;
  assign new_n24304_ = ~new_n24305_ & ~\all_features[2519] ;
  assign new_n24305_ = \all_features[2517]  & \all_features[2518]  & (\all_features[2516]  | (\all_features[2514]  & \all_features[2515]  & \all_features[2513] ));
  assign new_n24306_ = ~\all_features[2519]  & (~\all_features[2518]  | ~new_n24298_ | ~new_n24297_ | ~new_n24303_);
  assign new_n24307_ = \all_features[2519]  & (\all_features[2518]  | (\all_features[2517]  & (\all_features[2516]  | ~new_n24299_ | ~new_n24302_)));
  assign new_n24308_ = \all_features[2519]  & (\all_features[2517]  | \all_features[2518]  | \all_features[2516] );
  assign new_n24309_ = ~\all_features[2517]  & new_n24310_ & ((~\all_features[2514]  & new_n24302_) | ~\all_features[2516]  | ~\all_features[2515] );
  assign new_n24310_ = ~\all_features[2518]  & ~\all_features[2519] ;
  assign new_n24311_ = new_n24310_ & (~\all_features[2517]  | (~\all_features[2516]  & (~\all_features[2515]  | (~\all_features[2514]  & ~\all_features[2513] ))));
  assign new_n24312_ = new_n24310_ & (~\all_features[2515]  | ~new_n24297_ | (~\all_features[2514]  & ~new_n24298_));
  assign new_n24313_ = ~\all_features[2519]  & (~\all_features[2518]  | (~\all_features[2516]  & ~\all_features[2517]  & ~new_n24303_));
  assign new_n24314_ = ~\all_features[2519]  & ~\all_features[2518]  & ~\all_features[2517]  & ~\all_features[2515]  & ~\all_features[2516] ;
  assign new_n24315_ = ~new_n24309_ & ~new_n24314_ & (~new_n24320_ | (~new_n24316_ & new_n24321_));
  assign new_n24316_ = new_n24317_ & ((~new_n24319_ & new_n24318_ & new_n24296_) | ~new_n24308_ | ~new_n24307_);
  assign new_n24317_ = ~new_n24304_ & ~new_n24306_;
  assign new_n24318_ = new_n24300_ & (new_n24298_ | \all_features[2516]  | \all_features[2517]  | ~new_n24299_);
  assign new_n24319_ = new_n24300_ & \all_features[2517]  & ((~new_n24302_ & \all_features[2514] ) | \all_features[2516]  | \all_features[2515] );
  assign new_n24320_ = ~new_n24311_ & ~new_n24312_;
  assign new_n24321_ = ~new_n24313_ & ~new_n24301_;
  assign new_n24322_ = ~new_n24314_ & ~new_n24312_ & ~new_n24311_ & ~new_n24323_ & ~new_n24309_;
  assign new_n24323_ = new_n24321_ & new_n24317_ & (~new_n24318_ | ~new_n24308_ | ~new_n24307_ | ~new_n24296_);
  assign new_n24324_ = new_n24325_ & new_n24320_ & ~new_n24304_ & ~new_n24301_ & ~new_n24309_ & ~new_n24313_;
  assign new_n24325_ = ~new_n24306_ & ~new_n24314_;
  assign new_n24326_ = new_n24257_ ? ((new_n16410_ | ~new_n24292_ | ~new_n24008_) & (new_n24327_ | new_n24008_)) : new_n24258_;
  assign new_n24327_ = ~new_n19197_ & new_n23065_;
  assign new_n24328_ = new_n24329_ & (~new_n24343_ | ~new_n24340_ | ~new_n19238_);
  assign new_n24329_ = new_n24330_ & (new_n24342_ | ~new_n24331_ | ~new_n13523_) & (new_n19238_ | ~new_n24340_);
  assign new_n24330_ = (~new_n24337_ | ~new_n24333_) & (new_n24339_ | new_n13523_ | ~new_n24331_);
  assign new_n24331_ = ~new_n11130_ & new_n24332_;
  assign new_n24332_ = new_n18340_ & ~new_n18364_ & ~new_n18368_;
  assign new_n24333_ = new_n23765_ & ~new_n24334_ & ~new_n24336_;
  assign new_n24334_ = new_n18798_ & new_n24335_;
  assign new_n24335_ = ~new_n11274_ & ~new_n11301_;
  assign new_n24336_ = new_n23737_ & new_n23761_;
  assign new_n24337_ = ~new_n24332_ & ~new_n24338_;
  assign new_n24338_ = ~new_n24068_ & (~new_n24043_ | ~new_n24072_ | ~new_n24070_);
  assign new_n24339_ = new_n15745_ & (new_n15743_ | ~new_n16027_);
  assign new_n24340_ = ~new_n24077_ & new_n24341_;
  assign new_n24341_ = new_n11130_ & new_n24332_;
  assign new_n24342_ = ~new_n9163_ & ~new_n9165_;
  assign new_n24343_ = new_n24344_ & new_n24347_ & (~new_n24337_ | new_n24333_);
  assign new_n24344_ = (new_n24346_ | ~new_n21484_ | ~new_n24345_ | ~new_n12141_) & (~new_n24341_ | ~new_n24077_);
  assign new_n24345_ = ~new_n24332_ & new_n24338_;
  assign new_n24346_ = ~new_n12119_ & ~new_n12147_;
  assign new_n24347_ = ~new_n24348_ & (~new_n24331_ | (~new_n24339_ & ~new_n13523_) | (~new_n24342_ & new_n13523_));
  assign new_n24348_ = ~new_n21484_ & new_n24345_;
  assign new_n24349_ = ~new_n24350_ & ~new_n24351_ & (~new_n19717_ | ~new_n17214_ | new_n14162_ | new_n22423_);
  assign new_n24350_ = ~new_n17214_ & ~new_n8164_ & ~new_n14329_ & (~new_n11164_ | (~new_n11161_ & new_n11131_));
  assign new_n24351_ = new_n17214_ & new_n14162_ & (new_n22693_ ? (~new_n13360_ | ~new_n14724_) : ~new_n24352_);
  assign new_n24352_ = ~new_n6953_ & (~new_n6950_ | ~new_n18795_);
  assign new_n24353_ = ~new_n24354_ & new_n24364_;
  assign new_n24354_ = new_n24355_ & (~new_n24363_ | ~new_n24362_);
  assign new_n24355_ = new_n24356_ & (new_n24361_ | ~new_n24359_ | new_n24357_) & (new_n18189_ | new_n24360_ | ~new_n24357_);
  assign new_n24356_ = (~new_n23700_ | new_n24359_ | new_n24357_) & (~new_n24358_ | ~new_n18189_ | ~new_n9749_ | ~new_n24357_);
  assign new_n24357_ = new_n15755_ & new_n16143_;
  assign new_n24358_ = new_n13316_ & (new_n13285_ | new_n13314_);
  assign new_n24359_ = new_n19677_ & (new_n19673_ | new_n19651_);
  assign new_n24360_ = (~new_n13038_ | new_n22939_) & (~new_n22175_ | ~new_n22933_ | ~new_n22939_);
  assign new_n24361_ = ~new_n16282_ & (~new_n17544_ | ~new_n19548_);
  assign new_n24362_ = new_n18189_ & ~new_n24358_ & new_n24357_;
  assign new_n24363_ = ~new_n23196_ & new_n10603_;
  assign new_n24364_ = new_n24365_ & (new_n24363_ | ~new_n24362_);
  assign new_n24365_ = new_n24357_ | ((~new_n24361_ | ~new_n24359_) & (new_n23700_ | new_n12188_ | new_n24359_));
  assign new_n24366_ = new_n24367_ ? (~new_n24506_ ^ new_n24518_) : (new_n24506_ ^ new_n24518_);
  assign new_n24367_ = new_n24368_ ? (~new_n24492_ ^ new_n24493_) : (new_n24492_ ^ new_n24493_);
  assign new_n24368_ = new_n24369_ ? (~new_n24383_ ^ new_n24253_) : (new_n24383_ ^ new_n24253_);
  assign new_n24369_ = ~new_n24370_ & new_n24381_;
  assign new_n24370_ = new_n24371_ & (new_n22534_ | ~new_n24373_ | (new_n24380_ ? new_n12717_ : ~new_n21704_));
  assign new_n24371_ = new_n24372_ & (new_n24379_ | new_n23963_ | new_n24373_) & (~new_n22534_ | new_n24378_ | ~new_n24373_);
  assign new_n24372_ = new_n24373_ | ~new_n23963_ | (new_n24375_ ? new_n24377_ : new_n24376_);
  assign new_n24373_ = new_n19040_ & new_n24374_;
  assign new_n24374_ = new_n10830_ & new_n10833_;
  assign new_n24375_ = ~new_n9893_ & new_n20252_;
  assign new_n24376_ = ~new_n22878_ & new_n20483_;
  assign new_n24377_ = new_n10204_ & (new_n10201_ | new_n10190_);
  assign new_n24378_ = new_n23935_ & ~new_n13318_ & ~new_n19638_;
  assign new_n24379_ = ~new_n12792_ & ~new_n23548_;
  assign new_n24380_ = new_n13909_ & new_n13889_ & new_n22876_;
  assign new_n24381_ = new_n24382_ & (new_n24373_ | ((new_n24375_ | ~new_n24376_ | ~new_n23963_) & (~new_n24379_ | new_n23963_)));
  assign new_n24382_ = ~new_n24373_ | (new_n22534_ ? ~new_n24378_ : (new_n24380_ ? ~new_n12717_ : new_n21704_));
  assign new_n24383_ = new_n24384_ ? (new_n24396_ ^ new_n24449_) : (~new_n24396_ ^ new_n24449_);
  assign new_n24384_ = new_n24385_ & (~new_n24391_ | ~new_n24394_ | (new_n20102_ ? new_n24395_ : new_n16417_));
  assign new_n24385_ = ~new_n24390_ & (new_n24394_ | (new_n24386_ & new_n14392_) | (new_n24389_ & ~new_n14392_));
  assign new_n24386_ = (new_n24387_ & ~new_n14884_) | (~new_n16313_ & new_n14884_ & (~new_n16305_ | new_n24388_));
  assign new_n24387_ = ~new_n8097_ & (~new_n8094_ | new_n10368_);
  assign new_n24388_ = ~new_n16283_ & ~new_n16316_;
  assign new_n24389_ = new_n15441_ ? new_n19649_ : new_n23324_;
  assign new_n24390_ = ~new_n24391_ & new_n24394_ & (new_n24393_ ? (new_n15530_ | new_n24392_) : ~new_n12006_);
  assign new_n24391_ = new_n7946_ & ~new_n8409_ & new_n7943_;
  assign new_n24392_ = new_n23553_ & new_n15528_;
  assign new_n24393_ = ~new_n16450_ & new_n16446_;
  assign new_n24394_ = ~new_n9827_ & (~new_n9823_ | ~new_n9799_ | ~new_n9830_);
  assign new_n24395_ = new_n21602_ & new_n6528_;
  assign new_n24396_ = new_n24397_ & (~new_n24408_ | ((new_n24447_ | ~new_n12442_ | ~new_n10837_) & (new_n24444_ | new_n10837_)));
  assign new_n24397_ = ~new_n24399_ & (new_n24408_ ? ~new_n24398_ : (~new_n24409_ | (~new_n7221_ & new_n18093_)));
  assign new_n24398_ = new_n10837_ & new_n7832_ & new_n7830_ & ~new_n12442_ & new_n7805_;
  assign new_n24399_ = ~new_n24408_ & ~new_n24409_ & (new_n22837_ ? new_n24401_ : new_n24400_);
  assign new_n24400_ = new_n7192_ & (new_n7164_ | ~new_n11616_);
  assign new_n24401_ = new_n24402_ & new_n24403_;
  assign new_n24402_ = ~new_n20408_ & ~new_n20436_;
  assign new_n24403_ = ~new_n20431_ & ~new_n24404_;
  assign new_n24404_ = ~new_n24405_ & (\all_features[3875]  | \all_features[3876]  | \all_features[3877]  | \all_features[3878]  | \all_features[3879] );
  assign new_n24405_ = ~new_n20430_ & (new_n20428_ | (~new_n20426_ & (new_n20411_ | (~new_n20413_ & ~new_n24406_))));
  assign new_n24406_ = ~new_n20415_ & (new_n20417_ | (new_n20424_ & (~new_n20420_ | (~new_n24407_ & new_n20422_))));
  assign new_n24407_ = ~\all_features[3877]  & \all_features[3878]  & \all_features[3879]  & (\all_features[3876]  ? new_n20421_ : (new_n20418_ | ~new_n20421_));
  assign new_n24408_ = new_n20436_ & (new_n20408_ | (new_n20431_ & new_n24404_));
  assign new_n24409_ = new_n24442_ & new_n24441_ & new_n24410_ & new_n24433_;
  assign new_n24410_ = ~new_n24432_ & (new_n24431_ | new_n24411_);
  assign new_n24411_ = ~new_n24424_ & (new_n24426_ | (~new_n24427_ & (new_n24428_ | (~new_n24412_ & ~new_n24429_))));
  assign new_n24412_ = ~new_n24413_ & (~new_n24423_ | (new_n24417_ & (~new_n24420_ | (~new_n24422_ & new_n24421_))));
  assign new_n24413_ = ~\all_features[1055]  & (~\all_features[1054]  | ~new_n24414_ | ~new_n24415_ | ~new_n24416_);
  assign new_n24414_ = \all_features[1048]  & \all_features[1049] ;
  assign new_n24415_ = \all_features[1052]  & \all_features[1053] ;
  assign new_n24416_ = \all_features[1050]  & \all_features[1051] ;
  assign new_n24417_ = \all_features[1055]  & (\all_features[1054]  | (\all_features[1053]  & (\all_features[1052]  | ~new_n24419_ | ~new_n24418_)));
  assign new_n24418_ = ~\all_features[1048]  & ~\all_features[1049] ;
  assign new_n24419_ = ~\all_features[1050]  & ~\all_features[1051] ;
  assign new_n24420_ = \all_features[1055]  & (\all_features[1054]  | (new_n24415_ & (\all_features[1050]  | \all_features[1051]  | \all_features[1049] )));
  assign new_n24421_ = \all_features[1054]  & \all_features[1055]  & (\all_features[1052]  | \all_features[1053]  | new_n24414_ | ~new_n24419_);
  assign new_n24422_ = \all_features[1054]  & \all_features[1055]  & (\all_features[1053]  | (~new_n24419_ & \all_features[1052] ));
  assign new_n24423_ = \all_features[1055]  & (\all_features[1053]  | \all_features[1054]  | \all_features[1052] );
  assign new_n24424_ = new_n24425_ & (~\all_features[1053]  | (~\all_features[1052]  & (~\all_features[1051]  | (~\all_features[1050]  & ~\all_features[1049] ))));
  assign new_n24425_ = ~\all_features[1054]  & ~\all_features[1055] ;
  assign new_n24426_ = new_n24425_ & (~\all_features[1051]  | ~new_n24415_ | (~\all_features[1050]  & ~new_n24414_));
  assign new_n24427_ = ~\all_features[1055]  & (~\all_features[1054]  | (~\all_features[1052]  & ~\all_features[1053]  & ~new_n24416_));
  assign new_n24428_ = ~\all_features[1055]  & (~\all_features[1054]  | (~\all_features[1053]  & (new_n24418_ | ~new_n24416_ | ~\all_features[1052] )));
  assign new_n24429_ = ~new_n24430_ & ~\all_features[1055] ;
  assign new_n24430_ = \all_features[1053]  & \all_features[1054]  & (\all_features[1052]  | (\all_features[1050]  & \all_features[1051]  & \all_features[1049] ));
  assign new_n24431_ = ~\all_features[1053]  & new_n24425_ & ((~\all_features[1050]  & new_n24418_) | ~\all_features[1052]  | ~\all_features[1051] );
  assign new_n24432_ = ~\all_features[1055]  & ~\all_features[1054]  & ~\all_features[1053]  & ~\all_features[1051]  & ~\all_features[1052] ;
  assign new_n24433_ = new_n24438_ & (~new_n24439_ | (~new_n24434_ & new_n24440_));
  assign new_n24434_ = new_n24435_ & ((~new_n24436_ & new_n24420_ & new_n24421_) | ~new_n24423_ | ~new_n24417_);
  assign new_n24435_ = ~new_n24429_ & ~new_n24413_;
  assign new_n24436_ = \all_features[1055]  & \all_features[1054]  & ~new_n24437_ & \all_features[1053] ;
  assign new_n24437_ = ~\all_features[1051]  & ~\all_features[1052]  & (~\all_features[1050]  | new_n24418_);
  assign new_n24438_ = ~new_n24431_ & ~new_n24432_;
  assign new_n24439_ = ~new_n24424_ & ~new_n24426_;
  assign new_n24440_ = ~new_n24427_ & ~new_n24428_;
  assign new_n24441_ = new_n24435_ & new_n24440_ & new_n24438_ & new_n24439_;
  assign new_n24442_ = new_n24438_ & new_n24439_ & (~new_n24435_ | ~new_n24440_ | (new_n24443_ & new_n24417_));
  assign new_n24443_ = new_n24423_ & new_n24420_ & new_n24421_;
  assign new_n24444_ = (~new_n21015_ & new_n24445_) | (new_n12536_ & new_n24446_ & ~new_n24445_);
  assign new_n24445_ = new_n10677_ & (new_n10679_ | new_n20086_);
  assign new_n24446_ = new_n7661_ & new_n7665_;
  assign new_n24447_ = new_n24448_ & new_n7581_;
  assign new_n24448_ = new_n7559_ & new_n7583_;
  assign new_n24449_ = new_n24453_ & (new_n24450_ | new_n24458_) & (new_n12190_ | new_n18911_ | new_n24491_ | ~new_n24458_);
  assign new_n24450_ = (~new_n24452_ | ~new_n10128_ | (new_n15918_ & ~new_n15555_)) & (~new_n17151_ | new_n24451_ | new_n10128_);
  assign new_n24451_ = new_n14090_ & new_n17804_;
  assign new_n24452_ = ~new_n7396_ & new_n7591_;
  assign new_n24453_ = ~new_n24458_ | ~new_n18911_ | ((~new_n24455_ | ~new_n14845_) & (new_n24454_ | new_n15990_ | new_n14845_));
  assign new_n24454_ = new_n17216_ & new_n15986_;
  assign new_n24455_ = ~new_n24456_ & new_n24457_;
  assign new_n24456_ = new_n23786_ & new_n23810_;
  assign new_n24457_ = ~new_n23815_ & ~new_n23818_;
  assign new_n24458_ = new_n24489_ & (new_n24482_ | new_n24459_);
  assign new_n24459_ = ~new_n24481_ & ~new_n24480_ & ~new_n24479_ & ~new_n24460_ & ~new_n24477_;
  assign new_n24460_ = new_n24461_ & new_n24466_ & (~new_n24474_ | ~new_n24476_ | ~new_n24471_ | ~new_n24473_);
  assign new_n24461_ = ~new_n24462_ & ~new_n24464_;
  assign new_n24462_ = ~\all_features[5215]  & (~\all_features[5214]  | (~\all_features[5212]  & ~\all_features[5213]  & ~new_n24463_));
  assign new_n24463_ = \all_features[5210]  & \all_features[5211] ;
  assign new_n24464_ = ~\all_features[5215]  & (~\all_features[5214]  | (~\all_features[5213]  & (new_n24465_ | ~\all_features[5212]  | ~new_n24463_)));
  assign new_n24465_ = ~\all_features[5208]  & ~\all_features[5209] ;
  assign new_n24466_ = ~new_n24467_ & ~new_n24469_;
  assign new_n24467_ = ~new_n24468_ & ~\all_features[5215] ;
  assign new_n24468_ = \all_features[5213]  & \all_features[5214]  & (\all_features[5212]  | (\all_features[5210]  & \all_features[5211]  & \all_features[5209] ));
  assign new_n24469_ = ~\all_features[5215]  & (~new_n24470_ | ~\all_features[5208]  | ~\all_features[5209]  | ~\all_features[5214]  | ~new_n24463_);
  assign new_n24470_ = \all_features[5212]  & \all_features[5213] ;
  assign new_n24471_ = \all_features[5215]  & (\all_features[5214]  | (\all_features[5213]  & (\all_features[5212]  | ~new_n24472_ | ~new_n24465_)));
  assign new_n24472_ = ~\all_features[5210]  & ~\all_features[5211] ;
  assign new_n24473_ = \all_features[5215]  & (\all_features[5214]  | (new_n24470_ & (\all_features[5210]  | \all_features[5211]  | \all_features[5209] )));
  assign new_n24474_ = new_n24475_ & (\all_features[5212]  | \all_features[5213]  | ~new_n24472_ | (\all_features[5209]  & \all_features[5208] ));
  assign new_n24475_ = \all_features[5214]  & \all_features[5215] ;
  assign new_n24476_ = \all_features[5215]  & (\all_features[5213]  | \all_features[5214]  | \all_features[5212] );
  assign new_n24477_ = ~\all_features[5213]  & new_n24478_ & ((~\all_features[5210]  & new_n24465_) | ~\all_features[5212]  | ~\all_features[5211] );
  assign new_n24478_ = ~\all_features[5214]  & ~\all_features[5215] ;
  assign new_n24479_ = new_n24478_ & (~\all_features[5213]  | (~\all_features[5212]  & (~\all_features[5211]  | (~\all_features[5210]  & ~\all_features[5209] ))));
  assign new_n24480_ = new_n24478_ & (~new_n24470_ | ~\all_features[5211]  | (~\all_features[5210]  & (~\all_features[5208]  | ~\all_features[5209] )));
  assign new_n24481_ = ~\all_features[5215]  & ~\all_features[5214]  & ~\all_features[5213]  & ~\all_features[5211]  & ~\all_features[5212] ;
  assign new_n24482_ = ~new_n24479_ & new_n24488_ & (new_n24480_ | (~new_n24486_ & new_n24461_ & new_n24483_));
  assign new_n24483_ = ~new_n24462_ & (new_n24464_ | (~new_n24467_ & (new_n24469_ | new_n24484_)));
  assign new_n24484_ = new_n24476_ & (~new_n24471_ | (new_n24473_ & (new_n24485_ | ~new_n24474_)));
  assign new_n24485_ = new_n24475_ & (\all_features[5213]  | (~new_n24472_ & \all_features[5212] ));
  assign new_n24486_ = new_n24466_ & ((~new_n24487_ & new_n24474_ & new_n24473_) | ~new_n24476_ | ~new_n24471_);
  assign new_n24487_ = new_n24475_ & \all_features[5213]  & ((~new_n24465_ & \all_features[5210] ) | \all_features[5212]  | \all_features[5211] );
  assign new_n24488_ = ~new_n24477_ & ~new_n24481_;
  assign new_n24489_ = new_n24490_ & ~new_n24480_ & ~new_n24464_ & ~new_n24479_;
  assign new_n24490_ = ~new_n24481_ & ~new_n24477_ & ~new_n24462_ & ~new_n24467_ & ~new_n24469_;
  assign new_n24491_ = new_n9827_ & (new_n9830_ | ~new_n9798_);
  assign new_n24492_ = ~new_n24326_ & new_n24254_;
  assign new_n24493_ = ~new_n24497_ & (~new_n24498_ | (new_n24494_ & ~new_n24505_) | (~new_n24495_ & new_n24505_));
  assign new_n24494_ = new_n19244_ ? (new_n7221_ | (~new_n18094_ & new_n7194_)) : new_n22354_;
  assign new_n24495_ = new_n16336_ & ~new_n18260_ & new_n24496_;
  assign new_n24496_ = ~new_n18285_ & ~new_n18288_;
  assign new_n24497_ = ~new_n24498_ & (new_n24504_ | new_n24503_) & (new_n7159_ | ~new_n15714_ | ~new_n16282_ | ~new_n24503_);
  assign new_n24498_ = new_n20635_ & (~new_n20657_ | (~new_n24499_ & ~new_n20660_ & ~new_n20655_));
  assign new_n24499_ = ~new_n20653_ & ~new_n20647_ & (new_n20645_ | new_n20651_ | new_n24500_);
  assign new_n24500_ = new_n20643_ & ~new_n24501_ & new_n20648_;
  assign new_n24501_ = ~new_n20639_ & new_n20641_ & \all_features[5702]  & \all_features[5703]  & (~\all_features[5701]  | new_n24502_);
  assign new_n24502_ = ~\all_features[5699]  & ~\all_features[5700]  & (~\all_features[5698]  | new_n20650_);
  assign new_n24503_ = ~new_n14810_ & new_n21485_;
  assign new_n24504_ = ~new_n22052_ & ~new_n22083_;
  assign new_n24505_ = new_n19813_ & (new_n19811_ | ~new_n22549_);
  assign new_n24506_ = ~new_n24507_ & ~new_n24517_;
  assign new_n24507_ = new_n24508_ & ((new_n22456_ & new_n14206_) | ~new_n24512_ | new_n24515_);
  assign new_n24508_ = new_n24509_ & (~new_n24513_ | (~new_n24203_ & new_n24514_) | (~new_n23834_ & ~new_n24514_));
  assign new_n24509_ = (~new_n24511_ | ~new_n24512_ | (~new_n22947_ & ~new_n21615_)) & (~new_n24067_ | new_n24510_ | new_n24512_);
  assign new_n24510_ = (new_n16375_ | ~new_n23200_) & (new_n16108_ | new_n16140_ | new_n23200_);
  assign new_n24511_ = new_n22456_ & new_n14206_;
  assign new_n24512_ = ~new_n7866_ & (~new_n7863_ | ~new_n7835_);
  assign new_n24513_ = ~new_n24512_ & ~new_n24067_;
  assign new_n24514_ = ~new_n20205_ & (~new_n20202_ | new_n20172_);
  assign new_n24515_ = (new_n24516_ & new_n23556_) | (new_n9749_ & ~new_n23556_ & (new_n9727_ | ~new_n9750_));
  assign new_n24516_ = ~new_n24446_ & new_n7636_;
  assign new_n24517_ = new_n24514_ & ~new_n24203_ & new_n24513_;
  assign new_n24518_ = ~new_n24539_ & new_n24519_;
  assign new_n24519_ = new_n24525_ & (new_n24534_ | new_n24520_);
  assign new_n24520_ = (new_n24523_ | new_n8434_ | ~new_n12447_ | (new_n8438_ & new_n8412_)) & (new_n24521_ | new_n12447_);
  assign new_n24521_ = new_n24522_ ? new_n23934_ : (~new_n14461_ & (~new_n14465_ | ~new_n14437_ | ~new_n14463_));
  assign new_n24522_ = new_n17815_ & ~new_n8412_ & ~new_n8434_;
  assign new_n24523_ = ~new_n24524_ & new_n8201_;
  assign new_n24524_ = new_n8227_ & new_n12192_;
  assign new_n24525_ = ~new_n24532_ & ~new_n24538_ & (~new_n24536_ | (~new_n24526_ & ~new_n24537_));
  assign new_n24526_ = ~new_n23921_ & new_n24527_;
  assign new_n24527_ = ~new_n24528_ & new_n23450_;
  assign new_n24528_ = ~new_n24529_ & (\all_features[2643]  | \all_features[2644]  | \all_features[2645]  | \all_features[2646]  | \all_features[2647] );
  assign new_n24529_ = ~new_n23468_ & (new_n23471_ | (~new_n23472_ & (new_n23474_ | (~new_n23473_ & ~new_n24530_))));
  assign new_n24530_ = ~new_n23461_ & (new_n23463_ | (new_n23466_ & (~new_n23465_ | (~new_n24531_ & new_n23454_))));
  assign new_n24531_ = ~\all_features[2645]  & \all_features[2646]  & \all_features[2647]  & (\all_features[2644]  ? new_n23458_ : (new_n23457_ | ~new_n23458_));
  assign new_n24532_ = new_n24533_ & (new_n24041_ ? new_n22389_ : ~new_n24535_);
  assign new_n24533_ = new_n23735_ & new_n24534_;
  assign new_n24534_ = ~new_n24448_ & ~new_n7581_;
  assign new_n24535_ = ~new_n10767_ & new_n10738_;
  assign new_n24536_ = ~new_n23735_ & new_n24534_;
  assign new_n24537_ = ~new_n24527_ & (~new_n23955_ | ~new_n14164_ | ~new_n12354_);
  assign new_n24538_ = new_n24523_ & new_n12447_ & ~new_n16850_ & ~new_n24534_;
  assign new_n24539_ = ~new_n24540_ & ~new_n24541_ & (new_n24537_ | ~new_n24536_ | new_n24526_);
  assign new_n24540_ = ~new_n24534_ & ((new_n23934_ & new_n24522_ & ~new_n12447_) | (new_n16850_ & new_n24523_ & new_n12447_));
  assign new_n24541_ = new_n24533_ & (new_n24041_ ? ~new_n22389_ : new_n24535_);
  assign new_n24542_ = ~new_n24543_ & new_n24554_;
  assign new_n24543_ = new_n24544_ & (new_n22988_ | ((new_n21617_ | ~new_n7509_ | new_n20579_) & (~new_n24141_ | ~new_n20579_)));
  assign new_n24544_ = new_n24545_ & ~new_n24548_ & (new_n10773_ | new_n14336_ | new_n22988_ | ~new_n20579_);
  assign new_n24545_ = (~new_n24546_ | new_n24547_ | ~new_n22988_) & (new_n20579_ | new_n7509_ | ~new_n6354_ | new_n22988_);
  assign new_n24546_ = new_n7635_ & new_n21684_;
  assign new_n24547_ = new_n17414_ & (new_n17392_ | ~new_n19638_);
  assign new_n24548_ = new_n21525_ & new_n24547_ & ~new_n24549_ & new_n22988_;
  assign new_n24549_ = new_n7798_ & (new_n7772_ | ~new_n24550_);
  assign new_n24550_ = ~new_n7799_ & (new_n7792_ | (~new_n7791_ & (new_n7787_ | (~new_n24551_ & ~new_n7789_))));
  assign new_n24551_ = ~new_n7782_ & (new_n7783_ | (~new_n7775_ & ~new_n24552_));
  assign new_n24552_ = ~new_n7777_ & (~new_n7797_ | (new_n7796_ & (~new_n7793_ | (~new_n24553_ & new_n7794_))));
  assign new_n24553_ = \all_features[3686]  & \all_features[3687]  & (\all_features[3685]  | (~new_n7795_ & \all_features[3684] ));
  assign new_n24554_ = new_n24555_ & (~new_n22988_ | ((new_n24557_ | ~new_n24547_) & (new_n21684_ | new_n14884_ | new_n24547_)));
  assign new_n24555_ = new_n22988_ | (new_n20579_ ? new_n24556_ : (new_n7509_ ? ~new_n21617_ : new_n6354_));
  assign new_n24556_ = new_n14336_ ? new_n21692_ : ~new_n10773_;
  assign new_n24557_ = (~new_n24549_ | ~new_n21525_) & (new_n15367_ | ~new_n24558_ | new_n21525_);
  assign new_n24558_ = ~new_n15396_ & ~new_n15399_;
  assign new_n24559_ = ~new_n24575_ & new_n24560_;
  assign new_n24560_ = new_n24571_ & (new_n18577_ | (new_n24561_ & (new_n15329_ | new_n18892_ | new_n20800_)));
  assign new_n24561_ = (~new_n24562_ | new_n20800_) & (new_n24564_ | ~new_n7866_ | ~new_n20800_ | (~new_n7863_ & ~new_n7834_));
  assign new_n24562_ = new_n24563_ & new_n15329_ & new_n9550_;
  assign new_n24563_ = new_n9579_ & new_n9581_;
  assign new_n24564_ = new_n24565_ & ~new_n8134_ & ~new_n24566_;
  assign new_n24565_ = ~new_n8159_ & ~new_n8161_;
  assign new_n24566_ = ~new_n8136_ & (new_n8139_ | (~new_n8151_ & (new_n8150_ | (~new_n24567_ & ~new_n8153_))));
  assign new_n24567_ = ~new_n8155_ & (new_n8157_ | (~new_n8156_ & (~new_n24570_ | new_n24568_)));
  assign new_n24568_ = \all_features[4559]  & ((~new_n24569_ & ~\all_features[4557]  & \all_features[4558] ) | (~new_n8145_ & (\all_features[4558]  | (~new_n8143_ & \all_features[4557] ))));
  assign new_n24569_ = (~\all_features[4554]  & ~\all_features[4555]  & ~\all_features[4556]  & (~\all_features[4553]  | ~\all_features[4552] )) | (\all_features[4556]  & (\all_features[4554]  | \all_features[4555] ));
  assign new_n24570_ = \all_features[4559]  & (\all_features[4557]  | \all_features[4558]  | \all_features[4556] );
  assign new_n24571_ = ~new_n18577_ | (new_n24572_ & (new_n24574_ | ~new_n18174_ | ~new_n21529_) & (new_n6533_ | new_n21529_));
  assign new_n24572_ = (new_n18174_ | new_n12264_ | ~new_n21529_) & (~new_n6533_ | ~new_n24573_ | new_n21529_);
  assign new_n24573_ = ~new_n24442_ & ~new_n24433_ & ~new_n24441_;
  assign new_n24574_ = ~new_n7804_ & new_n7832_;
  assign new_n24575_ = ~new_n24576_ & (new_n18577_ | ((new_n15329_ | ~new_n18892_ | new_n20800_) & (~new_n24564_ | ~new_n20800_)));
  assign new_n24576_ = new_n18577_ & new_n24574_ & new_n18174_ & new_n21529_;
  assign \o[36]  = new_n24578_ ^ new_n24579_;
  assign new_n24578_ = new_n23438_ & new_n24559_;
  assign new_n24579_ = new_n24580_ ? (new_n24581_ ^ new_n24631_) : (~new_n24581_ ^ new_n24631_);
  assign new_n24580_ = (~new_n24366_ & new_n24542_) | (~new_n23439_ & (~new_n24366_ | new_n24542_));
  assign new_n24581_ = new_n24582_ ? (new_n24583_ ^ new_n24618_) : (~new_n24583_ ^ new_n24618_);
  assign new_n24582_ = (~new_n24124_ & new_n24353_) | (~new_n23440_ & (~new_n24124_ | new_n24353_));
  assign new_n24583_ = new_n24584_ ? (new_n24585_ ^ new_n24605_) : (~new_n24585_ ^ new_n24605_);
  assign new_n24584_ = (~new_n23940_ & new_n24114_) | (~new_n23441_ & (~new_n23940_ | new_n24114_));
  assign new_n24585_ = new_n24586_ ? (new_n24587_ ^ new_n24598_) : (~new_n24587_ ^ new_n24598_);
  assign new_n24586_ = (~new_n23773_ & new_n23931_) | (~new_n23442_ & (~new_n23773_ | new_n23931_));
  assign new_n24587_ = new_n24588_ ? (new_n24589_ ^ new_n24594_) : (~new_n24589_ ^ new_n24594_);
  assign new_n24588_ = (new_n23601_ & new_n23659_) | (new_n23443_ & (new_n23601_ | new_n23659_));
  assign new_n24589_ = new_n24590_ ^ new_n24591_;
  assign new_n24590_ = new_n23444_ & new_n23599_;
  assign new_n24591_ = ~new_n24593_ & new_n24592_;
  assign new_n24592_ = ~new_n23655_ & new_n23602_;
  assign new_n24593_ = ~new_n23658_ & new_n23656_;
  assign new_n24594_ = new_n24595_ ? (new_n24596_ ^ new_n24597_) : (~new_n24596_ ^ new_n24597_);
  assign new_n24595_ = new_n24543_ & new_n24554_;
  assign new_n24596_ = new_n24560_ & new_n24575_;
  assign new_n24597_ = new_n23660_ & new_n23772_;
  assign new_n24598_ = new_n24599_ ? (~new_n24600_ ^ new_n24604_) : (new_n24600_ ^ new_n24604_);
  assign new_n24599_ = (new_n23958_ & new_n24003_) | (new_n23942_ & (new_n23958_ | new_n24003_));
  assign new_n24600_ = new_n24601_ ? (new_n24602_ ^ new_n24603_) : (~new_n24602_ ^ new_n24603_);
  assign new_n24601_ = new_n23775_ & new_n23824_;
  assign new_n24602_ = new_n24519_ & new_n24539_;
  assign new_n24603_ = new_n23884_ & new_n23928_;
  assign new_n24604_ = (new_n23828_ & new_n23883_) | (new_n23774_ & (new_n23828_ | new_n23883_));
  assign new_n24605_ = new_n24606_ ? (~new_n24616_ ^ new_n24617_) : (new_n24616_ ^ new_n24617_);
  assign new_n24606_ = new_n24607_ ? (new_n24611_ ^ new_n24615_) : (~new_n24611_ ^ new_n24615_);
  assign new_n24607_ = new_n24608_ ? (new_n24609_ ^ new_n24610_) : (~new_n24609_ ^ new_n24610_);
  assign new_n24608_ = new_n24329_ & new_n24343_;
  assign new_n24609_ = new_n23943_ & new_n23956_;
  assign new_n24610_ = new_n23959_ & new_n23999_;
  assign new_n24611_ = new_n24612_ ? (new_n24613_ ^ new_n24614_) : (~new_n24613_ ^ new_n24614_);
  assign new_n24612_ = ~new_n24517_ & new_n24507_;
  assign new_n24613_ = new_n24354_ & new_n24364_;
  assign new_n24614_ = new_n23829_ & new_n23881_;
  assign new_n24615_ = (new_n24211_ & new_n24212_) | (new_n24196_ & (new_n24211_ | new_n24212_));
  assign new_n24616_ = (~new_n24195_ & new_n24253_) | (~new_n24126_ & (~new_n24195_ | new_n24253_));
  assign new_n24617_ = (new_n23931_ & new_n24036_) | (~new_n23941_ & (new_n23931_ | new_n24036_));
  assign new_n24618_ = new_n24619_ ? (~new_n24629_ ^ new_n24630_) : (new_n24629_ ^ new_n24630_);
  assign new_n24619_ = new_n24620_ ? (~new_n24627_ ^ new_n24628_) : (new_n24627_ ^ new_n24628_);
  assign new_n24620_ = new_n24621_ ? (~new_n24625_ ^ new_n24626_) : (new_n24625_ ^ new_n24626_);
  assign new_n24621_ = new_n24622_ ? (new_n24623_ ^ new_n24624_) : (~new_n24623_ ^ new_n24624_);
  assign new_n24622_ = new_n24370_ & new_n24381_;
  assign new_n24623_ = new_n24128_ & new_n24146_;
  assign new_n24624_ = new_n24213_ & new_n24251_;
  assign new_n24625_ = (new_n24149_ & new_n24175_) | (new_n24127_ & (new_n24149_ | new_n24175_));
  assign new_n24626_ = (new_n24396_ & new_n24449_) | (new_n24384_ & (new_n24396_ | new_n24449_));
  assign new_n24627_ = (~new_n24383_ & new_n24253_) | (new_n24369_ & (~new_n24383_ | new_n24253_));
  assign new_n24628_ = new_n24150_ & new_n24172_;
  assign new_n24629_ = (new_n24328_ & new_n24349_) | (~new_n24125_ & (new_n24328_ | new_n24349_));
  assign new_n24630_ = (new_n24492_ & new_n24493_) | (~new_n24368_ & (new_n24492_ | new_n24493_));
  assign new_n24631_ = (new_n24506_ & new_n24518_) | (~new_n24367_ & (new_n24506_ | new_n24518_));
  assign \o[37]  = ~new_n24633_ ^ new_n24634_;
  assign new_n24633_ = new_n24578_ & new_n24579_;
  assign new_n24634_ = new_n24635_ ^ new_n24636_;
  assign new_n24635_ = (~new_n24581_ & new_n24631_) | (new_n24580_ & (~new_n24581_ | new_n24631_));
  assign new_n24636_ = new_n24637_ ? (~new_n24638_ ^ new_n24664_) : (new_n24638_ ^ new_n24664_);
  assign new_n24637_ = (~new_n24583_ & ~new_n24618_) | (new_n24582_ & (~new_n24583_ | ~new_n24618_));
  assign new_n24638_ = new_n24639_ ? (new_n24640_ ^ new_n24656_) : (~new_n24640_ ^ new_n24656_);
  assign new_n24639_ = (~new_n24585_ & ~new_n24605_) | (new_n24584_ & (~new_n24585_ | ~new_n24605_));
  assign new_n24640_ = new_n24641_ ? (new_n24642_ ^ new_n24652_) : (~new_n24642_ ^ new_n24652_);
  assign new_n24641_ = (~new_n24587_ & ~new_n24598_) | (new_n24586_ & (~new_n24587_ | ~new_n24598_));
  assign new_n24642_ = new_n24643_ ? (new_n24644_ ^ new_n24649_) : (~new_n24644_ ^ new_n24649_);
  assign new_n24643_ = (~new_n24589_ & ~new_n24594_) | (new_n24588_ & (~new_n24589_ | ~new_n24594_));
  assign new_n24644_ = ~new_n24645_ ^ new_n24646_;
  assign new_n24645_ = ~new_n24590_ & ~new_n24591_;
  assign new_n24646_ = new_n24647_ ^ new_n24648_;
  assign new_n24647_ = new_n24592_ & new_n24593_;
  assign new_n24648_ = new_n23554_ & new_n23445_ & new_n23599_;
  assign new_n24649_ = ~new_n24650_ ^ new_n24651_;
  assign new_n24650_ = (new_n24596_ & new_n24597_) | (new_n24595_ & (new_n24596_ | new_n24597_));
  assign new_n24651_ = (new_n24602_ & new_n24603_) | (new_n24601_ & (new_n24602_ | new_n24603_));
  assign new_n24652_ = new_n24653_ ? (new_n24654_ ^ new_n24655_) : (~new_n24654_ ^ new_n24655_);
  assign new_n24653_ = (~new_n24611_ & new_n24615_) | (~new_n24607_ & (~new_n24611_ | new_n24615_));
  assign new_n24654_ = (~new_n24600_ & new_n24604_) | (new_n24599_ & (~new_n24600_ | new_n24604_));
  assign new_n24655_ = (new_n24613_ & new_n24614_) | (new_n24612_ & (new_n24613_ | new_n24614_));
  assign new_n24656_ = new_n24657_ ? (~new_n24662_ ^ new_n24663_) : (new_n24662_ ^ new_n24663_);
  assign new_n24657_ = ~new_n24658_ ^ new_n24661_;
  assign new_n24658_ = new_n24659_ ^ new_n24660_;
  assign new_n24659_ = (new_n24609_ & new_n24610_) | (new_n24608_ & (new_n24609_ | new_n24610_));
  assign new_n24660_ = (new_n24623_ & new_n24624_) | (new_n24622_ & (new_n24623_ | new_n24624_));
  assign new_n24661_ = (new_n24625_ & new_n24626_) | (~new_n24621_ & (new_n24625_ | new_n24626_));
  assign new_n24662_ = (new_n24616_ & new_n24617_) | (~new_n24606_ & (new_n24616_ | new_n24617_));
  assign new_n24663_ = (new_n24627_ & new_n24628_) | (~new_n24620_ & (new_n24627_ | new_n24628_));
  assign new_n24664_ = (new_n24629_ & new_n24630_) | (~new_n24619_ & (new_n24629_ | new_n24630_));
  assign \o[38]  = ((new_n24666_ | new_n24667_) & (new_n24668_ ^ new_n24669_)) | (~new_n24666_ & ~new_n24667_ & (~new_n24668_ ^ new_n24669_));
  assign new_n24666_ = ~new_n24634_ & new_n24633_;
  assign new_n24667_ = ~new_n24636_ & new_n24635_;
  assign new_n24668_ = (~new_n24638_ & new_n24664_) | (new_n24637_ & (~new_n24638_ | new_n24664_));
  assign new_n24669_ = new_n24670_ ? (~new_n24671_ ^ new_n24683_) : (new_n24671_ ^ new_n24683_);
  assign new_n24670_ = (~new_n24640_ & ~new_n24656_) | (new_n24639_ & (~new_n24640_ | ~new_n24656_));
  assign new_n24671_ = new_n24672_ ? (new_n24673_ ^ new_n24679_) : (~new_n24673_ ^ new_n24679_);
  assign new_n24672_ = (~new_n24642_ & ~new_n24652_) | (new_n24641_ & (~new_n24642_ | ~new_n24652_));
  assign new_n24673_ = new_n24674_ ? (~new_n24675_ ^ new_n24678_) : (new_n24675_ ^ new_n24678_);
  assign new_n24674_ = (~new_n24644_ & ~new_n24649_) | (new_n24643_ & (~new_n24644_ | ~new_n24649_));
  assign new_n24675_ = new_n24676_ ^ new_n24677_;
  assign new_n24676_ = ~new_n24645_ & ~new_n24646_;
  assign new_n24677_ = ~new_n24647_ & ~new_n24648_;
  assign new_n24678_ = new_n24650_ & new_n24651_;
  assign new_n24679_ = new_n24680_ ? (new_n24681_ ^ new_n24682_) : (~new_n24681_ ^ new_n24682_);
  assign new_n24680_ = new_n24658_ & new_n24661_;
  assign new_n24681_ = (new_n24654_ & new_n24655_) | (new_n24653_ & (new_n24654_ | new_n24655_));
  assign new_n24682_ = new_n24659_ & new_n24660_;
  assign new_n24683_ = (new_n24662_ & new_n24663_) | (~new_n24657_ & (new_n24662_ | new_n24663_));
  assign \o[39]  = ~new_n24685_ ^ new_n24686_;
  assign new_n24685_ = (new_n24668_ | (~new_n24669_ & (new_n24667_ | new_n24666_))) & (new_n24667_ | new_n24666_ | ~new_n24669_);
  assign new_n24686_ = new_n24687_ ^ new_n24688_;
  assign new_n24687_ = (~new_n24671_ & new_n24683_) | (new_n24670_ & (~new_n24671_ | new_n24683_));
  assign new_n24688_ = new_n24689_ ? (~new_n24690_ ^ new_n24693_) : (new_n24690_ ^ new_n24693_);
  assign new_n24689_ = (~new_n24673_ & ~new_n24679_) | (new_n24672_ & (~new_n24673_ | ~new_n24679_));
  assign new_n24690_ = ~new_n24691_ ^ new_n24692_;
  assign new_n24691_ = (~new_n24675_ & new_n24678_) | (new_n24674_ & (~new_n24675_ | new_n24678_));
  assign new_n24692_ = ~new_n24677_ & new_n24676_;
  assign new_n24693_ = (new_n24681_ & new_n24682_) | (new_n24680_ & (new_n24681_ | new_n24682_));
  assign \o[40]  = ((new_n24695_ | new_n24696_) & (~new_n24697_ ^ new_n24698_)) | (~new_n24695_ & ~new_n24696_ & (new_n24697_ ^ new_n24698_));
  assign new_n24695_ = ~new_n24686_ & new_n24685_;
  assign new_n24696_ = ~new_n24688_ & new_n24687_;
  assign new_n24697_ = (~new_n24690_ & new_n24693_) | (new_n24689_ & (~new_n24690_ | new_n24693_));
  assign new_n24698_ = new_n24691_ & new_n24692_;
  assign \o[41]  = (new_n24698_ | new_n24695_ | new_n24696_) & (new_n24697_ | (new_n24698_ & (new_n24695_ | new_n24696_)));
  assign \o[42]  = new_n24701_ ? (~new_n25372_ ^ new_n25401_) : (new_n25372_ ^ new_n25401_);
  assign new_n24701_ = new_n24702_ ? (new_n25333_ ^ new_n25353_) : (~new_n25333_ ^ new_n25353_);
  assign new_n24702_ = new_n24703_ ? (new_n25222_ ^ new_n25322_) : (~new_n25222_ ^ new_n25322_);
  assign new_n24703_ = new_n24704_ ? (new_n25004_ ^ new_n25211_) : (~new_n25004_ ^ new_n25211_);
  assign new_n24704_ = new_n24705_ ? (new_n24961_ ^ new_n24997_) : (~new_n24961_ ^ new_n24997_);
  assign new_n24705_ = new_n24706_ ? (new_n24849_ ^ new_n24944_) : (~new_n24849_ ^ new_n24944_);
  assign new_n24706_ = new_n24707_ ^ new_n24786_;
  assign new_n24707_ = ~new_n24708_ & new_n24756_;
  assign new_n24708_ = new_n24709_ & ((~new_n24715_ & new_n14162_ & new_n24714_) | (new_n24711_ & ~new_n20489_));
  assign new_n24709_ = ~new_n24751_ & ~new_n24753_ & new_n24710_ & (~new_n24755_ | ~new_n14278_ | ~new_n24712_);
  assign new_n24710_ = (~new_n20489_ | ~new_n24711_) & (~new_n24714_ | (new_n14162_ ? ~new_n24715_ : ~new_n24750_));
  assign new_n24711_ = ~new_n14278_ & new_n24712_;
  assign new_n24712_ = ~new_n18812_ & new_n24713_;
  assign new_n24713_ = ~new_n15037_ & new_n17804_;
  assign new_n24714_ = ~new_n24713_ & ~new_n18812_;
  assign new_n24715_ = new_n24716_ & ~new_n24745_ & ~new_n24749_;
  assign new_n24716_ = new_n24744_ | (~new_n24743_ & ~new_n24717_ & new_n24738_);
  assign new_n24717_ = ~new_n24731_ & (new_n24733_ | (~new_n24734_ & (new_n24735_ | (~new_n24718_ & ~new_n24736_))));
  assign new_n24718_ = ~new_n24725_ & (~new_n24729_ | (new_n24719_ & (~new_n24728_ | (~new_n24730_ & new_n24722_))));
  assign new_n24719_ = \all_features[1071]  & (\all_features[1070]  | new_n24720_);
  assign new_n24720_ = \all_features[1069]  & (\all_features[1066]  | \all_features[1067]  | \all_features[1068]  | ~new_n24721_);
  assign new_n24721_ = ~\all_features[1064]  & ~\all_features[1065] ;
  assign new_n24722_ = \all_features[1071]  & ~new_n24723_ & \all_features[1070] ;
  assign new_n24723_ = ~\all_features[1069]  & ~\all_features[1068]  & ~\all_features[1067]  & ~new_n24724_ & ~\all_features[1066] ;
  assign new_n24724_ = \all_features[1064]  & \all_features[1065] ;
  assign new_n24725_ = ~\all_features[1071]  & (~\all_features[1070]  | ~new_n24724_ | ~new_n24726_ | ~new_n24727_);
  assign new_n24726_ = \all_features[1068]  & \all_features[1069] ;
  assign new_n24727_ = \all_features[1066]  & \all_features[1067] ;
  assign new_n24728_ = \all_features[1071]  & (\all_features[1070]  | (new_n24726_ & (\all_features[1066]  | \all_features[1067]  | \all_features[1065] )));
  assign new_n24729_ = \all_features[1071]  & (\all_features[1069]  | \all_features[1070]  | \all_features[1068] );
  assign new_n24730_ = \all_features[1070]  & \all_features[1071]  & (\all_features[1069]  | (\all_features[1068]  & (\all_features[1067]  | \all_features[1066] )));
  assign new_n24731_ = new_n24732_ & (~\all_features[1069]  | (~\all_features[1068]  & (~\all_features[1067]  | (~\all_features[1066]  & ~\all_features[1065] ))));
  assign new_n24732_ = ~\all_features[1070]  & ~\all_features[1071] ;
  assign new_n24733_ = new_n24732_ & (~\all_features[1067]  | ~new_n24726_ | (~\all_features[1066]  & ~new_n24724_));
  assign new_n24734_ = ~\all_features[1071]  & (~\all_features[1070]  | (~\all_features[1068]  & ~\all_features[1069]  & ~new_n24727_));
  assign new_n24735_ = ~\all_features[1071]  & (~\all_features[1070]  | (~\all_features[1069]  & (new_n24721_ | ~new_n24727_ | ~\all_features[1068] )));
  assign new_n24736_ = ~new_n24737_ & ~\all_features[1071] ;
  assign new_n24737_ = \all_features[1069]  & \all_features[1070]  & (\all_features[1068]  | (\all_features[1066]  & \all_features[1067]  & \all_features[1065] ));
  assign new_n24738_ = new_n24742_ & (new_n24735_ | new_n24734_ | (~new_n24739_ & ~new_n24736_ & ~new_n24725_));
  assign new_n24739_ = new_n24729_ & ~new_n24740_ & new_n24719_;
  assign new_n24740_ = ~new_n24723_ & new_n24728_ & \all_features[1070]  & \all_features[1071]  & (~\all_features[1069]  | new_n24741_);
  assign new_n24741_ = ~\all_features[1067]  & ~\all_features[1068]  & (~\all_features[1066]  | new_n24721_);
  assign new_n24742_ = ~new_n24731_ & ~new_n24733_;
  assign new_n24743_ = ~\all_features[1069]  & new_n24732_ & ((~\all_features[1066]  & new_n24721_) | ~\all_features[1068]  | ~\all_features[1067] );
  assign new_n24744_ = ~\all_features[1071]  & ~\all_features[1070]  & ~\all_features[1069]  & ~\all_features[1067]  & ~\all_features[1068] ;
  assign new_n24745_ = new_n24742_ & new_n24747_ & (new_n24746_ | new_n24735_ | new_n24725_ | ~new_n24748_);
  assign new_n24746_ = new_n24729_ & new_n24728_ & new_n24719_ & new_n24722_;
  assign new_n24747_ = ~new_n24743_ & ~new_n24744_;
  assign new_n24748_ = ~new_n24734_ & ~new_n24736_;
  assign new_n24749_ = new_n24747_ & new_n24742_ & new_n24748_ & ~new_n24735_ & ~new_n24725_;
  assign new_n24750_ = new_n18775_ & new_n18780_ & ~new_n18771_ & ~new_n18782_ & ~new_n18770_;
  assign new_n24751_ = new_n18812_ & new_n23869_ & ~new_n24752_ & ~new_n15745_;
  assign new_n24752_ = ~new_n7407_ & (~new_n7396_ | ~new_n7405_);
  assign new_n24753_ = new_n24752_ & new_n18812_ & new_n14846_ & new_n24754_;
  assign new_n24754_ = ~new_n10648_ & new_n22838_;
  assign new_n24755_ = new_n13475_ & (~new_n18154_ | ~new_n13451_);
  assign new_n24756_ = ~new_n24757_ & (~new_n18812_ | (~new_n15745_ & new_n23869_ & ~new_n24752_) | (new_n24758_ & new_n24752_));
  assign new_n24757_ = new_n24714_ & ~new_n14162_ & ~new_n24750_;
  assign new_n24758_ = new_n24754_ ? new_n14846_ : ~new_n24759_;
  assign new_n24759_ = ~new_n24760_ & ~new_n24784_;
  assign new_n24760_ = new_n24778_ & ~new_n24783_ & ~new_n24761_ & ~new_n24782_;
  assign new_n24761_ = ~new_n24776_ & ~new_n24777_ & new_n24771_ & (~new_n24765_ | ~new_n24762_);
  assign new_n24762_ = \all_features[863]  & (\all_features[862]  | new_n24763_);
  assign new_n24763_ = \all_features[861]  & (\all_features[858]  | \all_features[859]  | \all_features[860]  | ~new_n24764_);
  assign new_n24764_ = ~\all_features[856]  & ~\all_features[857] ;
  assign new_n24765_ = new_n24770_ & new_n24766_ & new_n24768_;
  assign new_n24766_ = \all_features[863]  & (\all_features[862]  | (new_n24767_ & (\all_features[858]  | \all_features[859]  | \all_features[857] )));
  assign new_n24767_ = \all_features[860]  & \all_features[861] ;
  assign new_n24768_ = \all_features[863]  & ~new_n24769_ & \all_features[862] ;
  assign new_n24769_ = ~\all_features[858]  & ~\all_features[859]  & ~\all_features[860]  & ~\all_features[861]  & (~\all_features[857]  | ~\all_features[856] );
  assign new_n24770_ = \all_features[863]  & (\all_features[861]  | \all_features[862]  | \all_features[860] );
  assign new_n24771_ = ~new_n24772_ & ~new_n24774_;
  assign new_n24772_ = ~new_n24773_ & ~\all_features[863] ;
  assign new_n24773_ = \all_features[861]  & \all_features[862]  & (\all_features[860]  | (\all_features[858]  & \all_features[859]  & \all_features[857] ));
  assign new_n24774_ = ~\all_features[863]  & (~\all_features[862]  | (~\all_features[860]  & ~\all_features[861]  & ~new_n24775_));
  assign new_n24775_ = \all_features[858]  & \all_features[859] ;
  assign new_n24776_ = ~\all_features[863]  & (~\all_features[862]  | (~\all_features[861]  & (new_n24764_ | ~new_n24775_ | ~\all_features[860] )));
  assign new_n24777_ = ~\all_features[863]  & (~new_n24775_ | ~\all_features[856]  | ~\all_features[857]  | ~\all_features[862]  | ~new_n24767_);
  assign new_n24778_ = ~new_n24779_ & ~new_n24781_;
  assign new_n24779_ = ~\all_features[861]  & new_n24780_ & ((~\all_features[858]  & new_n24764_) | ~\all_features[860]  | ~\all_features[859] );
  assign new_n24780_ = ~\all_features[862]  & ~\all_features[863] ;
  assign new_n24781_ = ~\all_features[863]  & ~\all_features[862]  & ~\all_features[861]  & ~\all_features[859]  & ~\all_features[860] ;
  assign new_n24782_ = new_n24780_ & (~\all_features[861]  | (~\all_features[860]  & (~\all_features[859]  | (~\all_features[858]  & ~\all_features[857] ))));
  assign new_n24783_ = new_n24780_ & (~new_n24767_ | ~\all_features[859]  | (~\all_features[858]  & (~\all_features[856]  | ~\all_features[857] )));
  assign new_n24784_ = new_n24778_ & new_n24771_ & new_n24785_ & ~new_n24776_ & ~new_n24777_;
  assign new_n24785_ = ~new_n24782_ & ~new_n24783_;
  assign new_n24786_ = ~new_n24787_ & new_n24847_;
  assign new_n24787_ = new_n24788_ & new_n24807_ & ((new_n24804_ & new_n24805_) | (~new_n24811_ & new_n24846_));
  assign new_n24788_ = new_n24789_ & (new_n24805_ | new_n24806_ | ~new_n24804_);
  assign new_n24789_ = (new_n6603_ | ~new_n24790_ | ~new_n24803_) & (~new_n24802_ | ~new_n24801_);
  assign new_n24790_ = ~new_n24793_ & new_n24791_;
  assign new_n24791_ = new_n16815_ & new_n24792_;
  assign new_n24792_ = ~new_n16840_ & ~new_n16844_;
  assign new_n24793_ = ~new_n14568_ & ~new_n14552_ & (new_n14567_ | new_n24794_);
  assign new_n24794_ = new_n24800_ & (new_n14561_ | (~new_n14554_ & new_n24795_ & (new_n14557_ | new_n24798_)));
  assign new_n24795_ = ~new_n14557_ & ~new_n14559_ & (~new_n14574_ | ~new_n14569_ | new_n24796_);
  assign new_n24796_ = new_n14571_ & ~new_n24797_ & new_n14572_;
  assign new_n24797_ = new_n14573_ & \all_features[557]  & ((~new_n14556_ & \all_features[554] ) | \all_features[556]  | \all_features[555] );
  assign new_n24798_ = ~new_n14559_ & (~new_n14574_ | (new_n14569_ & (~new_n14571_ | (~new_n24799_ & new_n14572_))));
  assign new_n24799_ = new_n14573_ & (\all_features[557]  | (~new_n14570_ & \all_features[556] ));
  assign new_n24800_ = ~new_n14566_ & ~new_n14563_ & ~new_n14565_;
  assign new_n24801_ = ~new_n24451_ & ~new_n24791_;
  assign new_n24802_ = ~new_n14162_ & new_n16026_;
  assign new_n24803_ = ~new_n8083_ & new_n8093_;
  assign new_n24804_ = ~new_n24791_ & new_n24451_;
  assign new_n24805_ = new_n13367_ & (~new_n15530_ | (~new_n15528_ & new_n15497_));
  assign new_n24806_ = ~new_n13367_ & (~new_n15860_ | new_n19832_);
  assign new_n24807_ = (~new_n24809_ | ~new_n24801_) & (new_n24810_ | ~new_n24808_);
  assign new_n24808_ = ~new_n24803_ & new_n24790_;
  assign new_n24809_ = new_n16813_ & ~new_n15822_ & new_n14162_;
  assign new_n24810_ = new_n11373_ & new_n22952_;
  assign new_n24811_ = (~new_n24812_ & ~new_n23832_) | (~new_n24814_ & new_n24841_ & new_n23832_);
  assign new_n24812_ = new_n9313_ & new_n24813_;
  assign new_n24813_ = ~new_n9341_ & ~new_n15043_;
  assign new_n24814_ = ~new_n24840_ & (~new_n24833_ | (~new_n24838_ & (new_n24831_ | new_n24839_ | ~new_n24815_)));
  assign new_n24815_ = ~new_n24827_ & ~new_n24825_ & ((~new_n24822_ & new_n24816_) | ~new_n24830_ | ~new_n24829_);
  assign new_n24816_ = \all_features[535]  & \all_features[534]  & ~new_n24819_ & new_n24817_;
  assign new_n24817_ = \all_features[535]  & (\all_features[534]  | (new_n24818_ & (\all_features[530]  | \all_features[531]  | \all_features[529] )));
  assign new_n24818_ = \all_features[532]  & \all_features[533] ;
  assign new_n24819_ = new_n24821_ & ~\all_features[533]  & ~new_n24820_ & ~\all_features[532] ;
  assign new_n24820_ = \all_features[528]  & \all_features[529] ;
  assign new_n24821_ = ~\all_features[530]  & ~\all_features[531] ;
  assign new_n24822_ = \all_features[535]  & \all_features[534]  & ~new_n24823_ & \all_features[533] ;
  assign new_n24823_ = ~\all_features[531]  & ~\all_features[532]  & (~\all_features[530]  | new_n24824_);
  assign new_n24824_ = ~\all_features[528]  & ~\all_features[529] ;
  assign new_n24825_ = ~new_n24826_ & ~\all_features[535] ;
  assign new_n24826_ = \all_features[533]  & \all_features[534]  & (\all_features[532]  | (\all_features[530]  & \all_features[531]  & \all_features[529] ));
  assign new_n24827_ = ~\all_features[535]  & (~\all_features[534]  | ~new_n24828_ | ~new_n24820_ | ~new_n24818_);
  assign new_n24828_ = \all_features[530]  & \all_features[531] ;
  assign new_n24829_ = \all_features[535]  & (\all_features[534]  | (\all_features[533]  & (\all_features[532]  | ~new_n24821_ | ~new_n24824_)));
  assign new_n24830_ = \all_features[535]  & (\all_features[533]  | \all_features[534]  | \all_features[532] );
  assign new_n24831_ = ~new_n24825_ & (new_n24827_ | (new_n24830_ & (~new_n24829_ | (~new_n24832_ & new_n24817_))));
  assign new_n24832_ = ~\all_features[533]  & \all_features[534]  & \all_features[535]  & (\all_features[532]  ? new_n24821_ : (new_n24820_ | ~new_n24821_));
  assign new_n24833_ = ~new_n24837_ & ~new_n24834_ & ~new_n24836_;
  assign new_n24834_ = new_n24835_ & (~\all_features[533]  | (~\all_features[532]  & (~\all_features[531]  | (~\all_features[530]  & ~\all_features[529] ))));
  assign new_n24835_ = ~\all_features[534]  & ~\all_features[535] ;
  assign new_n24836_ = ~\all_features[533]  & new_n24835_ & ((~\all_features[530]  & new_n24824_) | ~\all_features[532]  | ~\all_features[531] );
  assign new_n24837_ = new_n24835_ & (~\all_features[531]  | ~new_n24818_ | (~\all_features[530]  & ~new_n24820_));
  assign new_n24838_ = ~\all_features[535]  & (~\all_features[534]  | (~\all_features[532]  & ~\all_features[533]  & ~new_n24828_));
  assign new_n24839_ = ~\all_features[535]  & (~\all_features[534]  | (~\all_features[533]  & (new_n24824_ | ~\all_features[532]  | ~new_n24828_)));
  assign new_n24840_ = ~\all_features[535]  & ~\all_features[534]  & ~\all_features[533]  & ~\all_features[531]  & ~\all_features[532] ;
  assign new_n24841_ = new_n24834_ | ~new_n24844_ | ((new_n24825_ | ~new_n24845_) & (new_n24842_ | new_n24837_));
  assign new_n24842_ = new_n24843_ & (~new_n24816_ | ~new_n24829_ | ~new_n24830_);
  assign new_n24843_ = ~new_n24827_ & ~new_n24825_ & ~new_n24838_ & ~new_n24839_;
  assign new_n24844_ = ~new_n24836_ & ~new_n24840_;
  assign new_n24845_ = ~new_n24837_ & ~new_n24827_ & ~new_n24838_ & ~new_n24839_;
  assign new_n24846_ = new_n24791_ & new_n24793_;
  assign new_n24847_ = new_n24848_ & (~new_n24810_ | ~new_n24808_) & (~new_n24806_ | ~new_n24804_);
  assign new_n24848_ = (~new_n24846_ | ~new_n24811_) & (new_n24802_ | new_n24809_ | ~new_n24801_);
  assign new_n24849_ = new_n24850_ ? (new_n24901_ ^ new_n24918_) : (~new_n24901_ ^ new_n24918_);
  assign new_n24850_ = ~new_n24851_ & new_n24899_;
  assign new_n24851_ = new_n24852_ & ((~new_n7269_ & new_n7226_ & new_n24857_) | (new_n24896_ & new_n24898_));
  assign new_n24852_ = new_n24853_ & (~new_n24896_ | (~new_n24895_ & ~new_n24897_) | (~new_n23088_ & new_n24897_));
  assign new_n24853_ = ~new_n24856_ & ~new_n24893_ & (~new_n24894_ | ~new_n14846_ | new_n24854_);
  assign new_n24854_ = new_n24855_ & new_n8132_;
  assign new_n24855_ = ~new_n19130_ & new_n20871_;
  assign new_n24856_ = new_n24857_ & (new_n7269_ ? new_n24892_ : ~new_n7226_);
  assign new_n24857_ = ~new_n14846_ & new_n24858_;
  assign new_n24858_ = ~new_n24890_ & ~new_n24887_ & ~new_n24859_ & ~new_n24881_;
  assign new_n24859_ = ~new_n24860_ & ~new_n24880_;
  assign new_n24860_ = ~new_n24874_ & (new_n24876_ | (~new_n24877_ & (new_n24878_ | (~new_n24861_ & ~new_n24879_))));
  assign new_n24861_ = ~new_n24862_ & (new_n24864_ | (new_n24873_ & (~new_n24868_ | (~new_n24872_ & new_n24871_))));
  assign new_n24862_ = ~new_n24863_ & ~\all_features[1319] ;
  assign new_n24863_ = \all_features[1317]  & \all_features[1318]  & (\all_features[1316]  | (\all_features[1314]  & \all_features[1315]  & \all_features[1313] ));
  assign new_n24864_ = ~\all_features[1319]  & (~\all_features[1318]  | ~new_n24865_ | ~new_n24866_ | ~new_n24867_);
  assign new_n24865_ = \all_features[1312]  & \all_features[1313] ;
  assign new_n24866_ = \all_features[1316]  & \all_features[1317] ;
  assign new_n24867_ = \all_features[1314]  & \all_features[1315] ;
  assign new_n24868_ = \all_features[1319]  & (\all_features[1318]  | (\all_features[1317]  & (\all_features[1316]  | ~new_n24870_ | ~new_n24869_)));
  assign new_n24869_ = ~\all_features[1312]  & ~\all_features[1313] ;
  assign new_n24870_ = ~\all_features[1314]  & ~\all_features[1315] ;
  assign new_n24871_ = \all_features[1319]  & (\all_features[1318]  | (new_n24866_ & (\all_features[1314]  | \all_features[1315]  | \all_features[1313] )));
  assign new_n24872_ = ~\all_features[1317]  & \all_features[1318]  & \all_features[1319]  & (\all_features[1316]  ? new_n24870_ : (new_n24865_ | ~new_n24870_));
  assign new_n24873_ = \all_features[1319]  & (\all_features[1317]  | \all_features[1318]  | \all_features[1316] );
  assign new_n24874_ = ~\all_features[1317]  & new_n24875_ & ((~\all_features[1314]  & new_n24869_) | ~\all_features[1316]  | ~\all_features[1315] );
  assign new_n24875_ = ~\all_features[1318]  & ~\all_features[1319] ;
  assign new_n24876_ = new_n24875_ & (~\all_features[1317]  | (~\all_features[1316]  & (~\all_features[1315]  | (~\all_features[1314]  & ~\all_features[1313] ))));
  assign new_n24877_ = new_n24875_ & (~\all_features[1315]  | ~new_n24866_ | (~\all_features[1314]  & ~new_n24865_));
  assign new_n24878_ = ~\all_features[1319]  & (~\all_features[1318]  | (~\all_features[1316]  & ~\all_features[1317]  & ~new_n24867_));
  assign new_n24879_ = ~\all_features[1319]  & (~\all_features[1318]  | (~\all_features[1317]  & (new_n24869_ | ~new_n24867_ | ~\all_features[1316] )));
  assign new_n24880_ = ~\all_features[1319]  & ~\all_features[1318]  & ~\all_features[1317]  & ~\all_features[1315]  & ~\all_features[1316] ;
  assign new_n24881_ = ~new_n24874_ & ~new_n24880_ & (~new_n24886_ | (~new_n24882_ & ~new_n24878_ & ~new_n24879_));
  assign new_n24882_ = ~new_n24862_ & ~new_n24864_ & (~new_n24873_ | ~new_n24868_ | new_n24883_);
  assign new_n24883_ = new_n24871_ & new_n24884_ & (new_n24885_ | ~\all_features[1317]  | ~\all_features[1318]  | ~\all_features[1319] );
  assign new_n24884_ = \all_features[1318]  & \all_features[1319]  & (\all_features[1316]  | \all_features[1317]  | new_n24865_ | ~new_n24870_);
  assign new_n24885_ = ~\all_features[1315]  & ~\all_features[1316]  & (~\all_features[1314]  | new_n24869_);
  assign new_n24886_ = ~new_n24876_ & ~new_n24877_;
  assign new_n24887_ = ~new_n24880_ & ~new_n24877_ & ~new_n24876_ & ~new_n24888_ & ~new_n24874_;
  assign new_n24888_ = new_n24889_ & (~new_n24884_ | ~new_n24873_ | ~new_n24868_ | ~new_n24871_);
  assign new_n24889_ = ~new_n24864_ & ~new_n24862_ & ~new_n24878_ & ~new_n24879_;
  assign new_n24890_ = new_n24891_ & new_n24886_ & ~new_n24862_ & ~new_n24879_ & ~new_n24874_ & ~new_n24878_;
  assign new_n24891_ = ~new_n24864_ & ~new_n24880_;
  assign new_n24892_ = ~new_n17844_ & new_n14337_;
  assign new_n24893_ = new_n23592_ & ~new_n13838_ & ~new_n24858_ & ~new_n14846_ & ~new_n23170_;
  assign new_n24894_ = ~new_n23581_ & (~new_n23558_ | ~new_n23584_ | ~new_n23588_);
  assign new_n24895_ = new_n10204_ & (new_n10201_ | ~new_n10168_);
  assign new_n24896_ = ~new_n24894_ & new_n14846_;
  assign new_n24897_ = ~new_n18985_ & (~new_n18962_ | new_n23549_);
  assign new_n24898_ = ~new_n23088_ & new_n24897_;
  assign new_n24899_ = new_n14846_ ? new_n24900_ : ((new_n24892_ | ~new_n7269_ | ~new_n24858_) & (new_n23592_ | new_n24858_));
  assign new_n24900_ = (~new_n24854_ | ~new_n24894_) & (new_n24895_ | new_n24897_ | new_n24894_);
  assign new_n24901_ = ~new_n24902_ & new_n24914_;
  assign new_n24902_ = new_n24912_ & new_n24903_ & (~new_n24755_ | new_n24908_ | ~new_n24907_);
  assign new_n24903_ = new_n12728_ | ((~new_n19773_ | ~new_n24906_ | new_n24387_) & (new_n24904_ | ~new_n24387_));
  assign new_n24904_ = (new_n7409_ & (~new_n7434_ | ~new_n7438_)) ? new_n24905_ : new_n9686_;
  assign new_n24905_ = ~new_n20730_ & new_n14923_;
  assign new_n24906_ = ~new_n15265_ & new_n21625_;
  assign new_n24907_ = ~new_n14162_ & new_n12728_;
  assign new_n24908_ = new_n22278_ & (new_n20918_ | (~new_n20916_ & (new_n20919_ | new_n24909_)));
  assign new_n24909_ = ~new_n20920_ & (new_n20911_ | (~new_n20913_ & (new_n20909_ | (~new_n24910_ & ~new_n20914_))));
  assign new_n24910_ = new_n20904_ & (~new_n20905_ | (new_n20902_ & (new_n24911_ | ~new_n20899_)));
  assign new_n24911_ = \all_features[782]  & \all_features[783]  & (\all_features[781]  | (\all_features[780]  & (\all_features[779]  | \all_features[778] )));
  assign new_n24912_ = ~new_n12728_ | ~new_n14162_ | (new_n7803_ ? new_n24913_ : ~new_n11337_);
  assign new_n24913_ = ~new_n10999_ & (~new_n13324_ | ~new_n10977_);
  assign new_n24914_ = new_n24915_ & (~new_n24907_ | (~new_n24908_ & new_n24755_) | (new_n19843_ & ~new_n24755_));
  assign new_n24915_ = (new_n24916_ | ~new_n14162_ | ~new_n12728_) & (new_n24387_ | ~new_n24917_ | new_n12728_);
  assign new_n24916_ = new_n7803_ ? ~new_n24913_ : new_n11337_;
  assign new_n24917_ = new_n24906_ ? ~new_n19773_ : ~new_n21964_;
  assign new_n24918_ = ~new_n24919_ & ~new_n24943_;
  assign new_n24919_ = new_n24922_ & ~new_n24940_ & ~new_n24920_ & ~new_n24939_;
  assign new_n24920_ = new_n24921_ & new_n24924_;
  assign new_n24921_ = new_n12756_ & ~new_n24923_ & new_n24922_;
  assign new_n24922_ = new_n15164_ & ~new_n14047_ & ~new_n14070_;
  assign new_n24923_ = ~new_n13271_ & new_n13244_;
  assign new_n24924_ = new_n24938_ | ~new_n24927_;
  assign new_n24925_ = ~\all_features[823]  & (~\all_features[822]  | new_n24926_);
  assign new_n24926_ = ~\all_features[821]  & (~\all_features[819]  | ~\all_features[820]  | ~\all_features[818]  | (~\all_features[817]  & ~\all_features[816] ));
  assign new_n24927_ = \all_features[822]  | \all_features[823]  | (~new_n24928_ & \all_features[821]  & new_n24930_);
  assign new_n24928_ = ~\all_features[820]  & (~\all_features[819]  | (~\all_features[818]  & ~\all_features[817] ));
  assign new_n24930_ = \all_features[819]  & \all_features[820]  & \all_features[821]  & (\all_features[818]  | (\all_features[817]  & \all_features[816] ));
  assign new_n24931_ = ~\all_features[823]  & (~new_n24932_ | (~\all_features[820]  & (~\all_features[818]  | ~\all_features[819]  | ~\all_features[817] )));
  assign new_n24932_ = \all_features[821]  & ~\all_features[823]  & \all_features[822] ;
  assign new_n24933_ = ~\all_features[823]  & (~\all_features[822]  | ~new_n24934_ | ~\all_features[820]  | ~\all_features[821] );
  assign new_n24934_ = \all_features[819]  & \all_features[818]  & \all_features[816]  & \all_features[817] ;
  assign new_n24938_ = ~\all_features[823]  & ~\all_features[822]  & ~\all_features[821]  & ~\all_features[819]  & ~\all_features[820] ;
  assign new_n24939_ = ~new_n12756_ & ~new_n24923_ & ~new_n13523_;
  assign new_n24940_ = new_n24923_ & new_n24922_ & (new_n24496_ | new_n20494_);
  assign new_n24943_ = ~new_n24924_ & new_n24921_;
  assign new_n24944_ = new_n24945_ & new_n24959_;
  assign new_n24945_ = new_n24956_ & new_n24946_ & new_n24949_ & (~new_n24958_ | ~new_n24957_);
  assign new_n24946_ = new_n24791_ | ((new_n24947_ | ~new_n24948_) & (new_n24023_ | ~new_n12864_ | new_n24948_));
  assign new_n24947_ = new_n18178_ & ~new_n18099_ & ~new_n12747_;
  assign new_n24948_ = new_n22899_ & new_n22922_;
  assign new_n24949_ = (~new_n24951_ | new_n24952_) & (~new_n24950_ | (new_n12864_ ? ~new_n24023_ : new_n24954_));
  assign new_n24950_ = ~new_n24791_ & ~new_n24948_;
  assign new_n24951_ = new_n24791_ & ~new_n16812_ & ~new_n23117_;
  assign new_n24952_ = ~new_n10833_ & (~new_n10830_ | new_n24953_);
  assign new_n24953_ = ~new_n19041_ & ~new_n10805_;
  assign new_n24954_ = new_n21855_ & new_n24955_;
  assign new_n24955_ = ~new_n21882_ & ~new_n21886_;
  assign new_n24956_ = ~new_n24791_ | ((new_n23218_ | ~new_n16812_) & (new_n18259_ | new_n18288_ | ~new_n23117_ | new_n16812_));
  assign new_n24957_ = ~new_n15920_ & ~new_n15953_;
  assign new_n24958_ = new_n24791_ & new_n16812_ & new_n23218_;
  assign new_n24959_ = new_n24960_ & (~new_n24958_ | new_n24957_);
  assign new_n24960_ = (new_n12864_ | ~new_n24950_ | ~new_n24954_) & (~new_n24952_ | ~new_n24951_);
  assign new_n24961_ = new_n24962_ ? (~new_n24944_ ^ new_n24988_) : (new_n24944_ ^ new_n24988_);
  assign new_n24962_ = new_n24963_ ? (new_n24978_ ^ new_n24982_) : (~new_n24978_ ^ new_n24982_);
  assign new_n24963_ = ~new_n24964_ & new_n24976_;
  assign new_n24964_ = ~new_n24965_ & new_n24969_ & (new_n21690_ | ~new_n21198_ | ~new_n24974_);
  assign new_n24965_ = new_n24966_ & (new_n9652_ ? new_n24967_ : new_n24968_);
  assign new_n24966_ = ~new_n19039_ & new_n21690_;
  assign new_n24967_ = ~new_n6591_ | (~new_n6569_ & new_n11061_);
  assign new_n24968_ = new_n16363_ & new_n20115_;
  assign new_n24969_ = (new_n21198_ | new_n21690_ | (~new_n24971_ & ~new_n24970_)) & (~new_n19039_ | new_n24972_ | ~new_n21690_);
  assign new_n24970_ = new_n11621_ & new_n17414_;
  assign new_n24971_ = ~new_n9422_ & ~new_n11621_;
  assign new_n24972_ = (new_n7097_ & new_n18288_) | (~new_n16101_ & new_n24973_ & ~new_n18288_);
  assign new_n24973_ = ~new_n16067_ & ~new_n16098_;
  assign new_n24974_ = new_n24975_ ? new_n6638_ : ~new_n23088_;
  assign new_n24975_ = new_n6448_ & (new_n6456_ | new_n6427_);
  assign new_n24976_ = new_n24977_ & (~new_n24966_ | (new_n24967_ & new_n9652_) | (new_n24968_ & ~new_n9652_));
  assign new_n24977_ = new_n21690_ | ((new_n24974_ | ~new_n21198_) & (new_n24971_ | new_n24970_ | new_n21198_));
  assign new_n24978_ = new_n19339_ ? new_n24979_ : ((~new_n24716_ & new_n24981_ & ~new_n18950_) | (new_n24980_ & new_n18950_));
  assign new_n24979_ = (new_n23765_ | ~new_n23122_ | new_n23771_) & (~new_n23771_ | (new_n22707_ ? new_n22796_ : ~new_n13976_));
  assign new_n24980_ = (~new_n11379_ & new_n13845_) ? new_n19343_ : new_n11699_;
  assign new_n24981_ = new_n24745_ & new_n24749_;
  assign new_n24982_ = ~new_n24983_ & ~new_n24987_;
  assign new_n24983_ = new_n11272_ & ((~new_n24984_ & ~new_n24985_ & ~new_n24791_) | (new_n14988_ & new_n7868_ & new_n24791_));
  assign new_n24984_ = ~new_n11615_ & new_n19195_;
  assign new_n24985_ = new_n11615_ & new_n24986_;
  assign new_n24986_ = ~new_n22633_ & (~new_n22635_ | ~new_n22611_);
  assign new_n24987_ = new_n11272_ & new_n11615_ & ~new_n24791_ & ~new_n24986_;
  assign new_n24988_ = new_n24989_ & (new_n24996_ | ~new_n19778_ | ~new_n24995_ | ~new_n13196_);
  assign new_n24989_ = (~new_n24992_ & ~new_n24990_ & new_n24995_) | (~new_n24995_ & (new_n6533_ ? ~new_n24993_ : new_n24455_));
  assign new_n24990_ = new_n24402_ & ~new_n24855_ & ~new_n24991_;
  assign new_n24991_ = new_n19778_ & new_n13196_;
  assign new_n24992_ = ~new_n24991_ & ~new_n24402_ & ~new_n21880_ & (~new_n21856_ | new_n24955_);
  assign new_n24993_ = new_n24994_ & ~new_n21251_ & ~new_n24792_;
  assign new_n24994_ = new_n16816_ & new_n16838_;
  assign new_n24995_ = new_n12933_ & (new_n12910_ | (new_n12936_ & new_n12940_));
  assign new_n24996_ = (~new_n10240_ & new_n12444_ & ~new_n13242_) | (new_n13242_ & (new_n19381_ | ~new_n15171_));
  assign new_n24997_ = new_n24998_ & new_n25000_ & (new_n16278_ | new_n24445_ | new_n22550_ | ~new_n13804_);
  assign new_n24998_ = ~new_n24999_ & (new_n13922_ | ~new_n22550_ | (new_n14786_ ? new_n15320_ : ~new_n20309_));
  assign new_n24999_ = new_n16840_ & new_n24994_ & ~new_n22550_ & ~new_n16278_ & ~new_n13804_;
  assign new_n25000_ = ~new_n25002_ & (new_n25001_ | new_n22550_ | ~new_n16278_);
  assign new_n25001_ = (new_n12453_ & ~new_n9550_ & new_n12373_) | (new_n16948_ & new_n12687_ & (new_n9550_ | ~new_n12373_));
  assign new_n25002_ = new_n13922_ & new_n22550_ & (new_n25003_ ? ~new_n13367_ : ~new_n18750_);
  assign new_n25003_ = new_n7101_ & ~new_n10609_ & new_n7098_;
  assign new_n25004_ = new_n25005_ ? (~new_n25149_ ^ new_n25202_) : (new_n25149_ ^ new_n25202_);
  assign new_n25005_ = new_n25006_ ? (new_n25072_ ^ new_n25143_) : (~new_n25072_ ^ new_n25143_);
  assign new_n25006_ = new_n25007_ ? (new_n25027_ ^ new_n25038_) : (~new_n25027_ ^ new_n25038_);
  assign new_n25007_ = ~new_n25008_ & new_n25025_;
  assign new_n25008_ = new_n25009_ & new_n25023_ & (~new_n17248_ | ~new_n25024_);
  assign new_n25009_ = new_n15318_ ? ((new_n25014_ | new_n25017_) & (~new_n8541_ | ~new_n25016_ | ~new_n25017_)) : new_n25010_;
  assign new_n25010_ = (new_n25011_ | ~new_n25012_ | (new_n19766_ & new_n19764_)) & (~new_n6389_ | new_n25013_ | new_n25012_);
  assign new_n25011_ = new_n6908_ & (new_n6886_ | new_n13805_);
  assign new_n25012_ = ~new_n14625_ & ~new_n13242_;
  assign new_n25013_ = new_n14210_ & new_n14182_ & new_n14207_;
  assign new_n25014_ = (new_n6448_ & (new_n6427_ | (new_n6450_ & new_n6456_))) ? ~new_n23218_ : ~new_n25015_;
  assign new_n25015_ = new_n24927_ & ~new_n24938_ & ~new_n24933_ & ~new_n24925_ & ~new_n24931_;
  assign new_n25016_ = new_n10240_ & (new_n10238_ | ~new_n10207_);
  assign new_n25017_ = new_n21278_ & (new_n21252_ | (new_n21274_ & new_n25018_));
  assign new_n25018_ = ~new_n21272_ & (new_n21273_ | (~new_n21270_ & (new_n21268_ | (~new_n21263_ & ~new_n25019_))));
  assign new_n25019_ = ~new_n21266_ & (new_n21261_ | (~new_n21265_ & (~new_n25022_ | new_n25020_)));
  assign new_n25020_ = \all_features[1287]  & ((~new_n25021_ & ~\all_features[1285]  & \all_features[1286] ) | (~new_n21258_ & (\all_features[1286]  | (~new_n21255_ & \all_features[1285] ))));
  assign new_n25021_ = (~\all_features[1282]  & ~\all_features[1283]  & ~\all_features[1284]  & (~\all_features[1281]  | ~\all_features[1280] )) | (\all_features[1284]  & (\all_features[1282]  | \all_features[1283] ));
  assign new_n25022_ = \all_features[1287]  & (\all_features[1285]  | \all_features[1286]  | \all_features[1284] );
  assign new_n25023_ = (new_n6389_ | new_n25012_ | new_n15318_) & (new_n25016_ | ~new_n25017_ | ~new_n15318_);
  assign new_n25024_ = new_n25012_ & ~new_n15318_ & new_n25011_;
  assign new_n25025_ = ~new_n25026_ & (~new_n15318_ | ((new_n8541_ | ~new_n25016_ | ~new_n25017_) & (~new_n25014_ | new_n25017_)));
  assign new_n25026_ = ~new_n17248_ & new_n25024_;
  assign new_n25027_ = ~new_n25036_ & new_n25028_;
  assign new_n25028_ = ~new_n25029_ & new_n25033_;
  assign new_n25029_ = ~new_n22937_ & new_n25030_;
  assign new_n25030_ = ~new_n25031_ & ~new_n21964_;
  assign new_n25031_ = ~new_n23857_ & (~new_n23835_ | ~new_n25032_);
  assign new_n25032_ = new_n23863_ & new_n23859_;
  assign new_n25033_ = new_n21964_ ? ((~new_n25034_ | ~new_n25035_ | new_n14242_) & (new_n19026_ | ~new_n14242_)) : ~new_n25031_;
  assign new_n25034_ = ~new_n10399_ & ~new_n8484_;
  assign new_n25035_ = new_n18991_ & new_n19017_;
  assign new_n25036_ = new_n25037_ & (~new_n22937_ | ~new_n25030_);
  assign new_n25037_ = ~new_n21964_ | ((new_n13243_ | ~new_n19026_ | ~new_n14242_) & (new_n14242_ | (new_n25035_ & new_n25034_)));
  assign new_n25038_ = ~new_n25070_ & new_n25039_;
  assign new_n25039_ = ~new_n25040_ & (new_n23640_ | ((new_n25061_ | ~new_n25062_ | ~new_n25060_) & (new_n25058_ | new_n25060_)));
  assign new_n25040_ = new_n6604_ & new_n23640_ & (new_n23832_ ? (new_n25057_ | new_n25041_) : ~new_n8985_);
  assign new_n25041_ = new_n25053_ & ~new_n25056_ & ~new_n25042_ & ~new_n25054_;
  assign new_n25042_ = ~new_n25043_ & ~new_n25046_ & ~new_n25048_ & (~new_n25050_ | (~new_n25052_ & ~\all_features[4878] ));
  assign new_n25043_ = ~\all_features[4879]  & (~\all_features[4878]  | (~\all_features[4877]  & (new_n25045_ | ~\all_features[4876]  | ~new_n25044_)));
  assign new_n25044_ = \all_features[4874]  & \all_features[4875] ;
  assign new_n25045_ = ~\all_features[4872]  & ~\all_features[4873] ;
  assign new_n25046_ = ~\all_features[4879]  & (~\all_features[4873]  | ~new_n25044_ | ~new_n25047_ | ~\all_features[4872] );
  assign new_n25047_ = \all_features[4878]  & \all_features[4876]  & \all_features[4877] ;
  assign new_n25048_ = ~\all_features[4879]  & (~\all_features[4878]  | ~\all_features[4877]  | (~new_n25049_ & ~\all_features[4876] ));
  assign new_n25049_ = \all_features[4875]  & \all_features[4873]  & \all_features[4874] ;
  assign new_n25050_ = \all_features[4878]  & \all_features[4879]  & (\all_features[4876]  | \all_features[4877]  | \all_features[4875]  | ~new_n25051_);
  assign new_n25051_ = ~\all_features[4874]  & (~\all_features[4873]  | ~\all_features[4872] );
  assign new_n25052_ = \all_features[4876]  & \all_features[4877]  & (\all_features[4875]  | \all_features[4874]  | \all_features[4873] );
  assign new_n25053_ = \all_features[4878]  | \all_features[4879]  | (~new_n25051_ & \all_features[4877]  & \all_features[4876]  & \all_features[4875] );
  assign new_n25054_ = ~\all_features[4877]  & new_n25055_ & ((~\all_features[4874]  & new_n25045_) | ~\all_features[4876]  | ~\all_features[4875] );
  assign new_n25055_ = ~\all_features[4878]  & ~\all_features[4879] ;
  assign new_n25056_ = new_n25055_ & (~\all_features[4877]  | (~\all_features[4876]  & (~\all_features[4875]  | (~\all_features[4874]  & ~\all_features[4873] ))));
  assign new_n25057_ = new_n25053_ & ~new_n25048_ & ~new_n25056_ & ~new_n25046_ & ~new_n25043_ & ~new_n25054_;
  assign new_n25058_ = (~new_n25059_ & new_n14330_ & new_n22365_) | (~new_n22365_ & (new_n7477_ | new_n7475_));
  assign new_n25059_ = new_n10801_ & new_n14331_;
  assign new_n25060_ = ~new_n24410_ & new_n24573_;
  assign new_n25061_ = new_n7000_ & new_n20097_ & new_n6998_;
  assign new_n25062_ = ~new_n25066_ & new_n24759_ & (new_n24781_ | (~new_n25063_ & ~new_n24779_));
  assign new_n25063_ = ~new_n24782_ & (new_n24783_ | (~new_n24774_ & (new_n24776_ | (~new_n24772_ & ~new_n25064_))));
  assign new_n25064_ = ~new_n24777_ & (~new_n24770_ | (new_n24762_ & (~new_n24766_ | (~new_n25065_ & new_n24768_))));
  assign new_n25065_ = \all_features[862]  & \all_features[863]  & (\all_features[861]  | (\all_features[860]  & (\all_features[859]  | \all_features[858] )));
  assign new_n25066_ = new_n24778_ & (~new_n24785_ | (~new_n25067_ & ~new_n24774_ & ~new_n24776_));
  assign new_n25067_ = ~new_n24777_ & ~new_n24772_ & (~new_n24770_ | new_n25068_ | ~new_n24762_);
  assign new_n25068_ = ~new_n24769_ & new_n24766_ & \all_features[862]  & \all_features[863]  & (~\all_features[861]  | new_n25069_);
  assign new_n25069_ = ~\all_features[859]  & ~\all_features[860]  & (~\all_features[858]  | new_n24764_);
  assign new_n25070_ = ~new_n6604_ & new_n23640_ & ((new_n9375_ & new_n22606_) ? ~new_n15030_ : ~new_n25071_);
  assign new_n25071_ = new_n15265_ & (new_n21636_ | (new_n21626_ & new_n24206_));
  assign new_n25072_ = new_n25073_ ? (new_n25106_ ^ new_n25140_) : (~new_n25106_ ^ new_n25140_);
  assign new_n25073_ = new_n25074_ & (new_n14337_ ? (~new_n25077_ | new_n25104_) : new_n25081_);
  assign new_n25074_ = ~new_n25075_ & (~new_n25078_ | ~new_n25079_) & (new_n16333_ | new_n14337_ | ~new_n25080_ | new_n25079_);
  assign new_n25075_ = new_n8595_ & new_n14337_ & ~new_n25076_ & ~new_n25077_;
  assign new_n25076_ = new_n7039_ & (new_n7036_ | new_n7003_);
  assign new_n25077_ = new_n23948_ & ~new_n22501_ & ~new_n23949_;
  assign new_n25078_ = new_n12447_ & ~new_n13328_ & ~new_n14337_;
  assign new_n25079_ = new_n18334_ & new_n20440_;
  assign new_n25080_ = new_n12717_ & new_n12709_;
  assign new_n25081_ = (~new_n25082_ | new_n25079_) & (new_n12447_ | ~new_n19048_ | ~new_n25079_);
  assign new_n25082_ = new_n25101_ & new_n25103_ & new_n25096_ & ~new_n25080_ & ~new_n25083_;
  assign new_n25083_ = ~new_n25095_ & ~new_n25094_ & ~new_n25092_ & ~new_n25084_ & ~new_n25090_;
  assign new_n25084_ = \all_features[2071]  & \all_features[2070]  & ~new_n25087_ & new_n25085_;
  assign new_n25085_ = \all_features[2071]  & (\all_features[2070]  | (new_n25086_ & (\all_features[2066]  | \all_features[2067]  | \all_features[2065] )));
  assign new_n25086_ = \all_features[2068]  & \all_features[2069] ;
  assign new_n25087_ = ~\all_features[2069]  & ~\all_features[2068]  & ~\all_features[2067]  & ~new_n25088_ & ~\all_features[2066] ;
  assign new_n25088_ = \all_features[2064]  & \all_features[2065] ;
  assign new_n25089_ = \all_features[2069]  & (\all_features[2065]  | \all_features[2066]  | \all_features[2067]  | \all_features[2068]  | \all_features[2064] );
  assign new_n25090_ = ~\all_features[2071]  & (~\all_features[2070]  | new_n25091_);
  assign new_n25091_ = ~\all_features[2069]  & (~\all_features[2067]  | ~\all_features[2068]  | ~\all_features[2066]  | (~\all_features[2065]  & ~\all_features[2064] ));
  assign new_n25092_ = ~new_n25093_ & ~\all_features[2071] ;
  assign new_n25093_ = \all_features[2069]  & \all_features[2070]  & (\all_features[2068]  | (\all_features[2066]  & \all_features[2067]  & \all_features[2065] ));
  assign new_n25094_ = ~\all_features[2071]  & (~new_n25088_ | ~\all_features[2066]  | ~\all_features[2067]  | ~\all_features[2070]  | ~new_n25086_);
  assign new_n25095_ = ~\all_features[2071]  & (~\all_features[2070]  | (~\all_features[2069]  & ~\all_features[2068]  & (~\all_features[2067]  | ~\all_features[2066] )));
  assign new_n25096_ = new_n25097_ & new_n25101_ & ~new_n25095_ & ~new_n25099_ & ~new_n25090_ & ~new_n25092_;
  assign new_n25097_ = ~new_n25094_ & (new_n25098_ | \all_features[2070]  | \all_features[2071] );
  assign new_n25098_ = new_n25086_ & \all_features[2067]  & (\all_features[2066]  | new_n25088_);
  assign new_n25099_ = ~\all_features[2071]  & ~new_n25100_ & ~\all_features[2070] ;
  assign new_n25100_ = \all_features[2069]  & (\all_features[2068]  | (\all_features[2067]  & (\all_features[2066]  | \all_features[2065] )));
  assign new_n25101_ = \all_features[2069]  | \all_features[2070]  | \all_features[2071]  | (\all_features[2068]  & \all_features[2067]  & ~new_n25102_);
  assign new_n25102_ = ~\all_features[2066]  & ~\all_features[2064]  & ~\all_features[2065] ;
  assign new_n25103_ = \all_features[2070]  | \all_features[2071]  | (new_n25100_ & new_n25098_);
  assign new_n25104_ = new_n25105_ ? (~new_n23032_ & (~new_n23003_ | ~new_n23025_ | ~new_n23594_)) : ~new_n7066_;
  assign new_n25105_ = ~new_n20785_ & new_n19434_;
  assign new_n25106_ = new_n14163_ ? new_n25107_ : ((new_n25111_ | new_n25137_ | ~new_n23450_) & (new_n25109_ | new_n23450_));
  assign new_n25107_ = (new_n25076_ | new_n25108_) & (new_n17898_ | ~new_n13807_ | ~new_n25108_);
  assign new_n25108_ = ~new_n23630_ & (~new_n23608_ | ~new_n23632_ | ~new_n23636_);
  assign new_n25109_ = (~new_n25110_ & ~new_n17840_) ? new_n18594_ : new_n17624_;
  assign new_n25110_ = new_n17817_ & new_n20160_;
  assign new_n25111_ = ~new_n25112_ & ~new_n25136_;
  assign new_n25112_ = new_n25130_ & (new_n25134_ | (~new_n25135_ & new_n25113_ & (new_n25122_ | new_n25128_)));
  assign new_n25113_ = ~new_n25122_ & ~new_n25124_ & (~new_n25127_ | ~new_n25126_ | new_n25114_);
  assign new_n25114_ = new_n25115_ & ~new_n25120_ & new_n25117_;
  assign new_n25115_ = \all_features[1327]  & (\all_features[1326]  | (new_n25116_ & (\all_features[1322]  | \all_features[1323]  | \all_features[1321] )));
  assign new_n25116_ = \all_features[1324]  & \all_features[1325] ;
  assign new_n25117_ = new_n25119_ & (\all_features[1324]  | \all_features[1325]  | ~new_n25118_ | (\all_features[1321]  & \all_features[1320] ));
  assign new_n25118_ = ~\all_features[1322]  & ~\all_features[1323] ;
  assign new_n25119_ = \all_features[1326]  & \all_features[1327] ;
  assign new_n25120_ = new_n25119_ & \all_features[1325]  & ((~new_n25121_ & \all_features[1322] ) | \all_features[1324]  | \all_features[1323] );
  assign new_n25121_ = ~\all_features[1320]  & ~\all_features[1321] ;
  assign new_n25122_ = ~new_n25123_ & ~\all_features[1327] ;
  assign new_n25123_ = \all_features[1325]  & \all_features[1326]  & (\all_features[1324]  | (\all_features[1322]  & \all_features[1323]  & \all_features[1321] ));
  assign new_n25124_ = ~\all_features[1327]  & (~new_n25116_ | ~\all_features[1320]  | ~\all_features[1321]  | ~\all_features[1326]  | ~new_n25125_);
  assign new_n25125_ = \all_features[1322]  & \all_features[1323] ;
  assign new_n25126_ = \all_features[1327]  & (\all_features[1326]  | (\all_features[1325]  & (\all_features[1324]  | ~new_n25118_ | ~new_n25121_)));
  assign new_n25127_ = \all_features[1327]  & (\all_features[1325]  | \all_features[1326]  | \all_features[1324] );
  assign new_n25128_ = ~new_n25124_ & (~new_n25127_ | (new_n25126_ & (~new_n25115_ | (~new_n25129_ & new_n25117_))));
  assign new_n25129_ = new_n25119_ & (\all_features[1325]  | (~new_n25118_ & \all_features[1324] ));
  assign new_n25130_ = \all_features[1326]  | \all_features[1327]  | (~new_n25133_ & new_n25132_ & \all_features[1325] );
  assign new_n25132_ = new_n25116_ & \all_features[1323]  & (\all_features[1322]  | (\all_features[1320]  & \all_features[1321] ));
  assign new_n25133_ = ~\all_features[1324]  & (~\all_features[1323]  | (~\all_features[1322]  & ~\all_features[1321] ));
  assign new_n25134_ = ~\all_features[1327]  & (~\all_features[1326]  | (~\all_features[1324]  & ~\all_features[1325]  & ~new_n25125_));
  assign new_n25135_ = ~\all_features[1327]  & (~\all_features[1326]  | (~\all_features[1325]  & (new_n25121_ | ~\all_features[1324]  | ~new_n25125_)));
  assign new_n25136_ = ~\all_features[1327]  & ~\all_features[1326]  & ~\all_features[1325]  & ~\all_features[1323]  & ~\all_features[1324] ;
  assign new_n25137_ = ~new_n25136_ & new_n25130_;
  assign new_n25140_ = new_n11272_ & (new_n25141_ | (~new_n7602_ & ~new_n10682_ & new_n21692_));
  assign new_n25141_ = new_n7602_ & ((~new_n12980_ & (new_n14045_ | ~new_n12978_)) ? ~new_n25142_ : new_n16762_);
  assign new_n25142_ = ~new_n20265_ & ~new_n12624_;
  assign new_n25143_ = (new_n23188_ | new_n25147_ | ~new_n25148_) & (new_n25148_ | (new_n7732_ ? new_n25144_ : new_n25145_));
  assign new_n25144_ = (new_n17391_ & new_n19638_) ? new_n10677_ : ~new_n22548_;
  assign new_n25145_ = new_n25146_ ? new_n18751_ : ~new_n18381_;
  assign new_n25146_ = new_n17215_ & new_n15958_;
  assign new_n25147_ = ~new_n22940_ & new_n21245_;
  assign new_n25148_ = new_n13471_ & new_n13467_ & new_n13476_ & ~new_n13464_ & ~new_n13474_;
  assign new_n25149_ = ~new_n25150_ & new_n25200_;
  assign new_n25150_ = new_n25151_ & (~new_n25198_ | ~new_n25196_) & (~new_n25197_ | ~new_n24563_);
  assign new_n25151_ = new_n25152_ & (new_n25163_ | ~new_n25162_) & (~new_n25160_ | ~new_n25159_);
  assign new_n25152_ = ~new_n25153_ & (new_n18953_ | ~new_n25158_ | ~new_n25157_ | (new_n18951_ & new_n18941_));
  assign new_n25153_ = ~new_n18914_ & new_n25154_ & (~new_n12301_ | ~new_n12298_ | new_n12268_);
  assign new_n25154_ = ~new_n25156_ & new_n25155_;
  assign new_n25155_ = new_n7736_ & (new_n7733_ | new_n19130_);
  assign new_n25156_ = ~new_n19822_ & new_n23072_;
  assign new_n25157_ = ~new_n25155_ & new_n25146_;
  assign new_n25158_ = new_n16411_ & new_n11896_;
  assign new_n25159_ = ~new_n25155_ & ~new_n25146_;
  assign new_n25160_ = (~new_n24855_ | ~new_n20115_) & (new_n16900_ | ~new_n25161_ | new_n20115_);
  assign new_n25161_ = new_n7830_ & new_n7832_;
  assign new_n25162_ = new_n25155_ & new_n25156_;
  assign new_n25163_ = (~new_n25077_ & new_n15753_ & new_n15596_) | (~new_n25164_ & new_n25191_ & (~new_n15753_ | ~new_n15596_));
  assign new_n25164_ = ~new_n25190_ & (~new_n25183_ | (~new_n25188_ & (new_n25181_ | new_n25189_ | ~new_n25165_)));
  assign new_n25165_ = ~new_n25177_ & ~new_n25175_ & ((~new_n25172_ & new_n25166_) | ~new_n25180_ | ~new_n25179_);
  assign new_n25166_ = \all_features[767]  & \all_features[766]  & ~new_n25169_ & new_n25167_;
  assign new_n25167_ = \all_features[767]  & (\all_features[766]  | (new_n25168_ & (\all_features[762]  | \all_features[763]  | \all_features[761] )));
  assign new_n25168_ = \all_features[764]  & \all_features[765] ;
  assign new_n25169_ = new_n25171_ & ~\all_features[765]  & ~new_n25170_ & ~\all_features[764] ;
  assign new_n25170_ = \all_features[760]  & \all_features[761] ;
  assign new_n25171_ = ~\all_features[762]  & ~\all_features[763] ;
  assign new_n25172_ = \all_features[767]  & \all_features[766]  & ~new_n25173_ & \all_features[765] ;
  assign new_n25173_ = ~\all_features[763]  & ~\all_features[764]  & (~\all_features[762]  | new_n25174_);
  assign new_n25174_ = ~\all_features[760]  & ~\all_features[761] ;
  assign new_n25175_ = ~new_n25176_ & ~\all_features[767] ;
  assign new_n25176_ = \all_features[765]  & \all_features[766]  & (\all_features[764]  | (\all_features[762]  & \all_features[763]  & \all_features[761] ));
  assign new_n25177_ = ~\all_features[767]  & (~\all_features[766]  | ~new_n25178_ | ~new_n25170_ | ~new_n25168_);
  assign new_n25178_ = \all_features[762]  & \all_features[763] ;
  assign new_n25179_ = \all_features[767]  & (\all_features[766]  | (\all_features[765]  & (\all_features[764]  | ~new_n25171_ | ~new_n25174_)));
  assign new_n25180_ = \all_features[767]  & (\all_features[765]  | \all_features[766]  | \all_features[764] );
  assign new_n25181_ = ~new_n25175_ & (new_n25177_ | (new_n25180_ & (~new_n25179_ | (~new_n25182_ & new_n25167_))));
  assign new_n25182_ = ~\all_features[765]  & \all_features[766]  & \all_features[767]  & (\all_features[764]  ? new_n25171_ : (new_n25170_ | ~new_n25171_));
  assign new_n25183_ = ~new_n25187_ & ~new_n25184_ & ~new_n25186_;
  assign new_n25184_ = new_n25185_ & (~\all_features[765]  | (~\all_features[764]  & (~\all_features[763]  | (~\all_features[762]  & ~\all_features[761] ))));
  assign new_n25185_ = ~\all_features[766]  & ~\all_features[767] ;
  assign new_n25186_ = ~\all_features[765]  & new_n25185_ & ((~\all_features[762]  & new_n25174_) | ~\all_features[764]  | ~\all_features[763] );
  assign new_n25187_ = new_n25185_ & (~\all_features[763]  | ~new_n25168_ | (~\all_features[762]  & ~new_n25170_));
  assign new_n25188_ = ~\all_features[767]  & (~\all_features[766]  | (~\all_features[764]  & ~\all_features[765]  & ~new_n25178_));
  assign new_n25189_ = ~\all_features[767]  & (~\all_features[766]  | (~\all_features[765]  & (new_n25174_ | ~\all_features[764]  | ~new_n25178_)));
  assign new_n25190_ = ~\all_features[767]  & ~\all_features[766]  & ~\all_features[765]  & ~\all_features[763]  & ~\all_features[764] ;
  assign new_n25191_ = new_n25184_ | ~new_n25194_ | ((new_n25175_ | ~new_n25195_) & (new_n25192_ | new_n25187_));
  assign new_n25192_ = new_n25193_ & (~new_n25166_ | ~new_n25179_ | ~new_n25180_);
  assign new_n25193_ = ~new_n25177_ & ~new_n25175_ & ~new_n25188_ & ~new_n25189_;
  assign new_n25194_ = ~new_n25186_ & ~new_n25190_;
  assign new_n25195_ = ~new_n25187_ & ~new_n25177_ & ~new_n25188_ & ~new_n25189_;
  assign new_n25196_ = ~new_n25158_ & new_n25157_;
  assign new_n25197_ = new_n25154_ & new_n18914_;
  assign new_n25198_ = ~new_n25199_ & new_n18950_;
  assign new_n25199_ = ~new_n18920_ & ~new_n18941_;
  assign new_n25200_ = new_n25201_ & (new_n24563_ | ~new_n25197_);
  assign new_n25201_ = (new_n25198_ | ~new_n25196_) & (~new_n25163_ | ~new_n25162_) & (new_n25160_ | ~new_n25159_);
  assign new_n25202_ = new_n25204_ & (new_n25203_ | new_n13804_ | new_n25206_);
  assign new_n25203_ = new_n7269_ ? new_n22275_ : (~new_n11333_ | (~new_n11335_ & new_n11304_));
  assign new_n25204_ = ~new_n25205_ & (~new_n13804_ | ((new_n25209_ | new_n15165_) & (~new_n23195_ | ~new_n19148_ | ~new_n15165_)));
  assign new_n25205_ = ~new_n13804_ & new_n25206_ & (new_n25208_ ? ~new_n10645_ : ~new_n25077_);
  assign new_n25206_ = ~new_n10906_ & (~new_n10908_ | ~new_n25207_);
  assign new_n25207_ = new_n10878_ & new_n10899_;
  assign new_n25208_ = new_n7771_ & new_n24550_;
  assign new_n25209_ = (new_n23880_ & ~new_n17896_ & new_n6766_) | (new_n19085_ & new_n25210_ & (new_n17896_ | ~new_n6766_));
  assign new_n25210_ = new_n19060_ & new_n19083_;
  assign new_n25211_ = new_n25212_ & ((~new_n9759_ & new_n25215_) | new_n21964_ | ~new_n25031_);
  assign new_n25212_ = ~new_n25029_ & (~new_n21964_ | ((new_n16230_ | ~new_n24041_ | ~new_n14329_) & (new_n25213_ | new_n14329_)));
  assign new_n25213_ = (~new_n24908_ | new_n12152_) & (new_n25214_ | ~new_n16058_ | ~new_n12152_);
  assign new_n25214_ = ~new_n16030_ & ~new_n16054_;
  assign new_n25215_ = \all_features[855]  | (~new_n25220_ & new_n25221_ & \all_features[854]  & new_n25218_);
  assign new_n25218_ = \all_features[854]  & \all_features[849]  & new_n25219_ & \all_features[848] ;
  assign new_n25219_ = \all_features[853]  & \all_features[852]  & \all_features[850]  & \all_features[851] ;
  assign new_n25220_ = ~\all_features[853]  & (~\all_features[851]  | ~\all_features[852]  | ~\all_features[850]  | (~\all_features[849]  & ~\all_features[848] ));
  assign new_n25221_ = \all_features[853]  & \all_features[854]  & (\all_features[852]  | (\all_features[850]  & \all_features[851]  & \all_features[849] ));
  assign new_n25222_ = new_n25223_ ? (~new_n25238_ ^ new_n25284_) : (new_n25238_ ^ new_n25284_);
  assign new_n25223_ = new_n25224_ ? (new_n25225_ ^ new_n25234_) : (~new_n25225_ ^ new_n25234_);
  assign new_n25224_ = ~new_n24945_ & new_n24959_;
  assign new_n25225_ = new_n25226_ & (new_n12373_ | ~new_n25228_ | (new_n18892_ ? ~new_n8355_ : ~new_n12802_));
  assign new_n25226_ = new_n25230_ & (~new_n25227_ | (~new_n23955_ & new_n14163_ & ~new_n25233_) | (new_n7303_ & new_n25233_));
  assign new_n25227_ = new_n25228_ & new_n12373_;
  assign new_n25228_ = ~new_n22558_ & new_n25229_;
  assign new_n25229_ = ~new_n10611_ & ~new_n10634_;
  assign new_n25230_ = new_n25228_ | ((~new_n21526_ | ~new_n25161_ | new_n25231_) & (new_n25232_ | ~new_n12908_ | ~new_n25231_));
  assign new_n25231_ = ~new_n21354_ & new_n17414_;
  assign new_n25232_ = new_n23338_ & new_n6921_;
  assign new_n25233_ = ~new_n15552_ & ~new_n14528_;
  assign new_n25234_ = (~new_n25235_ | new_n25237_) & (new_n8630_ | new_n25208_ | new_n8923_ | ~new_n25237_);
  assign new_n25235_ = new_n25236_ & (new_n19581_ | (new_n19553_ & new_n19577_));
  assign new_n25236_ = new_n19584_ & new_n22778_ & ~new_n16029_ & ~new_n16058_;
  assign new_n25237_ = new_n9207_ & (new_n9204_ | new_n13402_);
  assign new_n25238_ = ~new_n25239_ & new_n25281_;
  assign new_n25239_ = new_n25240_ & (new_n22548_ | new_n25280_ | ~new_n25279_);
  assign new_n25240_ = (new_n25279_ | ~new_n25276_ | new_n22548_) & (~new_n22548_ | (new_n25277_ ? ~new_n25241_ : new_n25275_));
  assign new_n25241_ = new_n25242_ ? ~new_n24755_ : ~new_n12908_;
  assign new_n25242_ = ~new_n25243_ & new_n25271_;
  assign new_n25243_ = ~new_n25270_ & (new_n25263_ | new_n25266_ | new_n25268_ | new_n25269_ | new_n25244_);
  assign new_n25244_ = ~new_n25257_ & ~new_n25262_ & ((~new_n25245_ & new_n25254_) | new_n25261_ | new_n25259_);
  assign new_n25245_ = new_n25246_ & (new_n25252_ | ~\all_features[749]  | ~\all_features[750]  | ~\all_features[751] );
  assign new_n25246_ = \all_features[751]  & \all_features[750]  & ~new_n25247_ & new_n25250_;
  assign new_n25247_ = new_n25248_ & ~\all_features[749]  & ~new_n25249_ & ~\all_features[748] ;
  assign new_n25248_ = ~\all_features[746]  & ~\all_features[747] ;
  assign new_n25249_ = \all_features[744]  & \all_features[745] ;
  assign new_n25250_ = \all_features[751]  & (\all_features[750]  | (new_n25251_ & (\all_features[746]  | \all_features[747]  | \all_features[745] )));
  assign new_n25251_ = \all_features[748]  & \all_features[749] ;
  assign new_n25252_ = ~\all_features[747]  & ~\all_features[748]  & (~\all_features[746]  | new_n25253_);
  assign new_n25253_ = ~\all_features[744]  & ~\all_features[745] ;
  assign new_n25254_ = new_n25255_ & new_n25256_;
  assign new_n25255_ = \all_features[751]  & (\all_features[750]  | (\all_features[749]  & (\all_features[748]  | ~new_n25253_ | ~new_n25248_)));
  assign new_n25256_ = \all_features[751]  & (\all_features[749]  | \all_features[750]  | \all_features[748] );
  assign new_n25257_ = ~\all_features[751]  & (~\all_features[750]  | (~\all_features[749]  & (new_n25253_ | ~new_n25258_ | ~\all_features[748] )));
  assign new_n25258_ = \all_features[746]  & \all_features[747] ;
  assign new_n25259_ = ~new_n25260_ & ~\all_features[751] ;
  assign new_n25260_ = \all_features[749]  & \all_features[750]  & (\all_features[748]  | (\all_features[746]  & \all_features[747]  & \all_features[745] ));
  assign new_n25261_ = ~\all_features[751]  & (~\all_features[750]  | ~new_n25249_ | ~new_n25251_ | ~new_n25258_);
  assign new_n25262_ = ~\all_features[751]  & (~\all_features[750]  | (~\all_features[748]  & ~\all_features[749]  & ~new_n25258_));
  assign new_n25263_ = ~new_n25262_ & (new_n25257_ | (~new_n25259_ & (new_n25261_ | new_n25264_)));
  assign new_n25264_ = new_n25256_ & (~new_n25255_ | (~new_n25265_ & new_n25250_));
  assign new_n25265_ = ~\all_features[749]  & \all_features[750]  & \all_features[751]  & (\all_features[748]  ? new_n25248_ : (new_n25249_ | ~new_n25248_));
  assign new_n25266_ = new_n25267_ & (~\all_features[749]  | (~\all_features[748]  & (~\all_features[747]  | (~\all_features[746]  & ~\all_features[745] ))));
  assign new_n25267_ = ~\all_features[750]  & ~\all_features[751] ;
  assign new_n25268_ = new_n25267_ & (~\all_features[747]  | ~new_n25251_ | (~\all_features[746]  & ~new_n25249_));
  assign new_n25269_ = ~\all_features[749]  & new_n25267_ & ((~\all_features[746]  & new_n25253_) | ~\all_features[748]  | ~\all_features[747] );
  assign new_n25270_ = ~\all_features[751]  & ~\all_features[750]  & ~\all_features[749]  & ~\all_features[747]  & ~\all_features[748] ;
  assign new_n25271_ = new_n25266_ | ~new_n25273_ | ((new_n25259_ | ~new_n25274_) & (new_n25272_ | new_n25268_));
  assign new_n25272_ = ~new_n25257_ & ~new_n25259_ & ~new_n25261_ & ~new_n25262_ & (~new_n25254_ | ~new_n25246_);
  assign new_n25273_ = ~new_n25269_ & ~new_n25270_;
  assign new_n25274_ = ~new_n25268_ & ~new_n25262_ & ~new_n25257_ & ~new_n25261_;
  assign new_n25275_ = new_n20262_ ? new_n19736_ : ~new_n21851_;
  assign new_n25276_ = new_n16313_ ? new_n22939_ : ~new_n21163_;
  assign new_n25277_ = ~new_n14786_ & (~new_n25278_ | new_n18081_);
  assign new_n25278_ = ~new_n14787_ & new_n14810_;
  assign new_n25279_ = new_n19457_ & (new_n19463_ | new_n19435_);
  assign new_n25280_ = (new_n7558_ | (~new_n23032_ & (new_n23593_ | ~new_n23003_))) & (~new_n13433_ | ~new_n21527_ | new_n23032_ | (~new_n23593_ & new_n23003_));
  assign new_n25281_ = ~new_n25283_ & ~new_n25282_ & (new_n22548_ | (new_n25276_ & ~new_n25279_) | (~new_n25280_ & new_n25279_));
  assign new_n25282_ = new_n24755_ & new_n25242_ & new_n22548_ & new_n25277_;
  assign new_n25283_ = ~new_n25277_ & new_n22548_ & (new_n20262_ ? new_n19736_ : ~new_n21851_);
  assign new_n25284_ = new_n25285_ & ((~new_n25290_ & new_n25321_) | new_n25320_ | ~new_n25291_);
  assign new_n25285_ = ~new_n25288_ | (new_n25286_ ? ~new_n25287_ : (new_n24033_ ? ~new_n23169_ : new_n25289_));
  assign new_n25286_ = new_n6498_ & new_n14159_;
  assign new_n25287_ = new_n15329_ ? ~new_n21527_ : ~new_n21535_;
  assign new_n25288_ = ~new_n7991_ & (~new_n7988_ | new_n14848_);
  assign new_n25289_ = ~new_n18985_ & (~new_n20447_ | ~new_n18962_);
  assign new_n25290_ = ~new_n25288_ | (new_n25286_ ? new_n25287_ : (new_n24033_ ? new_n23169_ : ~new_n25289_));
  assign new_n25291_ = ~new_n25288_ & new_n25292_;
  assign new_n25292_ = new_n25319_ | (~new_n25309_ & new_n25293_);
  assign new_n25293_ = new_n25309_ & (new_n25316_ | (~new_n25315_ & new_n25294_ & (new_n25303_ | new_n25313_)));
  assign new_n25294_ = ~new_n25303_ & ~new_n25305_ & (~new_n25308_ | ~new_n25307_ | new_n25295_);
  assign new_n25295_ = new_n25296_ & ~new_n25301_ & new_n25298_;
  assign new_n25296_ = \all_features[1551]  & (\all_features[1550]  | (new_n25297_ & (\all_features[1546]  | \all_features[1547]  | \all_features[1545] )));
  assign new_n25297_ = \all_features[1548]  & \all_features[1549] ;
  assign new_n25298_ = new_n25300_ & (\all_features[1548]  | \all_features[1549]  | ~new_n25299_ | (\all_features[1545]  & \all_features[1544] ));
  assign new_n25299_ = ~\all_features[1546]  & ~\all_features[1547] ;
  assign new_n25300_ = \all_features[1550]  & \all_features[1551] ;
  assign new_n25301_ = new_n25300_ & \all_features[1549]  & ((~new_n25302_ & \all_features[1546] ) | \all_features[1548]  | \all_features[1547] );
  assign new_n25302_ = ~\all_features[1544]  & ~\all_features[1545] ;
  assign new_n25303_ = ~new_n25304_ & ~\all_features[1551] ;
  assign new_n25304_ = \all_features[1549]  & \all_features[1550]  & (\all_features[1548]  | (\all_features[1546]  & \all_features[1547]  & \all_features[1545] ));
  assign new_n25305_ = ~\all_features[1551]  & (~new_n25297_ | ~\all_features[1544]  | ~\all_features[1545]  | ~\all_features[1550]  | ~new_n25306_);
  assign new_n25306_ = \all_features[1546]  & \all_features[1547] ;
  assign new_n25307_ = \all_features[1551]  & (\all_features[1550]  | (\all_features[1549]  & (\all_features[1548]  | ~new_n25299_ | ~new_n25302_)));
  assign new_n25308_ = \all_features[1551]  & (\all_features[1549]  | \all_features[1550]  | \all_features[1548] );
  assign new_n25309_ = \all_features[1550]  | \all_features[1551]  | (~new_n25312_ & new_n25311_ & \all_features[1549] );
  assign new_n25311_ = new_n25297_ & \all_features[1547]  & (\all_features[1546]  | (\all_features[1544]  & \all_features[1545] ));
  assign new_n25312_ = ~\all_features[1548]  & (~\all_features[1547]  | (~\all_features[1546]  & ~\all_features[1545] ));
  assign new_n25313_ = ~new_n25305_ & (~new_n25308_ | (new_n25307_ & (~new_n25296_ | (~new_n25314_ & new_n25298_))));
  assign new_n25314_ = new_n25300_ & (\all_features[1549]  | (~new_n25299_ & \all_features[1548] ));
  assign new_n25315_ = ~\all_features[1551]  & (~\all_features[1550]  | (~\all_features[1549]  & (new_n25302_ | ~\all_features[1548]  | ~new_n25306_)));
  assign new_n25316_ = ~\all_features[1551]  & (~\all_features[1550]  | (~\all_features[1548]  & ~\all_features[1549]  & ~new_n25306_));
  assign new_n25319_ = ~\all_features[1551]  & ~\all_features[1550]  & ~\all_features[1549]  & ~\all_features[1547]  & ~\all_features[1548] ;
  assign new_n25320_ = ~new_n24981_ & new_n22545_;
  assign new_n25321_ = new_n11169_ & ~new_n7994_ & new_n24981_;
  assign new_n25322_ = ~new_n25323_ & new_n25329_;
  assign new_n25323_ = new_n25324_ & (~new_n25328_ | (~new_n15668_ & new_n16101_) | (~new_n21106_ & ~new_n16101_));
  assign new_n25324_ = (~new_n11272_ | new_n25325_ | new_n22048_) & (new_n21695_ | ~new_n25326_ | ~new_n25327_ | ~new_n22048_);
  assign new_n25325_ = ~new_n12442_ & new_n18099_;
  assign new_n25326_ = new_n13055_ & ~new_n23070_ & new_n10438_;
  assign new_n25327_ = ~new_n9579_ & (~new_n9581_ | new_n12372_);
  assign new_n25328_ = ~new_n25326_ & new_n22048_;
  assign new_n25329_ = ~new_n25330_ & new_n25331_ & (new_n22048_ | (~new_n25325_ & new_n11272_));
  assign new_n25330_ = new_n25328_ & (new_n16101_ ? ~new_n15668_ : ~new_n21106_);
  assign new_n25331_ = ~new_n25326_ | ~new_n22048_ | (new_n25327_ ? ~new_n21695_ : new_n25332_);
  assign new_n25332_ = ~new_n9749_ & (~new_n9755_ | ~new_n9727_);
  assign new_n25333_ = ~new_n25350_ & new_n25334_;
  assign new_n25334_ = ~new_n25335_ & new_n25344_ & (new_n22048_ | (new_n25342_ & ~new_n25348_) | (~new_n25347_ & new_n25348_));
  assign new_n25335_ = new_n19059_ & new_n25336_ & new_n14336_ & (~new_n25338_ | ~new_n19085_);
  assign new_n25336_ = ~new_n25337_ & new_n22048_;
  assign new_n25337_ = new_n21077_ & ~new_n21106_ & ~new_n21108_;
  assign new_n25338_ = ~new_n25339_ & (\all_features[4107]  | \all_features[4108]  | \all_features[4109]  | \all_features[4110]  | \all_features[4111] );
  assign new_n25339_ = ~new_n19078_ & (new_n19082_ | (~new_n19081_ & (new_n19076_ | (~new_n19062_ & ~new_n25340_))));
  assign new_n25340_ = ~new_n19074_ & (new_n19073_ | (new_n19072_ & (~new_n19071_ | (~new_n25341_ & new_n19066_))));
  assign new_n25341_ = ~\all_features[4109]  & \all_features[4110]  & \all_features[4111]  & (\all_features[4108]  ? new_n19069_ : (new_n19070_ | ~new_n19069_));
  assign new_n25342_ = new_n18590_ ? new_n25343_ : ~new_n23879_;
  assign new_n25343_ = new_n11673_ & new_n13204_;
  assign new_n25344_ = ~new_n22048_ | ((new_n25345_ | ~new_n25337_) & (new_n14336_ | ~new_n25346_ | new_n25337_));
  assign new_n25345_ = new_n24975_ ? new_n18323_ : ~new_n25271_;
  assign new_n25346_ = ~new_n14810_ & (~new_n18086_ | ~new_n14787_);
  assign new_n25347_ = ~new_n21278_ & ~new_n25018_ & ~new_n21274_ & ~new_n15674_ & ~new_n21252_;
  assign new_n25348_ = ~new_n25349_ & new_n23124_;
  assign new_n25349_ = new_n6771_ & new_n6795_;
  assign new_n25350_ = new_n25351_ & (new_n14336_ | new_n25346_ | ~new_n25336_);
  assign new_n25351_ = new_n22048_ | (new_n25348_ ? ~new_n25352_ : (new_n18590_ ? ~new_n25343_ : new_n23879_));
  assign new_n25352_ = ~new_n13196_ & new_n15674_ & (~new_n13170_ | new_n13977_);
  assign new_n25353_ = new_n25364_ & new_n25354_ & (~new_n25368_ | (~new_n25369_ & ~new_n25371_));
  assign new_n25354_ = (new_n25363_ | ~new_n25360_) & (new_n15990_ | ~new_n25355_);
  assign new_n25355_ = new_n25358_ & ~new_n17214_ & ~new_n25356_;
  assign new_n25356_ = new_n15078_ & new_n25357_;
  assign new_n25357_ = ~new_n15050_ & ~new_n15074_;
  assign new_n25358_ = ~new_n23736_ & new_n25359_;
  assign new_n25359_ = new_n23766_ & new_n23769_;
  assign new_n25360_ = new_n17214_ & ~new_n25356_ & ~new_n25361_;
  assign new_n25361_ = ~new_n14125_ & new_n25362_;
  assign new_n25362_ = ~new_n14154_ & ~new_n14156_;
  assign new_n25363_ = new_n14607_ & new_n14609_;
  assign new_n25364_ = (new_n25365_ | new_n25356_) & (~new_n25367_ | ~new_n19500_ | ~new_n25356_);
  assign new_n25365_ = (new_n25358_ | new_n17214_) & (~new_n25361_ | ~new_n25366_ | ~new_n17214_);
  assign new_n25366_ = new_n20159_ & ~new_n17817_ & ~new_n17840_;
  assign new_n25367_ = new_n15550_ ? new_n21076_ : new_n25327_;
  assign new_n25368_ = ~new_n19500_ & new_n25356_;
  assign new_n25369_ = new_n25370_ & (new_n10127_ | (new_n10100_ & new_n10125_ & new_n18583_));
  assign new_n25370_ = new_n19432_ & (~new_n16482_ | ~new_n19427_);
  assign new_n25371_ = ~new_n24163_ & ~new_n25370_;
  assign new_n25372_ = new_n25373_ & (~new_n25398_ | (new_n25395_ & new_n25400_));
  assign new_n25373_ = ~new_n25381_ & new_n25374_ & (~new_n25389_ | ~new_n25387_);
  assign new_n25374_ = ~new_n25375_ & (~new_n25380_ | (new_n19342_ & new_n25062_) | (new_n23833_ & ~new_n25062_));
  assign new_n25375_ = new_n25376_ & (new_n25378_ ? ~new_n12490_ : new_n18153_);
  assign new_n25376_ = ~new_n25377_ & new_n22042_;
  assign new_n25377_ = new_n7407_ & (new_n7405_ | ~new_n18176_);
  assign new_n25378_ = new_n25379_ & new_n10677_;
  assign new_n25379_ = new_n10670_ & new_n10679_;
  assign new_n25380_ = ~new_n10737_ & ~new_n22042_;
  assign new_n25381_ = new_n25382_ & (new_n25383_ ? ~new_n25384_ : ~new_n25385_);
  assign new_n25382_ = ~new_n22042_ & new_n10737_;
  assign new_n25383_ = new_n7991_ & (new_n7988_ | ~new_n14848_);
  assign new_n25384_ = ~new_n8507_ & new_n8535_;
  assign new_n25385_ = ~new_n23200_ & new_n25386_;
  assign new_n25386_ = ~new_n23239_ & ~new_n23222_;
  assign new_n25387_ = ~new_n24535_ & new_n25388_;
  assign new_n25388_ = new_n22042_ & new_n25377_;
  assign new_n25389_ = new_n13799_ & (~new_n25390_ | (~new_n25391_ & ~new_n13792_));
  assign new_n25390_ = new_n13775_ & (\all_features[1083]  | \all_features[1084]  | \all_features[1085]  | \all_features[1086]  | \all_features[1087] );
  assign new_n25391_ = ~new_n13795_ & (new_n13796_ | (~new_n13797_ & (new_n13798_ | (~new_n13789_ & ~new_n25392_))));
  assign new_n25392_ = ~new_n13787_ & (~\all_features[1087]  | new_n25393_ | (~\all_features[1084]  & ~\all_features[1085]  & ~\all_features[1086] ));
  assign new_n25393_ = \all_features[1087]  & ((~new_n25394_ & ~\all_features[1085]  & \all_features[1086] ) | (~new_n13783_ & (\all_features[1086]  | (~new_n13778_ & \all_features[1085] ))));
  assign new_n25394_ = (\all_features[1084]  & (\all_features[1082]  | \all_features[1083] )) | (~new_n13786_ & ~\all_features[1082]  & ~\all_features[1083]  & ~\all_features[1084] );
  assign new_n25395_ = new_n25396_ & (~new_n25382_ | (~new_n25384_ & new_n25383_) | (~new_n25385_ & ~new_n25383_));
  assign new_n25396_ = (~new_n25397_ | new_n8267_) & (~new_n25376_ | ~new_n25378_ | ~new_n12490_);
  assign new_n25397_ = new_n25388_ & new_n24535_;
  assign new_n25398_ = new_n25399_ & (~new_n8267_ | ~new_n25397_);
  assign new_n25399_ = (new_n18153_ | new_n25378_ | ~new_n25376_) & (~new_n25380_ | ~new_n19342_ | ~new_n25062_);
  assign new_n25400_ = ~new_n25389_ & new_n25387_;
  assign new_n25401_ = ~new_n25402_ & new_n25416_;
  assign new_n25402_ = new_n25403_ & (~new_n25413_ | ~new_n15282_ | ~new_n23515_);
  assign new_n25403_ = (new_n25412_ | ~new_n25410_) & (new_n24755_ | ~new_n25404_);
  assign new_n25404_ = new_n25405_ & new_n25408_;
  assign new_n25405_ = ~new_n20786_ & new_n25406_;
  assign new_n25406_ = ~new_n16158_ & new_n25407_;
  assign new_n25407_ = ~new_n16188_ & ~new_n16190_;
  assign new_n25408_ = ~new_n18288_ & (~new_n18285_ | new_n25409_);
  assign new_n25409_ = ~new_n24165_ & ~new_n18260_;
  assign new_n25410_ = ~new_n10701_ & new_n25411_;
  assign new_n25411_ = ~new_n20786_ & ~new_n25406_;
  assign new_n25412_ = ~new_n21526_ & new_n16906_;
  assign new_n25413_ = new_n20786_ & new_n25414_;
  assign new_n25414_ = new_n8161_ & (new_n8159_ | new_n25415_);
  assign new_n25415_ = new_n8134_ & new_n24566_;
  assign new_n25416_ = new_n25417_ & new_n25419_ & (~new_n25421_ | ~new_n7161_) & (~new_n25420_ | new_n25422_);
  assign new_n25417_ = (~new_n24755_ | ~new_n25404_) & (~new_n25418_ | (new_n20895_ ? new_n18578_ : ~new_n24759_));
  assign new_n25418_ = ~new_n25414_ & new_n20786_;
  assign new_n25419_ = (~new_n25412_ | ~new_n25410_) & (~new_n25413_ | (new_n23515_ ? new_n15282_ : new_n25231_));
  assign new_n25420_ = ~new_n25408_ & new_n25405_;
  assign new_n25421_ = new_n25411_ & new_n10701_;
  assign new_n25422_ = new_n17414_ & (new_n17392_ | (new_n19639_ & new_n19644_));
  assign \o[43]  = new_n25424_ ? (new_n25425_ ^ new_n25475_) : (~new_n25425_ ^ new_n25475_);
  assign new_n25424_ = (new_n25372_ & new_n25401_) | (new_n24701_ & (new_n25372_ | new_n25401_));
  assign new_n25425_ = new_n25426_ ? (~new_n25473_ ^ new_n25474_) : (new_n25473_ ^ new_n25474_);
  assign new_n25426_ = new_n25427_ ? (new_n25465_ ^ new_n25466_) : (~new_n25465_ ^ new_n25466_);
  assign new_n25427_ = new_n25428_ ? (new_n25451_ ^ new_n25452_) : (~new_n25451_ ^ new_n25452_);
  assign new_n25428_ = new_n25429_ ? (new_n25441_ ^ new_n25442_) : (~new_n25441_ ^ new_n25442_);
  assign new_n25429_ = new_n25430_ ? (~new_n25431_ ^ new_n25437_) : (new_n25431_ ^ new_n25437_);
  assign new_n25430_ = ~new_n24707_ & ~new_n24786_;
  assign new_n25431_ = new_n25432_ ? (new_n25433_ ^ new_n25436_) : (~new_n25433_ ^ new_n25436_);
  assign new_n25432_ = new_n25334_ & new_n25350_;
  assign new_n25433_ = new_n25402_ & ~new_n25434_ & new_n25416_;
  assign new_n25434_ = new_n25435_ & (new_n7161_ | ~new_n25421_);
  assign new_n25435_ = (~new_n25422_ | ~new_n25420_) & (~new_n25418_ | (new_n20895_ ? ~new_n18578_ : new_n24759_));
  assign new_n25436_ = new_n24902_ & new_n24914_;
  assign new_n25437_ = new_n25438_ ? (new_n25439_ ^ new_n25440_) : (~new_n25439_ ^ new_n25440_);
  assign new_n25438_ = new_n25373_ & new_n25398_;
  assign new_n25439_ = new_n24847_ & new_n24788_;
  assign new_n25440_ = new_n24709_ & new_n24756_;
  assign new_n25441_ = (~new_n24849_ & new_n24944_) | (~new_n24706_ & (~new_n24849_ | new_n24944_));
  assign new_n25442_ = new_n25443_ ? (~new_n25444_ ^ new_n25445_) : (new_n25444_ ^ new_n25445_);
  assign new_n25443_ = (new_n24901_ & new_n24918_) | (new_n24850_ & (new_n24901_ | new_n24918_));
  assign new_n25444_ = (new_n24978_ & new_n24982_) | (new_n24963_ & (new_n24978_ | new_n24982_));
  assign new_n25445_ = new_n25446_ ? (new_n25447_ ^ new_n25450_) : (~new_n25447_ ^ new_n25450_);
  assign new_n25446_ = new_n24899_ & new_n24852_;
  assign new_n25447_ = new_n25353_ & new_n25448_;
  assign new_n25448_ = new_n25449_ & (new_n25367_ | ~new_n25356_ | ~new_n19500_) & (~new_n25360_ | ~new_n25363_);
  assign new_n25449_ = (~new_n15990_ | ~new_n25355_) & (new_n25371_ | new_n25369_ | ~new_n25368_);
  assign new_n25450_ = ~new_n24943_ & new_n24919_;
  assign new_n25451_ = (~new_n24961_ & new_n24997_) | (~new_n24705_ & (~new_n24961_ | new_n24997_));
  assign new_n25452_ = new_n25453_ ? (~new_n25463_ ^ new_n25464_) : (new_n25463_ ^ new_n25464_);
  assign new_n25453_ = new_n25454_ ? (new_n25458_ ^ new_n25459_) : (~new_n25458_ ^ new_n25459_);
  assign new_n25454_ = new_n25455_ ? (new_n25456_ ^ new_n25457_) : (~new_n25456_ ^ new_n25457_);
  assign new_n25455_ = new_n25323_ & new_n25329_;
  assign new_n25456_ = new_n24964_ & new_n24976_;
  assign new_n25457_ = new_n25290_ & new_n25285_ & (~new_n25291_ | (~new_n25320_ & new_n25321_));
  assign new_n25458_ = (new_n25027_ & new_n25038_) | (new_n25007_ & (new_n25027_ | new_n25038_));
  assign new_n25459_ = new_n25460_ ? (new_n25461_ ^ new_n25462_) : (~new_n25461_ ^ new_n25462_);
  assign new_n25460_ = new_n25239_ & new_n25281_;
  assign new_n25461_ = new_n25028_ & new_n25036_;
  assign new_n25462_ = ~new_n24987_ & new_n24983_;
  assign new_n25463_ = (~new_n25072_ & new_n25143_) | (~new_n25006_ & (~new_n25072_ | new_n25143_));
  assign new_n25464_ = (new_n24944_ & new_n24988_) | (~new_n24962_ & (new_n24944_ | new_n24988_));
  assign new_n25465_ = (~new_n25004_ & new_n25211_) | (~new_n24704_ & (~new_n25004_ | new_n25211_));
  assign new_n25466_ = new_n25467_ ? (~new_n25471_ ^ new_n25472_) : (new_n25471_ ^ new_n25472_);
  assign new_n25467_ = new_n25468_ ? (new_n25469_ ^ new_n25470_) : (~new_n25469_ ^ new_n25470_);
  assign new_n25468_ = new_n25150_ & new_n25200_;
  assign new_n25469_ = new_n25008_ & new_n25025_;
  assign new_n25470_ = (new_n25106_ & new_n25140_) | (new_n25073_ & (new_n25106_ | new_n25140_));
  assign new_n25471_ = (new_n25149_ & new_n25202_) | (~new_n25005_ & (new_n25149_ | new_n25202_));
  assign new_n25472_ = (new_n25225_ & new_n25234_) | (new_n25224_ & (new_n25225_ | new_n25234_));
  assign new_n25473_ = (~new_n25222_ & new_n25322_) | (~new_n24703_ & (~new_n25222_ | new_n25322_));
  assign new_n25474_ = (new_n25238_ & new_n25284_) | (~new_n25223_ & (new_n25238_ | new_n25284_));
  assign new_n25475_ = (new_n25333_ & new_n25353_) | (~new_n24702_ & (new_n25333_ | new_n25353_));
  assign \o[44]  = ~new_n25477_ ^ new_n25478_;
  assign new_n25477_ = (~new_n25425_ & new_n25475_) | (new_n25424_ & (~new_n25425_ | new_n25475_));
  assign new_n25478_ = new_n25479_ ^ new_n25480_;
  assign new_n25479_ = (new_n25473_ & new_n25474_) | (~new_n25426_ & (new_n25473_ | new_n25474_));
  assign new_n25480_ = new_n25481_ ? (~new_n25482_ ^ new_n25505_) : (new_n25482_ ^ new_n25505_);
  assign new_n25481_ = (~new_n25466_ & new_n25465_) | (~new_n25427_ & (~new_n25466_ | new_n25465_));
  assign new_n25482_ = new_n25483_ ? (new_n25484_ ^ new_n25501_) : (~new_n25484_ ^ new_n25501_);
  assign new_n25483_ = (~new_n25452_ & new_n25451_) | (~new_n25428_ & (~new_n25452_ | new_n25451_));
  assign new_n25484_ = new_n25485_ ? (new_n25486_ ^ new_n25497_) : (~new_n25486_ ^ new_n25497_);
  assign new_n25485_ = (~new_n25442_ & new_n25441_) | (~new_n25429_ & (~new_n25442_ | new_n25441_));
  assign new_n25486_ = new_n25487_ ? (new_n25488_ ^ new_n25494_) : (~new_n25488_ ^ new_n25494_);
  assign new_n25487_ = (~new_n25431_ & ~new_n25437_) | (~new_n25430_ & (~new_n25431_ | ~new_n25437_));
  assign new_n25488_ = new_n25489_ ? (~new_n25492_ ^ new_n25493_) : (new_n25492_ ^ new_n25493_);
  assign new_n25489_ = new_n25490_ ^ new_n25491_;
  assign new_n25490_ = new_n25438_ & ~new_n25400_ & new_n25395_;
  assign new_n25491_ = new_n25439_ & new_n24807_;
  assign new_n25492_ = (new_n25439_ & new_n25440_) | (new_n25438_ & (new_n25439_ | new_n25440_));
  assign new_n25493_ = new_n25434_ & new_n25402_ & new_n25416_;
  assign new_n25494_ = ~new_n25495_ ^ new_n25496_;
  assign new_n25495_ = (new_n25433_ & new_n25436_) | (new_n25432_ & (new_n25433_ | new_n25436_));
  assign new_n25496_ = (new_n25447_ & new_n25450_) | (new_n25446_ & (new_n25447_ | new_n25450_));
  assign new_n25497_ = new_n25498_ ? (new_n25499_ ^ new_n25500_) : (~new_n25499_ ^ new_n25500_);
  assign new_n25498_ = (~new_n25445_ & new_n25444_) | (new_n25443_ & (~new_n25445_ | new_n25444_));
  assign new_n25499_ = (~new_n25459_ & new_n25458_) | (~new_n25454_ & (~new_n25459_ | new_n25458_));
  assign new_n25500_ = (new_n25456_ & new_n25457_) | (new_n25455_ & (new_n25456_ | new_n25457_));
  assign new_n25501_ = new_n25502_ ? (new_n25503_ ^ new_n25504_) : (~new_n25503_ ^ new_n25504_);
  assign new_n25502_ = (new_n25463_ & new_n25464_) | (~new_n25453_ & (new_n25463_ | new_n25464_));
  assign new_n25503_ = (new_n25469_ & new_n25470_) | (new_n25468_ & (new_n25469_ | new_n25470_));
  assign new_n25504_ = (new_n25461_ & new_n25462_) | (new_n25460_ & (new_n25461_ | new_n25462_));
  assign new_n25505_ = (new_n25471_ & new_n25472_) | (~new_n25467_ & (new_n25471_ | new_n25472_));
  assign \o[45]  = ((new_n25507_ | new_n25508_) & (new_n25509_ ^ new_n25510_)) | (~new_n25507_ & ~new_n25508_ & (~new_n25509_ ^ new_n25510_));
  assign new_n25507_ = ~new_n25478_ & new_n25477_;
  assign new_n25508_ = ~new_n25480_ & new_n25479_;
  assign new_n25509_ = (~new_n25482_ & new_n25505_) | (new_n25481_ & (~new_n25482_ | new_n25505_));
  assign new_n25510_ = new_n25511_ ? (~new_n25512_ ^ new_n25521_) : (new_n25512_ ^ new_n25521_);
  assign new_n25511_ = (~new_n25484_ & ~new_n25501_) | (new_n25483_ & (~new_n25484_ | ~new_n25501_));
  assign new_n25512_ = new_n25513_ ? (~new_n25514_ ^ new_n25520_) : (new_n25514_ ^ new_n25520_);
  assign new_n25513_ = (~new_n25486_ & ~new_n25497_) | (new_n25485_ & (~new_n25486_ | ~new_n25497_));
  assign new_n25514_ = new_n25515_ ? (~new_n25516_ ^ new_n25519_) : (new_n25516_ ^ new_n25519_);
  assign new_n25515_ = (~new_n25488_ & ~new_n25494_) | (new_n25487_ & (~new_n25488_ | ~new_n25494_));
  assign new_n25516_ = new_n25517_ ^ new_n25518_;
  assign new_n25517_ = (new_n25492_ & new_n25493_) | (~new_n25489_ & (new_n25492_ | new_n25493_));
  assign new_n25518_ = ~new_n25490_ & ~new_n25491_;
  assign new_n25519_ = new_n25495_ & new_n25496_;
  assign new_n25520_ = (new_n25499_ & new_n25500_) | (new_n25498_ & (new_n25499_ | new_n25500_));
  assign new_n25521_ = (new_n25503_ & new_n25504_) | (new_n25502_ & (new_n25503_ | new_n25504_));
  assign \o[46]  = ~new_n25523_ ^ new_n25524_;
  assign new_n25523_ = (new_n25509_ | (~new_n25510_ & (new_n25508_ | new_n25507_))) & (new_n25508_ | new_n25507_ | ~new_n25510_);
  assign new_n25524_ = new_n25525_ ^ new_n25526_;
  assign new_n25525_ = (~new_n25512_ & new_n25521_) | (new_n25511_ & (~new_n25512_ | new_n25521_));
  assign new_n25526_ = new_n25527_ ^ new_n25528_;
  assign new_n25527_ = (~new_n25514_ & new_n25520_) | (new_n25513_ & (~new_n25514_ | new_n25520_));
  assign new_n25528_ = ~new_n25529_ ^ new_n25530_;
  assign new_n25529_ = (~new_n25516_ & new_n25519_) | (new_n25515_ & (~new_n25516_ | new_n25519_));
  assign new_n25530_ = ~new_n25518_ & new_n25517_;
  assign \o[47]  = ((new_n25532_ | new_n25533_) & (~new_n25534_ ^ new_n25535_)) | (~new_n25532_ & ~new_n25533_ & (new_n25534_ ^ new_n25535_));
  assign new_n25532_ = ~new_n25524_ & new_n25523_;
  assign new_n25533_ = ~new_n25526_ & new_n25525_;
  assign new_n25534_ = ~new_n25528_ & new_n25527_;
  assign new_n25535_ = new_n25529_ & new_n25530_;
  assign \o[48]  = (new_n25535_ | new_n25532_ | new_n25533_) & (new_n25534_ | (new_n25535_ & (new_n25532_ | new_n25533_)));
  assign \o[49]  = new_n25538_ ^ new_n26391_;
  assign new_n25538_ = new_n25539_ ? (new_n26368_ ^ new_n26386_) : (~new_n26368_ ^ new_n26386_);
  assign new_n25539_ = new_n25540_ ? (~new_n26292_ ^ new_n26305_) : (new_n26292_ ^ new_n26305_);
  assign new_n25540_ = new_n25541_ ? (new_n26204_ ^ new_n26291_) : (~new_n26204_ ^ new_n26291_);
  assign new_n25541_ = new_n25542_ ? (new_n26046_ ^ new_n26157_) : (~new_n26046_ ^ new_n26157_);
  assign new_n25542_ = new_n25543_ ? (new_n25926_ ^ new_n26045_) : (~new_n25926_ ^ new_n26045_);
  assign new_n25543_ = new_n25544_ ? (new_n25759_ ^ new_n25910_) : (~new_n25759_ ^ new_n25910_);
  assign new_n25544_ = new_n25545_ ? (new_n25648_ ^ new_n25703_) : (~new_n25648_ ^ new_n25703_);
  assign new_n25545_ = new_n25546_ & (new_n25624_ | ~new_n25623_);
  assign new_n25546_ = new_n25547_ & new_n25612_ & (~new_n25614_ | ~new_n25613_);
  assign new_n25547_ = new_n25550_ & (~new_n25610_ | ~new_n25548_) & (~new_n25609_ | ~new_n25611_);
  assign new_n25548_ = new_n20233_ & ~new_n18578_ & new_n25549_;
  assign new_n25549_ = ~new_n14877_ & new_n11725_;
  assign new_n25550_ = (new_n25578_ | ~new_n25553_) & (~new_n25551_ | ~new_n20235_);
  assign new_n25551_ = new_n25552_ & ~new_n20233_ & new_n14384_;
  assign new_n25552_ = new_n19090_ & new_n15702_;
  assign new_n25553_ = new_n25554_ & ~new_n14384_ & ~new_n20233_;
  assign new_n25554_ = ~new_n25574_ & (new_n25555_ | new_n25576_ | new_n25577_);
  assign new_n25555_ = ~new_n25573_ & new_n25568_ & (~new_n25558_ | ~new_n25562_) & (new_n25556_ | new_n25571_);
  assign new_n25556_ = ~new_n25566_ & ~new_n25557_ & ~new_n25564_;
  assign new_n25557_ = new_n25558_ & (~new_n25562_ | (~new_n25561_ & \all_features[2717]  & \all_features[2718]  & \all_features[2719] ));
  assign new_n25558_ = \all_features[2719]  & (\all_features[2718]  | (\all_features[2717]  & (\all_features[2716]  | ~new_n25560_ | ~new_n25559_)));
  assign new_n25559_ = ~\all_features[2712]  & ~\all_features[2713] ;
  assign new_n25560_ = ~\all_features[2714]  & ~\all_features[2715] ;
  assign new_n25561_ = ~\all_features[2715]  & ~\all_features[2716]  & (~\all_features[2714]  | new_n25559_);
  assign new_n25562_ = \all_features[2718]  & \all_features[2719]  & (\all_features[2716]  | \all_features[2717]  | new_n25563_ | ~new_n25560_);
  assign new_n25563_ = \all_features[2712]  & \all_features[2713] ;
  assign new_n25564_ = ~new_n25565_ & ~\all_features[2719] ;
  assign new_n25565_ = \all_features[2717]  & \all_features[2718]  & (\all_features[2716]  | (\all_features[2714]  & \all_features[2715]  & \all_features[2713] ));
  assign new_n25566_ = ~\all_features[2719]  & (~new_n25567_ | ~\all_features[2716]  | ~\all_features[2717]  | ~\all_features[2718]  | ~new_n25563_);
  assign new_n25567_ = \all_features[2714]  & \all_features[2715] ;
  assign new_n25568_ = ~new_n25572_ & ~new_n25571_ & ~new_n25566_ & ~new_n25564_ & ~new_n25569_;
  assign new_n25569_ = new_n25570_ & (~\all_features[2717]  | (~\all_features[2716]  & (~\all_features[2715]  | (~\all_features[2714]  & ~\all_features[2713] ))));
  assign new_n25570_ = ~\all_features[2718]  & ~\all_features[2719] ;
  assign new_n25571_ = ~\all_features[2719]  & (~\all_features[2718]  | (~\all_features[2716]  & ~\all_features[2717]  & ~new_n25567_));
  assign new_n25572_ = new_n25570_ & (~\all_features[2715]  | ~\all_features[2716]  | ~\all_features[2717]  | (~\all_features[2714]  & ~new_n25563_));
  assign new_n25573_ = ~\all_features[2719]  & (~\all_features[2718]  | (~\all_features[2717]  & (new_n25559_ | ~\all_features[2716]  | ~new_n25567_)));
  assign new_n25574_ = new_n25575_ & ~new_n25577_ & ~new_n25566_ & ~new_n25564_ & ~new_n25569_;
  assign new_n25575_ = ~new_n25572_ & ~new_n25576_ & ~new_n25573_ & ~new_n25571_;
  assign new_n25576_ = ~\all_features[2717]  & new_n25570_ & ((~\all_features[2714]  & new_n25559_) | ~\all_features[2716]  | ~\all_features[2715] );
  assign new_n25577_ = ~\all_features[2719]  & ~\all_features[2718]  & ~\all_features[2717]  & ~\all_features[2715]  & ~\all_features[2716] ;
  assign new_n25578_ = ~new_n25579_ & new_n25601_ & (new_n25608_ | new_n25584_ | new_n25586_ | ~new_n25606_);
  assign new_n25579_ = ~new_n25594_ & (new_n25596_ | (~new_n25598_ & (new_n25599_ | (~new_n25580_ & ~new_n25600_))));
  assign new_n25580_ = ~new_n25584_ & (new_n25586_ | (new_n25593_ & (~new_n25581_ | (~new_n25590_ & new_n25592_))));
  assign new_n25581_ = \all_features[5935]  & (\all_features[5934]  | new_n25582_);
  assign new_n25582_ = \all_features[5933]  & (\all_features[5930]  | \all_features[5931]  | \all_features[5932]  | ~new_n25583_);
  assign new_n25583_ = ~\all_features[5928]  & ~\all_features[5929] ;
  assign new_n25584_ = ~new_n25585_ & ~\all_features[5935] ;
  assign new_n25585_ = \all_features[5933]  & \all_features[5934]  & (\all_features[5932]  | (\all_features[5930]  & \all_features[5931]  & \all_features[5929] ));
  assign new_n25586_ = ~\all_features[5935]  & (~\all_features[5934]  | ~new_n25587_ | ~new_n25588_ | ~new_n25589_);
  assign new_n25587_ = \all_features[5928]  & \all_features[5929] ;
  assign new_n25588_ = \all_features[5932]  & \all_features[5933] ;
  assign new_n25589_ = \all_features[5930]  & \all_features[5931] ;
  assign new_n25590_ = ~\all_features[5933]  & new_n25591_ & ((~\all_features[5932]  & (new_n25587_ | \all_features[5930]  | \all_features[5931] )) | (~\all_features[5930]  & ~\all_features[5931]  & \all_features[5932] ));
  assign new_n25591_ = \all_features[5934]  & \all_features[5935] ;
  assign new_n25592_ = \all_features[5935]  & (\all_features[5934]  | (new_n25588_ & (\all_features[5930]  | \all_features[5931]  | \all_features[5929] )));
  assign new_n25593_ = \all_features[5935]  & (\all_features[5933]  | \all_features[5934]  | \all_features[5932] );
  assign new_n25594_ = new_n25595_ & ((~\all_features[5930]  & new_n25583_) | ~\all_features[5932]  | ~\all_features[5931] );
  assign new_n25595_ = ~\all_features[5935]  & ~\all_features[5933]  & ~\all_features[5934] ;
  assign new_n25596_ = ~\all_features[5935]  & ~new_n25597_ & ~\all_features[5934] ;
  assign new_n25597_ = \all_features[5933]  & (\all_features[5932]  | (\all_features[5931]  & (\all_features[5930]  | \all_features[5929] )));
  assign new_n25598_ = ~\all_features[5934]  & ~\all_features[5935]  & (~\all_features[5931]  | ~new_n25588_ | (~\all_features[5930]  & ~new_n25587_));
  assign new_n25599_ = ~\all_features[5935]  & (~\all_features[5934]  | (~\all_features[5932]  & ~\all_features[5933]  & ~new_n25589_));
  assign new_n25600_ = ~\all_features[5935]  & (~\all_features[5934]  | (~\all_features[5933]  & (new_n25583_ | ~new_n25589_ | ~\all_features[5932] )));
  assign new_n25601_ = ~new_n25596_ & ~new_n25584_ & new_n25607_ & new_n25606_ & (new_n25586_ | new_n25602_);
  assign new_n25602_ = new_n25593_ & ~new_n25603_ & new_n25581_;
  assign new_n25603_ = new_n25592_ & new_n25604_ & (~\all_features[5933]  | ~new_n25591_ | new_n25605_);
  assign new_n25604_ = new_n25591_ & (new_n25587_ | \all_features[5930]  | \all_features[5931]  | \all_features[5932]  | \all_features[5933] );
  assign new_n25605_ = ~\all_features[5931]  & ~\all_features[5932]  & (~\all_features[5930]  | new_n25583_);
  assign new_n25606_ = ~new_n25599_ & ~new_n25600_;
  assign new_n25607_ = ~new_n25594_ & ~new_n25598_ & ~new_n25586_ & (\all_features[5932]  | \all_features[5931]  | ~new_n25595_);
  assign new_n25608_ = new_n25593_ & new_n25592_ & new_n25581_ & new_n25604_;
  assign new_n25609_ = ~new_n25554_ & ~new_n14384_ & ~new_n20233_;
  assign new_n25610_ = ~new_n21189_ & ~new_n17734_;
  assign new_n25611_ = new_n16562_ & (new_n16559_ | new_n16528_);
  assign new_n25612_ = ~new_n20233_ | ((new_n25549_ | new_n18578_) & (new_n12371_ | new_n23550_ | ~new_n18578_));
  assign new_n25613_ = new_n14384_ & ~new_n20233_ & ~new_n25552_;
  assign new_n25614_ = ~new_n25619_ & ~new_n21111_ & ~new_n25615_;
  assign new_n25615_ = ~new_n25616_ & (\all_features[5667]  | \all_features[5668]  | \all_features[5669]  | \all_features[5670]  | \all_features[5671] );
  assign new_n25616_ = ~new_n21113_ & (new_n21116_ | (~new_n21117_ & (new_n21131_ | (~new_n21126_ & ~new_n25617_))));
  assign new_n25617_ = ~new_n21128_ & (new_n21130_ | (new_n21124_ & (~new_n21132_ | (~new_n25618_ & new_n21121_))));
  assign new_n25618_ = ~\all_features[5669]  & \all_features[5670]  & \all_features[5671]  & (\all_features[5668]  ? new_n21123_ : (new_n21119_ | ~new_n21123_));
  assign new_n25619_ = new_n21112_ & (new_n21117_ | new_n21116_ | (~new_n21126_ & ~new_n21131_ & ~new_n25620_));
  assign new_n25620_ = ~new_n21130_ & ~new_n21128_ & (~new_n21124_ | ~new_n21132_ | new_n25621_);
  assign new_n25621_ = new_n21121_ & new_n21122_ & (new_n25622_ | ~\all_features[5669]  | ~\all_features[5670]  | ~\all_features[5671] );
  assign new_n25622_ = ~\all_features[5667]  & ~\all_features[5668]  & (~\all_features[5666]  | new_n21114_);
  assign new_n25623_ = (new_n25610_ | ~new_n25548_) & (~new_n25553_ | ~new_n25578_) & (new_n25614_ | ~new_n25613_);
  assign new_n25624_ = ~new_n25625_ & (new_n20235_ | ~new_n25551_);
  assign new_n25625_ = new_n18578_ & new_n20233_ & (new_n12371_ ? ~new_n25626_ : new_n23550_);
  assign new_n25626_ = ~new_n25627_ & ~new_n25645_ & (new_n25647_ | \all_features[5981]  | \all_features[5982]  | \all_features[5983] );
  assign new_n25627_ = new_n25628_ & (~new_n25643_ | (~new_n25641_ & ~new_n25644_ & ~new_n25638_ & new_n25645_));
  assign new_n25628_ = ~new_n25629_ & ~new_n25632_ & ~new_n25638_ & new_n25640_ & (~new_n25637_ | ~new_n25635_);
  assign new_n25629_ = ~\all_features[5983]  & ~new_n25630_ & ~\all_features[5982] ;
  assign new_n25630_ = \all_features[5979]  & \all_features[5980]  & \all_features[5981]  & (\all_features[5978]  | new_n25631_);
  assign new_n25631_ = \all_features[5976]  & \all_features[5977] ;
  assign new_n25632_ = ~\all_features[5983]  & (~\all_features[5982]  | (~\all_features[5981]  & (new_n25634_ | ~\all_features[5980]  | ~new_n25633_)));
  assign new_n25633_ = \all_features[5978]  & \all_features[5979] ;
  assign new_n25634_ = ~\all_features[5976]  & ~\all_features[5977] ;
  assign new_n25635_ = \all_features[5983]  & (\all_features[5982]  | (\all_features[5981]  & (\all_features[5980]  | ~new_n25636_ | ~new_n25634_)));
  assign new_n25636_ = ~\all_features[5978]  & ~\all_features[5979] ;
  assign new_n25637_ = \all_features[5982]  & \all_features[5983]  & (\all_features[5980]  | \all_features[5981]  | new_n25631_ | ~new_n25636_);
  assign new_n25638_ = ~new_n25639_ & ~\all_features[5983] ;
  assign new_n25639_ = \all_features[5981]  & \all_features[5982]  & (\all_features[5980]  | (\all_features[5978]  & \all_features[5979]  & \all_features[5977] ));
  assign new_n25640_ = \all_features[5983]  | (new_n25631_ & \all_features[5980]  & \all_features[5981]  & \all_features[5982]  & new_n25633_);
  assign new_n25641_ = new_n25635_ & (~new_n25637_ | (~new_n25642_ & \all_features[5981]  & \all_features[5982]  & \all_features[5983] ));
  assign new_n25642_ = ~\all_features[5979]  & ~\all_features[5980]  & (~\all_features[5978]  | new_n25634_);
  assign new_n25643_ = \all_features[5983]  | (\all_features[5982]  & (\all_features[5981]  | (~new_n25634_ & \all_features[5980]  & new_n25633_)));
  assign new_n25644_ = ~\all_features[5983]  & (~new_n25631_ | ~\all_features[5980]  | ~\all_features[5981]  | ~\all_features[5982]  | ~new_n25633_);
  assign new_n25645_ = ~\all_features[5983]  & ~\all_features[5982]  & ~\all_features[5981]  & ~\all_features[5979]  & ~\all_features[5980] ;
  assign new_n25647_ = \all_features[5979]  & \all_features[5980]  & (\all_features[5978]  | ~new_n25634_);
  assign new_n25648_ = ~new_n25649_ & new_n25702_;
  assign new_n25649_ = ~new_n25664_ & new_n25650_ & (new_n23188_ | ~new_n10645_ | new_n25667_);
  assign new_n25650_ = ~new_n25651_ & (new_n10645_ | (~new_n24132_ & new_n25656_ & new_n25662_) | (~new_n25654_ & ~new_n25662_));
  assign new_n25651_ = ~new_n25653_ & new_n25652_;
  assign new_n25652_ = new_n10645_ & new_n23188_;
  assign new_n25653_ = new_n6662_ & (new_n6640_ | ~new_n6665_);
  assign new_n25654_ = ~new_n25655_ & new_n23550_;
  assign new_n25655_ = ~new_n7251_ & (~new_n7253_ | ~new_n7229_);
  assign new_n25656_ = new_n21536_ & new_n25657_;
  assign new_n25657_ = ~new_n22786_ & ~new_n25658_;
  assign new_n25658_ = ~new_n25659_ & (\all_features[4635]  | \all_features[4636]  | \all_features[4637]  | \all_features[4638]  | \all_features[4639] );
  assign new_n25659_ = ~new_n21540_ & (new_n21543_ | (~new_n21544_ & (new_n21553_ | (~new_n21548_ & ~new_n25660_))));
  assign new_n25660_ = ~new_n21550_ & (new_n21552_ | (new_n21558_ & (~new_n21554_ | (~new_n25661_ & new_n21556_))));
  assign new_n25661_ = ~\all_features[4637]  & \all_features[4638]  & \all_features[4639]  & (\all_features[4636]  ? new_n21555_ : (new_n21546_ | ~new_n21555_));
  assign new_n25662_ = new_n25663_ & new_n8132_;
  assign new_n25663_ = new_n8121_ & new_n8129_;
  assign new_n25664_ = new_n25665_ & (new_n25655_ ? new_n25666_ : ~new_n23550_);
  assign new_n25665_ = ~new_n10645_ & ~new_n25662_;
  assign new_n25666_ = ~new_n15332_ & (~new_n20465_ | new_n20473_);
  assign new_n25667_ = new_n7339_ ? new_n25208_ : (new_n25700_ | (new_n25668_ & new_n25690_ & new_n25696_));
  assign new_n25668_ = ~new_n25669_ & ~new_n25689_;
  assign new_n25669_ = ~new_n25687_ & (new_n25684_ | (~new_n25686_ & (new_n25688_ | (~new_n25670_ & ~new_n25673_))));
  assign new_n25670_ = ~\all_features[2063]  & (~\all_features[2062]  | new_n25671_);
  assign new_n25671_ = ~\all_features[2061]  & (new_n25672_ | ~\all_features[2059]  | ~\all_features[2060]  | ~\all_features[2058] );
  assign new_n25672_ = ~\all_features[2056]  & ~\all_features[2057] ;
  assign new_n25673_ = ~new_n25674_ & (new_n25676_ | (new_n25683_ & (~new_n25679_ | (~new_n25682_ & new_n25681_))));
  assign new_n25674_ = ~new_n25675_ & ~\all_features[2063] ;
  assign new_n25675_ = \all_features[2061]  & \all_features[2062]  & (\all_features[2060]  | (\all_features[2058]  & \all_features[2059]  & \all_features[2057] ));
  assign new_n25676_ = ~\all_features[2063]  & (~new_n25678_ | ~\all_features[2058]  | ~\all_features[2059]  | ~\all_features[2062]  | ~new_n25677_);
  assign new_n25677_ = \all_features[2056]  & \all_features[2057] ;
  assign new_n25678_ = \all_features[2060]  & \all_features[2061] ;
  assign new_n25679_ = \all_features[2063]  & (\all_features[2062]  | (\all_features[2061]  & (\all_features[2060]  | ~new_n25680_ | ~new_n25672_)));
  assign new_n25680_ = ~\all_features[2058]  & ~\all_features[2059] ;
  assign new_n25681_ = \all_features[2063]  & (\all_features[2062]  | (new_n25678_ & (\all_features[2058]  | \all_features[2059]  | \all_features[2057] )));
  assign new_n25682_ = ~\all_features[2061]  & \all_features[2062]  & \all_features[2063]  & (\all_features[2060]  ? new_n25680_ : (new_n25677_ | ~new_n25680_));
  assign new_n25683_ = \all_features[2063]  & (\all_features[2061]  | \all_features[2062]  | \all_features[2060] );
  assign new_n25684_ = new_n25685_ & (~\all_features[2061]  | (~\all_features[2060]  & (~\all_features[2059]  | (~\all_features[2058]  & ~\all_features[2057] ))));
  assign new_n25685_ = ~\all_features[2062]  & ~\all_features[2063] ;
  assign new_n25686_ = new_n25685_ & (~\all_features[2059]  | ~new_n25678_ | (~\all_features[2058]  & ~new_n25677_));
  assign new_n25687_ = ~\all_features[2061]  & new_n25685_ & ((~\all_features[2058]  & new_n25672_) | ~\all_features[2060]  | ~\all_features[2059] );
  assign new_n25688_ = ~\all_features[2063]  & (~\all_features[2062]  | (~\all_features[2061]  & ~\all_features[2060]  & (~\all_features[2059]  | ~\all_features[2058] )));
  assign new_n25689_ = ~\all_features[2063]  & ~\all_features[2062]  & ~\all_features[2061]  & ~\all_features[2059]  & ~\all_features[2060] ;
  assign new_n25690_ = new_n25695_ & ~new_n25691_ & new_n25694_;
  assign new_n25691_ = ~new_n25688_ & ~new_n25676_ & ~new_n25674_ & ~new_n25670_ & ~new_n25692_;
  assign new_n25692_ = new_n25683_ & new_n25693_ & new_n25679_ & new_n25681_;
  assign new_n25693_ = \all_features[2062]  & \all_features[2063]  & (\all_features[2060]  | \all_features[2061]  | new_n25677_ | ~new_n25680_);
  assign new_n25694_ = ~new_n25687_ & ~new_n25689_;
  assign new_n25695_ = ~new_n25684_ & ~new_n25686_;
  assign new_n25696_ = new_n25694_ & (~new_n25695_ | (~new_n25670_ & ~new_n25697_ & ~new_n25688_));
  assign new_n25697_ = ~new_n25674_ & ~new_n25676_ & (~new_n25683_ | ~new_n25679_ | new_n25698_);
  assign new_n25698_ = new_n25681_ & new_n25693_ & (new_n25699_ | ~\all_features[2061]  | ~\all_features[2062]  | ~\all_features[2063] );
  assign new_n25699_ = ~\all_features[2059]  & ~\all_features[2060]  & (~\all_features[2058]  | new_n25672_);
  assign new_n25700_ = new_n25701_ & ~new_n25688_ & ~new_n25687_ & ~new_n25670_ & ~new_n25686_;
  assign new_n25701_ = ~new_n25689_ & ~new_n25676_ & ~new_n25674_ & ~new_n25684_;
  assign new_n25702_ = (new_n15282_ | ~new_n25653_ | ~new_n25652_) & (new_n25666_ | ~new_n25665_ | ~new_n25655_);
  assign new_n25703_ = new_n25704_ & (~new_n25748_ | (new_n25757_ & (new_n25758_ | new_n25754_)));
  assign new_n25704_ = new_n25705_ & (new_n25746_ | ~new_n25744_) & (~new_n11824_ | ~new_n25710_);
  assign new_n25705_ = (~new_n25706_ | ~new_n25708_) & (~new_n25707_ | ~new_n25709_);
  assign new_n25706_ = new_n20233_ & ~new_n21355_ & ~new_n7771_;
  assign new_n25707_ = ~new_n21355_ & ~new_n17931_ & ~new_n20233_;
  assign new_n25708_ = ~new_n15147_ & (~new_n15144_ | new_n15114_);
  assign new_n25709_ = ~new_n20402_ & ~new_n20405_;
  assign new_n25710_ = new_n25711_ & new_n21355_ & new_n21689_;
  assign new_n25711_ = ~new_n25712_ & new_n25739_;
  assign new_n25712_ = ~new_n25738_ & (~new_n25731_ | (~new_n25736_ & (new_n25729_ | new_n25737_ | ~new_n25713_)));
  assign new_n25713_ = ~new_n25725_ & ~new_n25723_ & ((~new_n25720_ & new_n25714_) | ~new_n25728_ | ~new_n25727_);
  assign new_n25714_ = \all_features[5951]  & \all_features[5950]  & ~new_n25717_ & new_n25715_;
  assign new_n25715_ = \all_features[5951]  & (\all_features[5950]  | (new_n25716_ & (\all_features[5946]  | \all_features[5947]  | \all_features[5945] )));
  assign new_n25716_ = \all_features[5948]  & \all_features[5949] ;
  assign new_n25717_ = new_n25719_ & ~\all_features[5949]  & ~new_n25718_ & ~\all_features[5948] ;
  assign new_n25718_ = \all_features[5944]  & \all_features[5945] ;
  assign new_n25719_ = ~\all_features[5946]  & ~\all_features[5947] ;
  assign new_n25720_ = \all_features[5951]  & \all_features[5950]  & ~new_n25721_ & \all_features[5949] ;
  assign new_n25721_ = ~\all_features[5947]  & ~\all_features[5948]  & (~\all_features[5946]  | new_n25722_);
  assign new_n25722_ = ~\all_features[5944]  & ~\all_features[5945] ;
  assign new_n25723_ = ~new_n25724_ & ~\all_features[5951] ;
  assign new_n25724_ = \all_features[5949]  & \all_features[5950]  & (\all_features[5948]  | (\all_features[5946]  & \all_features[5947]  & \all_features[5945] ));
  assign new_n25725_ = ~\all_features[5951]  & (~\all_features[5950]  | ~new_n25726_ | ~new_n25718_ | ~new_n25716_);
  assign new_n25726_ = \all_features[5946]  & \all_features[5947] ;
  assign new_n25727_ = \all_features[5951]  & (\all_features[5950]  | (\all_features[5949]  & (\all_features[5948]  | ~new_n25719_ | ~new_n25722_)));
  assign new_n25728_ = \all_features[5951]  & (\all_features[5949]  | \all_features[5950]  | \all_features[5948] );
  assign new_n25729_ = ~new_n25723_ & (new_n25725_ | (new_n25728_ & (~new_n25727_ | (~new_n25730_ & new_n25715_))));
  assign new_n25730_ = ~\all_features[5949]  & \all_features[5950]  & \all_features[5951]  & (\all_features[5948]  ? new_n25719_ : (new_n25718_ | ~new_n25719_));
  assign new_n25731_ = ~new_n25735_ & ~new_n25732_ & ~new_n25734_;
  assign new_n25732_ = new_n25733_ & (~\all_features[5949]  | (~\all_features[5948]  & (~\all_features[5947]  | (~\all_features[5946]  & ~\all_features[5945] ))));
  assign new_n25733_ = ~\all_features[5950]  & ~\all_features[5951] ;
  assign new_n25734_ = ~\all_features[5949]  & new_n25733_ & ((~\all_features[5946]  & new_n25722_) | ~\all_features[5948]  | ~\all_features[5947] );
  assign new_n25735_ = new_n25733_ & (~\all_features[5947]  | ~new_n25716_ | (~\all_features[5946]  & ~new_n25718_));
  assign new_n25736_ = ~\all_features[5951]  & (~\all_features[5950]  | (~\all_features[5948]  & ~\all_features[5949]  & ~new_n25726_));
  assign new_n25737_ = ~\all_features[5951]  & (~\all_features[5950]  | (~\all_features[5949]  & (new_n25722_ | ~\all_features[5948]  | ~new_n25726_)));
  assign new_n25738_ = ~\all_features[5951]  & ~\all_features[5950]  & ~\all_features[5949]  & ~\all_features[5947]  & ~\all_features[5948] ;
  assign new_n25739_ = new_n25732_ | ~new_n25742_ | ((new_n25723_ | ~new_n25743_) & (new_n25740_ | new_n25735_));
  assign new_n25740_ = new_n25741_ & (~new_n25714_ | ~new_n25727_ | ~new_n25728_);
  assign new_n25741_ = ~new_n25725_ & ~new_n25723_ & ~new_n25736_ & ~new_n25737_;
  assign new_n25742_ = ~new_n25734_ & ~new_n25738_;
  assign new_n25743_ = ~new_n25735_ & ~new_n25725_ & ~new_n25736_ & ~new_n25737_;
  assign new_n25744_ = new_n21355_ & ~new_n21689_ & ~new_n25745_;
  assign new_n25745_ = new_n16558_ & new_n21391_;
  assign new_n25746_ = new_n18164_ & new_n25747_;
  assign new_n25747_ = new_n12601_ & new_n12624_;
  assign new_n25748_ = new_n25749_ & (new_n14084_ | ~new_n25752_) & (~new_n25751_ | new_n25753_);
  assign new_n25749_ = (new_n15757_ | ~new_n25750_) & (~new_n25744_ | ~new_n25746_);
  assign new_n25750_ = new_n17931_ & ~new_n20233_ & ~new_n21355_;
  assign new_n25751_ = new_n25745_ & ~new_n21689_ & new_n21355_;
  assign new_n25752_ = new_n21355_ & ~new_n25711_ & new_n21689_;
  assign new_n25753_ = ~new_n12029_ & (~new_n12007_ | new_n16652_);
  assign new_n25754_ = ~new_n25755_ & (new_n25756_ | ((~new_n25753_ | ~new_n25751_) & (~new_n25752_ | ~new_n14084_)));
  assign new_n25755_ = ~new_n25708_ & new_n25706_;
  assign new_n25756_ = new_n25750_ & new_n15757_;
  assign new_n25757_ = (new_n25709_ | ~new_n25707_) & (new_n11824_ | ~new_n25710_);
  assign new_n25758_ = new_n7771_ & new_n20233_ & ~new_n9689_ & ~new_n21355_;
  assign new_n25759_ = new_n25760_ ? (new_n25812_ ^ new_n25906_) : (~new_n25812_ ^ new_n25906_);
  assign new_n25760_ = ~new_n25809_ & new_n25761_;
  assign new_n25761_ = new_n25762_ & ((new_n14290_ & new_n25807_) | new_n25806_ | ~new_n25805_);
  assign new_n25762_ = new_n25763_ & (new_n25767_ | ((new_n10037_ | new_n24447_) & (new_n25765_ | new_n9761_ | ~new_n24447_)));
  assign new_n25763_ = (~new_n25770_ | ~new_n25764_) & (~new_n25768_ | (new_n12908_ ? new_n16282_ : new_n25804_));
  assign new_n25764_ = new_n24447_ & ~new_n25767_ & new_n25765_;
  assign new_n25765_ = ~new_n15247_ & (~new_n20103_ | new_n25766_);
  assign new_n25766_ = ~new_n22444_ & ~new_n22448_;
  assign new_n25767_ = ~new_n21524_ & new_n21493_;
  assign new_n25768_ = ~new_n25769_ & new_n25767_;
  assign new_n25769_ = ~new_n12354_ & (~new_n14177_ | ~new_n14164_);
  assign new_n25770_ = new_n25771_ & ~new_n25796_ & ~new_n25800_;
  assign new_n25771_ = ~new_n25772_ & ~new_n25794_;
  assign new_n25772_ = new_n25789_ & ~new_n25793_ & ~new_n25773_ & ~new_n25792_;
  assign new_n25773_ = new_n25774_ & (~new_n25787_ | ~new_n25788_ | ~new_n25784_ | ~new_n25786_);
  assign new_n25774_ = ~new_n25781_ & ~new_n25779_ & ~new_n25775_ & ~new_n25777_;
  assign new_n25775_ = ~\all_features[1623]  & (~\all_features[1622]  | (~\all_features[1620]  & ~\all_features[1621]  & ~new_n25776_));
  assign new_n25776_ = \all_features[1618]  & \all_features[1619] ;
  assign new_n25777_ = ~\all_features[1623]  & (~\all_features[1622]  | (~\all_features[1621]  & (new_n25778_ | ~new_n25776_ | ~\all_features[1620] )));
  assign new_n25778_ = ~\all_features[1616]  & ~\all_features[1617] ;
  assign new_n25779_ = ~new_n25780_ & ~\all_features[1623] ;
  assign new_n25780_ = \all_features[1621]  & \all_features[1622]  & (\all_features[1620]  | (\all_features[1618]  & \all_features[1619]  & \all_features[1617] ));
  assign new_n25781_ = ~\all_features[1623]  & (~\all_features[1622]  | ~new_n25782_ | ~new_n25783_ | ~new_n25776_);
  assign new_n25782_ = \all_features[1616]  & \all_features[1617] ;
  assign new_n25783_ = \all_features[1620]  & \all_features[1621] ;
  assign new_n25784_ = \all_features[1623]  & (\all_features[1622]  | (\all_features[1621]  & (\all_features[1620]  | ~new_n25785_ | ~new_n25778_)));
  assign new_n25785_ = ~\all_features[1618]  & ~\all_features[1619] ;
  assign new_n25786_ = \all_features[1623]  & (\all_features[1622]  | (new_n25783_ & (\all_features[1618]  | \all_features[1619]  | \all_features[1617] )));
  assign new_n25787_ = \all_features[1622]  & \all_features[1623]  & (\all_features[1620]  | \all_features[1621]  | new_n25782_ | ~new_n25785_);
  assign new_n25788_ = \all_features[1623]  & (\all_features[1621]  | \all_features[1622]  | \all_features[1620] );
  assign new_n25789_ = ~new_n25790_ & (\all_features[1619]  | \all_features[1620]  | \all_features[1621]  | \all_features[1622]  | \all_features[1623] );
  assign new_n25790_ = ~\all_features[1621]  & new_n25791_ & ((~\all_features[1618]  & new_n25778_) | ~\all_features[1620]  | ~\all_features[1619] );
  assign new_n25791_ = ~\all_features[1622]  & ~\all_features[1623] ;
  assign new_n25792_ = new_n25791_ & (~\all_features[1621]  | (~\all_features[1620]  & (~\all_features[1619]  | (~\all_features[1618]  & ~\all_features[1617] ))));
  assign new_n25793_ = new_n25791_ & (~\all_features[1619]  | ~new_n25783_ | (~\all_features[1618]  & ~new_n25782_));
  assign new_n25794_ = new_n25795_ & new_n25789_ & ~new_n25792_ & ~new_n25779_;
  assign new_n25795_ = ~new_n25781_ & ~new_n25777_ & ~new_n25793_ & ~new_n25775_;
  assign new_n25796_ = ~new_n25797_ & (\all_features[1619]  | \all_features[1620]  | \all_features[1621]  | \all_features[1622]  | \all_features[1623] );
  assign new_n25797_ = ~new_n25790_ & (new_n25792_ | (~new_n25793_ & (new_n25775_ | (~new_n25798_ & ~new_n25777_))));
  assign new_n25798_ = ~new_n25779_ & (new_n25781_ | (new_n25788_ & (~new_n25784_ | (~new_n25799_ & new_n25786_))));
  assign new_n25799_ = ~\all_features[1621]  & \all_features[1622]  & \all_features[1623]  & (\all_features[1620]  ? new_n25785_ : (new_n25782_ | ~new_n25785_));
  assign new_n25800_ = new_n25789_ & (new_n25793_ | new_n25792_ | (~new_n25801_ & ~new_n25775_ & ~new_n25777_));
  assign new_n25801_ = ~new_n25779_ & ~new_n25781_ & (~new_n25788_ | ~new_n25784_ | new_n25802_);
  assign new_n25802_ = new_n25786_ & new_n25787_ & (new_n25803_ | ~\all_features[1621]  | ~\all_features[1622]  | ~\all_features[1623] );
  assign new_n25803_ = ~\all_features[1619]  & ~\all_features[1620]  & (~\all_features[1618]  | new_n25778_);
  assign new_n25804_ = new_n12112_ & new_n12115_;
  assign new_n25805_ = new_n25767_ & new_n25769_;
  assign new_n25806_ = ~new_n25807_ & (new_n17802_ | ~new_n25808_);
  assign new_n25807_ = ~new_n10432_ & (~new_n10409_ | ~new_n23071_);
  assign new_n25808_ = ~new_n17800_ & ~new_n17791_;
  assign new_n25809_ = new_n25811_ & new_n25810_ & (new_n25770_ | ~new_n25764_);
  assign new_n25810_ = (~new_n25806_ | ~new_n25805_) & (~new_n25768_ | (new_n12908_ ? ~new_n16282_ : ~new_n25804_));
  assign new_n25811_ = (~new_n10037_ | new_n24447_ | new_n25767_) & (~new_n25807_ | ~new_n14290_ | ~new_n25769_ | ~new_n25767_);
  assign new_n25812_ = ~new_n25813_ & new_n25901_;
  assign new_n25813_ = ~new_n25855_ & new_n25814_ & (new_n25900_ | ~new_n25865_);
  assign new_n25814_ = (new_n14426_ | new_n25823_ | new_n25817_) & (~new_n25817_ | (new_n25656_ ? ~new_n25816_ : ~new_n25815_));
  assign new_n25815_ = new_n13887_ & new_n19604_;
  assign new_n25816_ = ~new_n9209_ & ~new_n20155_;
  assign new_n25817_ = ~new_n21524_ & ~new_n21521_ & ~new_n25818_ & ~new_n21494_;
  assign new_n25818_ = ~new_n21509_ & (new_n21507_ | (~new_n21512_ & (new_n21511_ | new_n25819_)));
  assign new_n25819_ = ~new_n21514_ & (new_n21516_ | (~new_n21519_ & (new_n21518_ | new_n25820_)));
  assign new_n25820_ = ~new_n25821_ & \all_features[1271]  & (\all_features[1270]  | \all_features[1269]  | \all_features[1268] );
  assign new_n25821_ = \all_features[1271]  & ((~new_n25822_ & ~\all_features[1269]  & \all_features[1270] ) | (~new_n21501_ & (\all_features[1270]  | (~new_n21497_ & \all_features[1269] ))));
  assign new_n25822_ = (\all_features[1268]  & ~new_n21499_) | (~new_n21504_ & ~\all_features[1268]  & new_n21499_);
  assign new_n25823_ = ~new_n25853_ & (new_n25850_ | new_n25824_ | new_n25844_ | new_n25847_ | ~new_n25854_);
  assign new_n25824_ = new_n25843_ & (new_n25849_ | (~new_n25848_ & new_n25838_ & (new_n25841_ | new_n25825_)));
  assign new_n25825_ = ~new_n25832_ & (~new_n25836_ | (new_n25826_ & (~new_n25835_ | (~new_n25837_ & new_n25829_))));
  assign new_n25826_ = \all_features[5415]  & (\all_features[5414]  | new_n25827_);
  assign new_n25827_ = \all_features[5413]  & (\all_features[5410]  | \all_features[5411]  | \all_features[5412]  | ~new_n25828_);
  assign new_n25828_ = ~\all_features[5408]  & ~\all_features[5409] ;
  assign new_n25829_ = \all_features[5415]  & ~new_n25830_ & \all_features[5414] ;
  assign new_n25830_ = ~\all_features[5413]  & ~\all_features[5412]  & ~\all_features[5411]  & ~new_n25831_ & ~\all_features[5410] ;
  assign new_n25831_ = \all_features[5408]  & \all_features[5409] ;
  assign new_n25832_ = ~\all_features[5415]  & (~\all_features[5414]  | ~new_n25833_ | ~new_n25831_ | ~new_n25834_);
  assign new_n25833_ = \all_features[5410]  & \all_features[5411] ;
  assign new_n25834_ = \all_features[5412]  & \all_features[5413] ;
  assign new_n25835_ = \all_features[5415]  & (\all_features[5414]  | (new_n25834_ & (\all_features[5410]  | \all_features[5411]  | \all_features[5409] )));
  assign new_n25836_ = \all_features[5415]  & (\all_features[5413]  | \all_features[5414]  | \all_features[5412] );
  assign new_n25837_ = \all_features[5414]  & \all_features[5415]  & (\all_features[5413]  | (\all_features[5412]  & (\all_features[5411]  | \all_features[5410] )));
  assign new_n25838_ = ~new_n25832_ & ~new_n25841_ & (~new_n25836_ | new_n25839_ | ~new_n25826_);
  assign new_n25839_ = ~new_n25830_ & new_n25835_ & \all_features[5414]  & \all_features[5415]  & (~\all_features[5413]  | new_n25840_);
  assign new_n25840_ = ~\all_features[5411]  & ~\all_features[5412]  & (~\all_features[5410]  | new_n25828_);
  assign new_n25841_ = ~new_n25842_ & ~\all_features[5415] ;
  assign new_n25842_ = \all_features[5413]  & \all_features[5414]  & (\all_features[5412]  | (\all_features[5410]  & \all_features[5411]  & \all_features[5409] ));
  assign new_n25843_ = ~new_n25847_ & ~new_n25844_ & ~new_n25846_;
  assign new_n25844_ = new_n25845_ & (~\all_features[5413]  | (~\all_features[5412]  & (~\all_features[5411]  | (~\all_features[5410]  & ~\all_features[5409] ))));
  assign new_n25845_ = ~\all_features[5414]  & ~\all_features[5415] ;
  assign new_n25846_ = ~\all_features[5413]  & new_n25845_ & ((~\all_features[5410]  & new_n25828_) | ~\all_features[5412]  | ~\all_features[5411] );
  assign new_n25847_ = new_n25845_ & (~\all_features[5411]  | ~new_n25834_ | (~\all_features[5410]  & ~new_n25831_));
  assign new_n25848_ = ~\all_features[5415]  & (~\all_features[5414]  | (~\all_features[5413]  & (new_n25828_ | ~new_n25833_ | ~\all_features[5412] )));
  assign new_n25849_ = ~\all_features[5415]  & (~\all_features[5414]  | (~\all_features[5412]  & ~\all_features[5413]  & ~new_n25833_));
  assign new_n25850_ = ~new_n25841_ & ~new_n25848_ & new_n25852_ & (~new_n25826_ | ~new_n25851_);
  assign new_n25851_ = new_n25836_ & new_n25829_ & new_n25835_;
  assign new_n25852_ = ~new_n25832_ & ~new_n25849_;
  assign new_n25853_ = new_n25852_ & new_n25854_ & ~new_n25847_ & ~new_n25848_ & ~new_n25841_ & ~new_n25844_;
  assign new_n25854_ = ~new_n25846_ & (\all_features[5411]  | \all_features[5412]  | \all_features[5413]  | \all_features[5414]  | \all_features[5415] );
  assign new_n25855_ = new_n25656_ & new_n25817_ & ((new_n20155_ & ~new_n9209_) | (new_n23034_ & new_n25856_ & new_n9209_));
  assign new_n25856_ = ~new_n25857_ & ~new_n25861_;
  assign new_n25857_ = new_n23053_ & (~new_n23059_ | (~new_n25858_ & ~new_n23047_ & ~new_n23051_));
  assign new_n25858_ = ~new_n23052_ & ~new_n23045_ & (~new_n23043_ | ~new_n23049_ | new_n25859_);
  assign new_n25859_ = new_n23038_ & new_n23040_ & (new_n25860_ | ~\all_features[2293]  | ~\all_features[2294]  | ~\all_features[2295] );
  assign new_n25860_ = ~\all_features[2291]  & ~\all_features[2292]  & (~\all_features[2290]  | new_n23050_);
  assign new_n25861_ = ~new_n25862_ & (\all_features[2291]  | \all_features[2292]  | \all_features[2293]  | \all_features[2294]  | \all_features[2295] );
  assign new_n25862_ = ~new_n23054_ & (new_n23056_ | (~new_n23057_ & (new_n23047_ | (~new_n23051_ & ~new_n25863_))));
  assign new_n25863_ = ~new_n23045_ & (new_n23052_ | (new_n23043_ & (~new_n23049_ | (~new_n25864_ & new_n23038_))));
  assign new_n25864_ = ~\all_features[2293]  & \all_features[2294]  & \all_features[2295]  & (\all_features[2292]  ? new_n23041_ : (new_n23042_ | ~new_n23041_));
  assign new_n25865_ = new_n25866_ & ~new_n25817_ & new_n14426_;
  assign new_n25866_ = new_n25867_ & ~new_n25896_ & ~new_n25899_;
  assign new_n25867_ = ~new_n25868_ & ~new_n25892_;
  assign new_n25868_ = new_n25889_ & (~new_n25883_ | (~new_n25869_ & ~new_n25887_ & ~new_n25891_));
  assign new_n25869_ = ~new_n25880_ & ~new_n25879_ & (~new_n25882_ | ~new_n25878_ | new_n25870_);
  assign new_n25870_ = new_n25871_ & new_n25873_ & (new_n25876_ | ~\all_features[1637]  | ~\all_features[1638]  | ~\all_features[1639] );
  assign new_n25871_ = \all_features[1639]  & (\all_features[1638]  | (new_n25872_ & (\all_features[1634]  | \all_features[1635]  | \all_features[1633] )));
  assign new_n25872_ = \all_features[1636]  & \all_features[1637] ;
  assign new_n25873_ = \all_features[1638]  & \all_features[1639]  & (\all_features[1636]  | \all_features[1637]  | new_n25874_ | ~new_n25875_);
  assign new_n25874_ = \all_features[1632]  & \all_features[1633] ;
  assign new_n25875_ = ~\all_features[1634]  & ~\all_features[1635] ;
  assign new_n25876_ = ~\all_features[1635]  & ~\all_features[1636]  & (~\all_features[1634]  | new_n25877_);
  assign new_n25877_ = ~\all_features[1632]  & ~\all_features[1633] ;
  assign new_n25878_ = \all_features[1639]  & (\all_features[1638]  | (\all_features[1637]  & (\all_features[1636]  | ~new_n25877_ | ~new_n25875_)));
  assign new_n25879_ = ~\all_features[1639]  & (~new_n25872_ | ~\all_features[1634]  | ~\all_features[1635]  | ~\all_features[1638]  | ~new_n25874_);
  assign new_n25880_ = ~new_n25881_ & ~\all_features[1639] ;
  assign new_n25881_ = \all_features[1637]  & \all_features[1638]  & (\all_features[1636]  | (\all_features[1634]  & \all_features[1635]  & \all_features[1633] ));
  assign new_n25882_ = \all_features[1639]  & (\all_features[1637]  | \all_features[1638]  | \all_features[1636] );
  assign new_n25883_ = ~new_n25884_ & ~new_n25886_;
  assign new_n25884_ = new_n25885_ & (~\all_features[1635]  | ~new_n25872_ | (~\all_features[1634]  & ~new_n25874_));
  assign new_n25885_ = ~\all_features[1638]  & ~\all_features[1639] ;
  assign new_n25886_ = new_n25885_ & (~\all_features[1637]  | (~\all_features[1636]  & (~\all_features[1635]  | (~\all_features[1634]  & ~\all_features[1633] ))));
  assign new_n25887_ = ~\all_features[1639]  & (~\all_features[1638]  | new_n25888_);
  assign new_n25888_ = ~\all_features[1637]  & (new_n25877_ | ~\all_features[1635]  | ~\all_features[1636]  | ~\all_features[1634] );
  assign new_n25889_ = ~new_n25890_ & (\all_features[1635]  | \all_features[1636]  | \all_features[1637]  | \all_features[1638]  | \all_features[1639] );
  assign new_n25890_ = ~\all_features[1637]  & new_n25885_ & ((~\all_features[1634]  & new_n25877_) | ~\all_features[1636]  | ~\all_features[1635] );
  assign new_n25891_ = ~\all_features[1639]  & (~\all_features[1638]  | (~\all_features[1637]  & ~\all_features[1636]  & (~\all_features[1635]  | ~\all_features[1634] )));
  assign new_n25892_ = ~new_n25893_ & (\all_features[1635]  | \all_features[1636]  | \all_features[1637]  | \all_features[1638]  | \all_features[1639] );
  assign new_n25893_ = ~new_n25890_ & (new_n25886_ | (~new_n25884_ & (new_n25891_ | (~new_n25887_ & ~new_n25894_))));
  assign new_n25894_ = ~new_n25880_ & (new_n25879_ | (new_n25882_ & (~new_n25878_ | (~new_n25895_ & new_n25871_))));
  assign new_n25895_ = ~\all_features[1637]  & \all_features[1638]  & \all_features[1639]  & (\all_features[1636]  ? new_n25875_ : (new_n25874_ | ~new_n25875_));
  assign new_n25896_ = new_n25883_ & new_n25889_ & (new_n25887_ | new_n25897_ | new_n25879_ | ~new_n25898_);
  assign new_n25897_ = new_n25882_ & new_n25878_ & new_n25871_ & new_n25873_;
  assign new_n25898_ = ~new_n25880_ & ~new_n25891_;
  assign new_n25899_ = new_n25883_ & new_n25898_ & new_n25889_ & ~new_n25887_ & ~new_n25879_;
  assign new_n25900_ = ~new_n11062_ & ~new_n11094_;
  assign new_n25901_ = ~new_n25904_ & ~new_n25902_ & (~new_n25900_ | ~new_n25865_);
  assign new_n25902_ = ~new_n25656_ & new_n25817_ & (new_n19604_ ? ~new_n13887_ : ~new_n25903_);
  assign new_n25903_ = new_n20246_ & ~new_n15473_ & ~new_n15477_;
  assign new_n25904_ = ~new_n25817_ & ((new_n25823_ & ~new_n14426_) | (~new_n25866_ & new_n14426_ & (new_n25905_ | ~new_n14759_)));
  assign new_n25905_ = new_n21953_ & new_n21957_;
  assign new_n25906_ = ~new_n25907_ & ~new_n25909_;
  assign new_n25907_ = new_n21705_ & ((~new_n21689_ & new_n25908_) | (~new_n15674_ & new_n11897_ & ~new_n25908_));
  assign new_n25908_ = ~new_n12187_ & (~new_n12185_ | new_n16566_);
  assign new_n25909_ = new_n21705_ & new_n25908_ & ~new_n21689_ & ~new_n25746_;
  assign new_n25910_ = ~new_n25925_ & new_n25911_;
  assign new_n25911_ = new_n25921_ ? ((~new_n25912_ & ~new_n25914_ & new_n25922_) | (~new_n25923_ & ~new_n25922_)) : new_n25916_;
  assign new_n25912_ = ~new_n22548_ & new_n25913_;
  assign new_n25913_ = ~new_n24459_ & ~new_n24489_;
  assign new_n25914_ = ~new_n25915_ & ~new_n25913_;
  assign new_n25915_ = new_n15366_ & new_n24558_;
  assign new_n25916_ = (new_n25919_ | new_n7803_ | ~new_n25917_) & (~new_n13406_ | new_n25917_ | (new_n25920_ & new_n12733_));
  assign new_n25917_ = ~new_n11623_ & new_n25918_;
  assign new_n25918_ = ~new_n8963_ & ~new_n8985_;
  assign new_n25919_ = new_n14679_ & (new_n14656_ | (new_n14682_ & new_n14686_));
  assign new_n25920_ = new_n8924_ & new_n8927_;
  assign new_n25921_ = ~new_n21387_ | (~new_n21388_ & new_n21356_);
  assign new_n25922_ = new_n13503_ & (new_n13480_ | new_n13505_);
  assign new_n25923_ = ~new_n9967_ & new_n9995_ & (new_n6908_ | ~new_n25924_);
  assign new_n25924_ = ~new_n6886_ & ~new_n6910_;
  assign new_n25925_ = ~new_n13406_ & ~new_n25921_ & ~new_n25917_;
  assign new_n25926_ = new_n25927_ ? (~new_n25999_ ^ new_n25910_) : (new_n25999_ ^ new_n25910_);
  assign new_n25927_ = new_n25928_ ? (new_n25952_ ^ new_n25970_) : (~new_n25952_ ^ new_n25970_);
  assign new_n25928_ = new_n25948_ & (new_n25951_ | ~new_n25929_);
  assign new_n25929_ = ~new_n25943_ & new_n25930_ & (~new_n25947_ | ~new_n20499_ | ~new_n25946_);
  assign new_n25930_ = ~new_n25931_ & (~new_n25942_ | (~new_n12758_ & ~new_n19501_));
  assign new_n25931_ = new_n25932_ & new_n25935_ & new_n20852_ & (new_n24010_ | ~new_n25936_);
  assign new_n25932_ = ~new_n19162_ & new_n25933_;
  assign new_n25933_ = new_n25794_ & new_n25934_ & new_n25772_;
  assign new_n25934_ = new_n25796_ & new_n25800_;
  assign new_n25935_ = new_n9234_ & new_n23153_ & new_n9211_;
  assign new_n25936_ = ~new_n24019_ & ~new_n25937_;
  assign new_n25937_ = ~new_n20866_ & (new_n20860_ | (~new_n20864_ & (new_n20857_ | (~new_n25938_ & ~new_n20861_))));
  assign new_n25938_ = ~new_n20854_ & (new_n20862_ | (~new_n20865_ & (~new_n25941_ | new_n25939_)));
  assign new_n25939_ = \all_features[3527]  & ((~new_n25940_ & ~\all_features[3525]  & \all_features[3526] ) | (~new_n24015_ & (\all_features[3526]  | (~new_n24013_ & \all_features[3525] ))));
  assign new_n25940_ = (~\all_features[3522]  & ~\all_features[3523]  & ~\all_features[3524]  & (~\all_features[3521]  | ~\all_features[3520] )) | (\all_features[3524]  & (\all_features[3522]  | \all_features[3523] ));
  assign new_n25941_ = \all_features[3527]  & (\all_features[3525]  | \all_features[3526]  | \all_features[3524] );
  assign new_n25942_ = ~new_n20405_ & new_n19162_;
  assign new_n25943_ = new_n25944_ & (new_n20116_ ? new_n25945_ : new_n23174_);
  assign new_n25944_ = new_n19162_ & new_n20405_;
  assign new_n25945_ = new_n19599_ & (~new_n19600_ | ~new_n14008_);
  assign new_n25946_ = ~new_n19162_ & ~new_n25933_;
  assign new_n25947_ = ~new_n22423_ & (~new_n22420_ | ~new_n22391_);
  assign new_n25948_ = new_n25950_ & new_n25949_ & (new_n25945_ | ~new_n20116_ | ~new_n25944_);
  assign new_n25949_ = (~new_n25932_ | new_n25935_) & (new_n12758_ | new_n19501_ | ~new_n25942_);
  assign new_n25950_ = ~new_n25946_ | (new_n25947_ ? new_n20499_ : new_n18109_);
  assign new_n25951_ = (new_n25947_ | ~new_n25946_ | ~new_n18109_) & (new_n20116_ | new_n23174_ | ~new_n25944_);
  assign new_n25952_ = ~new_n25966_ & new_n25953_;
  assign new_n25953_ = ~new_n25960_ & new_n25954_ & (~new_n25965_ | ~new_n25964_);
  assign new_n25954_ = new_n25957_ | ((new_n25933_ | ~new_n25956_) & (new_n25959_ | ~new_n25955_));
  assign new_n25955_ = ~new_n16267_ & new_n16956_;
  assign new_n25956_ = ~new_n16956_ & (new_n15195_ | (new_n15172_ & new_n15198_));
  assign new_n25957_ = ~new_n25958_ & new_n25210_;
  assign new_n25958_ = ~new_n19085_ & ~new_n25338_;
  assign new_n25959_ = ~new_n6908_ & (~new_n6886_ | new_n6909_);
  assign new_n25960_ = new_n25957_ & ((~new_n25961_ & ~new_n23324_) | (~new_n19821_ & new_n25963_ & new_n23324_));
  assign new_n25961_ = (~new_n25962_ & ~new_n16282_) | (new_n20974_ & new_n10739_ & new_n10761_ & new_n16282_);
  assign new_n25962_ = ~new_n7769_ & (~new_n7767_ | new_n18589_);
  assign new_n25963_ = new_n15244_ & new_n15237_ & new_n15264_;
  assign new_n25964_ = new_n23324_ & ~new_n25963_ & new_n25957_;
  assign new_n25965_ = new_n23785_ & new_n24457_;
  assign new_n25966_ = ~new_n25969_ & ~new_n25968_ & (new_n25957_ | (new_n25967_ & ~new_n25956_) | (~new_n25933_ & new_n25956_));
  assign new_n25967_ = ~new_n25959_ & new_n25955_;
  assign new_n25968_ = ~new_n25965_ & new_n25964_;
  assign new_n25969_ = new_n25957_ & ~new_n16282_ & ~new_n23324_ & ~new_n25962_;
  assign new_n25970_ = new_n25971_ & new_n25998_;
  assign new_n25971_ = new_n18902_ & ((new_n25933_ & new_n25997_ & ~new_n25972_) | (new_n25972_ & (new_n25988_ | ~new_n25974_)));
  assign new_n25972_ = ~new_n25973_ & ~new_n17659_;
  assign new_n25973_ = new_n17637_ & new_n17667_;
  assign new_n25974_ = ~new_n25986_ & new_n16612_ & (~new_n25983_ | (~new_n25984_ & new_n25975_));
  assign new_n25975_ = new_n25976_ & ~new_n25983_ & ~new_n25979_ & ~new_n25981_;
  assign new_n25976_ = \all_features[2495]  | (\all_features[2494]  & (\all_features[2493]  | (~new_n25978_ & \all_features[2492]  & new_n25977_)));
  assign new_n25977_ = \all_features[2490]  & \all_features[2491] ;
  assign new_n25978_ = ~\all_features[2488]  & ~\all_features[2489] ;
  assign new_n25979_ = ~\all_features[2495]  & (~new_n25980_ | ~\all_features[2492]  | ~\all_features[2493]  | ~\all_features[2494]  | ~new_n25977_);
  assign new_n25980_ = \all_features[2488]  & \all_features[2489] ;
  assign new_n25981_ = ~new_n25982_ & ~\all_features[2495] ;
  assign new_n25982_ = \all_features[2493]  & \all_features[2494]  & (\all_features[2492]  | (\all_features[2490]  & \all_features[2491]  & \all_features[2489] ));
  assign new_n25983_ = ~\all_features[2495]  & ~\all_features[2494]  & ~\all_features[2493]  & ~\all_features[2491]  & ~\all_features[2492] ;
  assign new_n25984_ = ~\all_features[2495]  & ~new_n25985_ & ~\all_features[2494] ;
  assign new_n25985_ = \all_features[2491]  & \all_features[2492]  & \all_features[2493]  & (\all_features[2490]  | new_n25980_);
  assign new_n25986_ = ~\all_features[2495]  & ~\all_features[2494]  & ~new_n25987_ & ~\all_features[2493] ;
  assign new_n25987_ = \all_features[2491]  & \all_features[2492]  & (\all_features[2490]  | ~new_n25978_);
  assign new_n25988_ = new_n25989_ & (~new_n25976_ | (~new_n25995_ & ~new_n25979_ & ~new_n25981_ & new_n25983_));
  assign new_n25989_ = ~new_n25984_ & ~new_n25990_ & ~new_n25981_ & new_n25994_ & (~new_n25993_ | ~new_n25991_);
  assign new_n25990_ = ~\all_features[2495]  & (~\all_features[2494]  | (~\all_features[2493]  & (new_n25978_ | ~\all_features[2492]  | ~new_n25977_)));
  assign new_n25991_ = \all_features[2495]  & (\all_features[2494]  | (\all_features[2493]  & (\all_features[2492]  | ~new_n25992_ | ~new_n25978_)));
  assign new_n25992_ = ~\all_features[2490]  & ~\all_features[2491] ;
  assign new_n25993_ = \all_features[2494]  & \all_features[2495]  & (\all_features[2492]  | \all_features[2493]  | new_n25980_ | ~new_n25992_);
  assign new_n25994_ = \all_features[2495]  | (new_n25980_ & \all_features[2492]  & \all_features[2493]  & \all_features[2494]  & new_n25977_);
  assign new_n25995_ = new_n25991_ & (~new_n25993_ | (~new_n25996_ & \all_features[2493]  & \all_features[2494]  & \all_features[2495] ));
  assign new_n25996_ = ~\all_features[2491]  & ~\all_features[2492]  & (~\all_features[2490]  | new_n25978_);
  assign new_n25997_ = ~\all_features[5774]  & ~\all_features[5775]  & (~\all_features[5773]  | ~\all_features[5772]  | ~\all_features[5771] );
  assign new_n25998_ = new_n18902_ & (new_n25972_ | (new_n25933_ & new_n25997_) | (new_n16998_ & ~new_n25997_));
  assign new_n25999_ = ~new_n26000_ & new_n26043_;
  assign new_n26000_ = ~new_n26039_ & ~new_n26001_ & new_n26003_ & (~new_n26042_ | ~new_n26041_);
  assign new_n26001_ = new_n26002_ & new_n6884_;
  assign new_n26002_ = ~new_n19279_ & new_n13887_;
  assign new_n26003_ = ~new_n26004_ | (new_n26038_ ? new_n26005_ : ~new_n19195_);
  assign new_n26004_ = ~new_n13887_ & ~new_n19279_;
  assign new_n26005_ = ~new_n26037_ & ~new_n26034_ & ~new_n26006_ & ~new_n26027_;
  assign new_n26006_ = ~new_n26007_ & (\all_features[2051]  | \all_features[2052]  | \all_features[2053]  | \all_features[2054]  | \all_features[2055] );
  assign new_n26007_ = ~new_n26021_ & (new_n26023_ | (~new_n26024_ & (new_n26025_ | (~new_n26008_ & ~new_n26026_))));
  assign new_n26008_ = ~new_n26009_ & (new_n26011_ | (new_n26020_ & (~new_n26015_ | (~new_n26019_ & new_n26018_))));
  assign new_n26009_ = ~new_n26010_ & ~\all_features[2055] ;
  assign new_n26010_ = \all_features[2053]  & \all_features[2054]  & (\all_features[2052]  | (\all_features[2050]  & \all_features[2051]  & \all_features[2049] ));
  assign new_n26011_ = ~\all_features[2055]  & (~\all_features[2054]  | ~new_n26012_ | ~new_n26013_ | ~new_n26014_);
  assign new_n26012_ = \all_features[2048]  & \all_features[2049] ;
  assign new_n26013_ = \all_features[2052]  & \all_features[2053] ;
  assign new_n26014_ = \all_features[2050]  & \all_features[2051] ;
  assign new_n26015_ = \all_features[2055]  & (\all_features[2054]  | (\all_features[2053]  & (\all_features[2052]  | ~new_n26017_ | ~new_n26016_)));
  assign new_n26016_ = ~\all_features[2048]  & ~\all_features[2049] ;
  assign new_n26017_ = ~\all_features[2050]  & ~\all_features[2051] ;
  assign new_n26018_ = \all_features[2055]  & (\all_features[2054]  | (new_n26013_ & (\all_features[2050]  | \all_features[2051]  | \all_features[2049] )));
  assign new_n26019_ = ~\all_features[2053]  & \all_features[2054]  & \all_features[2055]  & (\all_features[2052]  ? new_n26017_ : (new_n26012_ | ~new_n26017_));
  assign new_n26020_ = \all_features[2055]  & (\all_features[2053]  | \all_features[2054]  | \all_features[2052] );
  assign new_n26021_ = ~\all_features[2053]  & new_n26022_ & ((~\all_features[2050]  & new_n26016_) | ~\all_features[2052]  | ~\all_features[2051] );
  assign new_n26022_ = ~\all_features[2054]  & ~\all_features[2055] ;
  assign new_n26023_ = new_n26022_ & (~\all_features[2053]  | (~\all_features[2052]  & (~\all_features[2051]  | (~\all_features[2050]  & ~\all_features[2049] ))));
  assign new_n26024_ = new_n26022_ & (~\all_features[2051]  | ~new_n26013_ | (~\all_features[2050]  & ~new_n26012_));
  assign new_n26025_ = ~\all_features[2055]  & (~\all_features[2054]  | (~\all_features[2052]  & ~\all_features[2053]  & ~new_n26014_));
  assign new_n26026_ = ~\all_features[2055]  & (~\all_features[2054]  | (~\all_features[2053]  & (new_n26016_ | ~new_n26014_ | ~\all_features[2052] )));
  assign new_n26027_ = new_n26033_ & (~new_n26032_ | (~new_n26028_ & ~new_n26025_ & ~new_n26026_));
  assign new_n26028_ = ~new_n26009_ & ~new_n26011_ & (~new_n26020_ | ~new_n26015_ | new_n26029_);
  assign new_n26029_ = new_n26018_ & new_n26030_ & (new_n26031_ | ~\all_features[2053]  | ~\all_features[2054]  | ~\all_features[2055] );
  assign new_n26030_ = \all_features[2054]  & \all_features[2055]  & (\all_features[2052]  | \all_features[2053]  | new_n26012_ | ~new_n26017_);
  assign new_n26031_ = ~\all_features[2051]  & ~\all_features[2052]  & (~\all_features[2050]  | new_n26016_);
  assign new_n26032_ = ~new_n26023_ & ~new_n26024_;
  assign new_n26033_ = ~new_n26021_ & (\all_features[2051]  | \all_features[2052]  | \all_features[2053]  | \all_features[2054]  | \all_features[2055] );
  assign new_n26034_ = new_n26032_ & new_n26033_ & (new_n26035_ | new_n26026_ | new_n26011_ | ~new_n26036_);
  assign new_n26035_ = new_n26020_ & new_n26030_ & new_n26015_ & new_n26018_;
  assign new_n26036_ = ~new_n26025_ & ~new_n26009_;
  assign new_n26037_ = new_n26033_ & new_n26032_ & new_n26036_ & ~new_n26026_ & ~new_n26011_;
  assign new_n26038_ = ~new_n19190_ & (~new_n19164_ | ~new_n19191_);
  assign new_n26039_ = new_n19279_ & (new_n21722_ ? new_n26040_ : (~new_n15762_ | ~new_n9833_));
  assign new_n26040_ = ~new_n10204_ & (~new_n10201_ | new_n10168_);
  assign new_n26041_ = new_n21722_ & ~new_n26040_ & new_n19279_;
  assign new_n26042_ = ~new_n20580_ & new_n11906_;
  assign new_n26043_ = new_n26044_ & (new_n26042_ | ~new_n26041_) & (~new_n26002_ | new_n6884_);
  assign new_n26044_ = ~new_n26004_ | (new_n26038_ ? ~new_n26005_ : new_n19195_);
  assign new_n26045_ = new_n25953_ & new_n25966_;
  assign new_n26046_ = new_n26047_ ? (~new_n26045_ ^ new_n26156_) : (new_n26045_ ^ new_n26156_);
  assign new_n26047_ = new_n26048_ ? (new_n26081_ ^ new_n26150_) : (~new_n26081_ ^ new_n26150_);
  assign new_n26048_ = new_n26049_ ? (new_n26057_ ^ new_n26076_) : (~new_n26057_ ^ new_n26076_);
  assign new_n26049_ = new_n26050_ & (~new_n25903_ | new_n26055_);
  assign new_n26050_ = ~new_n26051_ & (new_n25903_ | ((new_n26054_ | new_n9966_) & (new_n23319_ | new_n26042_ | ~new_n9966_)));
  assign new_n26051_ = new_n25903_ & ~new_n26053_ & ~new_n24395_ & ~new_n26052_;
  assign new_n26052_ = new_n24158_ & new_n25918_;
  assign new_n26053_ = new_n18752_ & new_n19315_;
  assign new_n26054_ = (~new_n9936_ & ~new_n8132_ & (~new_n8099_ | ~new_n8129_)) | (~new_n20966_ & new_n18575_ & (new_n8132_ | (new_n8099_ & new_n8129_)));
  assign new_n26055_ = (new_n26056_ | new_n18797_ | new_n21245_ | ~new_n24395_) & (~new_n25422_ | ~new_n26052_ | new_n24395_);
  assign new_n26056_ = ~new_n21211_ & new_n21242_;
  assign new_n26057_ = ~new_n26058_ & ~new_n26075_;
  assign new_n26058_ = new_n26059_ & (~new_n26074_ | ~new_n19813_) & (~new_n19888_ | (new_n26070_ & new_n26073_));
  assign new_n26059_ = ~new_n26060_ & (new_n19888_ | (~new_n26062_ & new_n26063_ & new_n10906_) | (new_n26064_ & ~new_n10906_));
  assign new_n26060_ = new_n19888_ & new_n25770_ & ~new_n26061_ & new_n20578_;
  assign new_n26061_ = ~new_n18396_ & new_n20584_;
  assign new_n26062_ = ~new_n6848_ & new_n8542_;
  assign new_n26063_ = ~new_n13196_ & (~new_n13170_ | ~new_n20801_);
  assign new_n26064_ = new_n13130_ & ~new_n26065_ & new_n13127_;
  assign new_n26065_ = ~new_n13100_ & (new_n13115_ | (~new_n13113_ & (new_n13118_ | (~new_n13117_ & ~new_n26066_))));
  assign new_n26066_ = ~new_n13120_ & (new_n13122_ | (~new_n13125_ & (new_n13124_ | (~new_n26067_ & new_n26069_))));
  assign new_n26067_ = \all_features[5687]  & ((~new_n26068_ & ~\all_features[5685]  & \all_features[5686] ) | (~new_n13107_ & (\all_features[5686]  | (~new_n13103_ & \all_features[5685] ))));
  assign new_n26068_ = (\all_features[5684]  & ~new_n13105_) | (~new_n13110_ & ~\all_features[5684]  & new_n13105_);
  assign new_n26069_ = \all_features[5687]  & (\all_features[5685]  | \all_features[5686]  | \all_features[5684] );
  assign new_n26070_ = (~new_n26071_ | new_n20578_) & (new_n23598_ | ~new_n26061_ | ~new_n20578_);
  assign new_n26071_ = new_n26072_ & new_n6953_ & (new_n6950_ | new_n6921_);
  assign new_n26072_ = new_n16448_ & new_n16418_ & new_n16446_;
  assign new_n26073_ = (new_n26072_ | new_n20578_) & (new_n25770_ | new_n26061_ | ~new_n20578_);
  assign new_n26074_ = new_n26064_ & ~new_n19888_ & ~new_n10906_;
  assign new_n26075_ = ~new_n19813_ & new_n26074_;
  assign new_n26076_ = new_n18582_ & (new_n26077_ | (~new_n26078_ & (new_n15588_ ? new_n26080_ : new_n22837_)));
  assign new_n26077_ = new_n26078_ & ((new_n14679_ & new_n20241_ & (new_n14656_ | ~new_n14681_)) | (new_n26079_ & ~new_n20241_));
  assign new_n26078_ = ~new_n14751_ & new_n14726_;
  assign new_n26079_ = ~new_n15990_ & (~new_n15986_ | new_n15957_);
  assign new_n26080_ = new_n20767_ & new_n20761_ & new_n20768_ & new_n20739_;
  assign new_n26081_ = new_n26082_ ? (new_n26129_ ^ new_n26142_) : (~new_n26129_ ^ new_n26142_);
  assign new_n26082_ = ~new_n26083_ & new_n26127_;
  assign new_n26083_ = new_n26093_ & (new_n26125_ | (new_n26084_ & ~new_n26126_) | (~new_n26091_ & new_n26126_));
  assign new_n26084_ = new_n16646_ ? (new_n20080_ | (~new_n26086_ & new_n20077_)) : new_n26085_;
  assign new_n26085_ = ~new_n11333_ & (~new_n11335_ | ~new_n12265_);
  assign new_n26086_ = ~new_n20052_ & ~new_n26087_;
  assign new_n26087_ = ~new_n26088_ & (\all_features[5427]  | \all_features[5428]  | \all_features[5429]  | \all_features[5430]  | \all_features[5431] );
  assign new_n26088_ = ~new_n20073_ & (new_n20069_ | (~new_n20071_ & (new_n20065_ | (~new_n20067_ & ~new_n26089_))));
  assign new_n26089_ = ~new_n20074_ & (new_n20076_ | (new_n20063_ & (~new_n20062_ | (~new_n26090_ & new_n20057_))));
  assign new_n26090_ = ~\all_features[5429]  & \all_features[5430]  & \all_features[5431]  & (\all_features[5428]  ? new_n20061_ : (new_n20060_ | ~new_n20061_));
  assign new_n26091_ = new_n26092_ ? ~new_n13063_ : new_n15530_;
  assign new_n26092_ = new_n23035_ & new_n23058_;
  assign new_n26093_ = ~new_n26125_ | (new_n16997_ ? (new_n22545_ ? ~new_n23548_ : ~new_n14276_) : new_n26094_);
  assign new_n26094_ = (new_n11783_ | ~new_n19139_ | (new_n25059_ & new_n18192_)) & (new_n26095_ | new_n26122_ | (~new_n11783_ & new_n19139_));
  assign new_n26095_ = ~new_n26119_ & ~new_n26117_ & ~new_n26121_ & (new_n26120_ | (new_n26114_ & new_n26096_));
  assign new_n26096_ = ~new_n26108_ & ~new_n26113_ & (new_n26112_ | new_n26110_ | new_n26097_);
  assign new_n26097_ = new_n26101_ & new_n26107_ & (~new_n26105_ | ~new_n26103_ | new_n26098_);
  assign new_n26098_ = \all_features[2263]  & \all_features[2262]  & ~new_n26099_ & \all_features[2261] ;
  assign new_n26099_ = ~\all_features[2259]  & ~\all_features[2260]  & (~\all_features[2258]  | new_n26100_);
  assign new_n26100_ = ~\all_features[2256]  & ~\all_features[2257] ;
  assign new_n26101_ = \all_features[2263]  & (\all_features[2262]  | (\all_features[2261]  & (\all_features[2260]  | ~new_n26102_ | ~new_n26100_)));
  assign new_n26102_ = ~\all_features[2258]  & ~\all_features[2259] ;
  assign new_n26103_ = \all_features[2263]  & (\all_features[2262]  | (new_n26104_ & (\all_features[2258]  | \all_features[2259]  | \all_features[2257] )));
  assign new_n26104_ = \all_features[2260]  & \all_features[2261] ;
  assign new_n26105_ = \all_features[2262]  & \all_features[2263]  & (\all_features[2260]  | \all_features[2261]  | new_n26106_ | ~new_n26102_);
  assign new_n26106_ = \all_features[2256]  & \all_features[2257] ;
  assign new_n26107_ = \all_features[2263]  & (\all_features[2261]  | \all_features[2262]  | \all_features[2260] );
  assign new_n26108_ = ~\all_features[2263]  & (~\all_features[2262]  | (~\all_features[2261]  & (new_n26100_ | ~\all_features[2260]  | ~new_n26109_)));
  assign new_n26109_ = \all_features[2258]  & \all_features[2259] ;
  assign new_n26110_ = ~new_n26111_ & ~\all_features[2263] ;
  assign new_n26111_ = \all_features[2261]  & \all_features[2262]  & (\all_features[2260]  | (\all_features[2258]  & \all_features[2259]  & \all_features[2257] ));
  assign new_n26112_ = ~\all_features[2263]  & (~\all_features[2262]  | ~new_n26109_ | ~new_n26106_ | ~new_n26104_);
  assign new_n26113_ = ~\all_features[2263]  & (~\all_features[2262]  | (~\all_features[2260]  & ~\all_features[2261]  & ~new_n26109_));
  assign new_n26114_ = ~new_n26113_ & (new_n26108_ | (~new_n26115_ & ~new_n26110_));
  assign new_n26115_ = ~new_n26112_ & (~new_n26107_ | (new_n26101_ & (~new_n26103_ | (~new_n26116_ & new_n26105_))));
  assign new_n26116_ = \all_features[2262]  & \all_features[2263]  & (\all_features[2261]  | (~new_n26102_ & \all_features[2260] ));
  assign new_n26117_ = new_n26118_ & (~\all_features[2261]  | (~\all_features[2260]  & (~\all_features[2259]  | (~\all_features[2258]  & ~\all_features[2257] ))));
  assign new_n26118_ = ~\all_features[2262]  & ~\all_features[2263] ;
  assign new_n26119_ = ~\all_features[2261]  & new_n26118_ & ((~\all_features[2258]  & new_n26100_) | ~\all_features[2260]  | ~\all_features[2259] );
  assign new_n26120_ = new_n26118_ & (~\all_features[2259]  | ~new_n26104_ | (~\all_features[2258]  & ~new_n26106_));
  assign new_n26121_ = ~\all_features[2263]  & ~\all_features[2262]  & ~\all_features[2261]  & ~\all_features[2259]  & ~\all_features[2260] ;
  assign new_n26122_ = ~new_n26121_ & ~new_n26120_ & ~new_n26117_ & ~new_n26119_;
  assign new_n26125_ = ~new_n14119_ & (~new_n14122_ | ~new_n14091_);
  assign new_n26126_ = new_n11884_ & (new_n11861_ | new_n11886_);
  assign new_n26127_ = (~new_n26128_ | ~new_n26126_ | new_n26125_) & (new_n22545_ | new_n14276_ | ~new_n16997_ | ~new_n26125_);
  assign new_n26128_ = ~new_n26092_ & ~new_n15530_;
  assign new_n26129_ = new_n26137_ & (new_n26140_ | new_n26130_);
  assign new_n26130_ = ~new_n25903_ & (new_n26136_ ? (new_n26132_ ? ~new_n26134_ : new_n26133_) : ~new_n26131_);
  assign new_n26131_ = new_n16899_ & new_n20482_;
  assign new_n26132_ = ~new_n11901_ & (~new_n21842_ | ~new_n17013_);
  assign new_n26133_ = ~new_n6597_ & new_n18577_;
  assign new_n26134_ = new_n22711_ & new_n26135_;
  assign new_n26135_ = ~new_n14505_ & ~new_n14528_;
  assign new_n26136_ = new_n23879_ & (~new_n16356_ | ~new_n9968_);
  assign new_n26137_ = (new_n18574_ | new_n16899_ | new_n26136_ | new_n25903_) & (~new_n26139_ | ~new_n26138_ | ~new_n25903_);
  assign new_n26138_ = ~new_n7557_ & (~new_n8701_ | ~new_n9688_);
  assign new_n26139_ = new_n18421_ & (~new_n18451_ | ~new_n18447_);
  assign new_n26140_ = new_n25903_ & (new_n26141_ | new_n26139_ | (new_n6908_ & (new_n6886_ | ~new_n6909_)));
  assign new_n26141_ = new_n20080_ & (new_n20077_ | (new_n20052_ & new_n26087_));
  assign new_n26142_ = new_n26143_ & new_n26149_;
  assign new_n26143_ = new_n21705_ & (new_n26144_ | (new_n15170_ & new_n26148_));
  assign new_n26144_ = ~new_n26145_ & (new_n10774_ | ~new_n26147_ | ~new_n18324_);
  assign new_n26145_ = new_n26146_ & new_n26006_ & new_n26027_;
  assign new_n26146_ = new_n26034_ & new_n26037_;
  assign new_n26147_ = ~new_n11497_ & ~new_n11496_ & ~new_n11493_ & ~new_n11494_;
  assign new_n26148_ = new_n10911_ & new_n26145_;
  assign new_n26149_ = new_n21705_ & (new_n26148_ | new_n26144_);
  assign new_n26150_ = new_n26151_ & new_n26155_;
  assign new_n26151_ = new_n26153_ & (~new_n26152_ | ~new_n21917_ | ~new_n24042_);
  assign new_n26152_ = (~new_n12562_ & (new_n14046_ | (new_n15163_ & new_n14072_))) | (new_n25973_ & new_n17659_ & ~new_n14046_ & (~new_n15163_ | ~new_n14072_));
  assign new_n26153_ = (new_n21917_ & new_n24042_) | (new_n26154_ & ~new_n24042_ & (new_n22443_ ? ~new_n16758_ : new_n23133_));
  assign new_n26154_ = new_n11301_ & (new_n11274_ | new_n13767_);
  assign new_n26155_ = (~new_n21917_ | new_n26152_ | ~new_n24042_) & (new_n16758_ | ~new_n26154_ | ~new_n22443_ | new_n24042_);
  assign new_n26156_ = ~new_n26155_ & new_n26151_;
  assign new_n26157_ = new_n26158_ & new_n26173_;
  assign new_n26158_ = new_n26159_ & (~new_n26171_ | (new_n18887_ & new_n26170_) | (new_n26172_ & ~new_n26170_));
  assign new_n26159_ = ~new_n26160_ & (new_n15549_ | ~new_n26163_ | (new_n6884_ ? new_n13516_ : new_n26169_));
  assign new_n26160_ = new_n26164_ & ~new_n26161_ & new_n26162_;
  assign new_n26161_ = new_n22923_ & new_n24948_ & new_n24027_;
  assign new_n26162_ = ~new_n14923_ & ~new_n26163_;
  assign new_n26163_ = ~new_n25700_ & ~new_n25690_ & ~new_n25696_;
  assign new_n26164_ = new_n16023_ & (new_n15993_ | new_n26165_);
  assign new_n26165_ = ~new_n16017_ & new_n16018_ & (new_n16016_ | (~new_n26166_ & ~new_n16014_));
  assign new_n26166_ = ~new_n16012_ & (new_n16002_ | (~new_n16004_ & (new_n16005_ | (~new_n26167_ & ~new_n16007_))));
  assign new_n26167_ = new_n16010_ & (~new_n15995_ | (new_n16009_ & (new_n26168_ | ~new_n15998_)));
  assign new_n26168_ = \all_features[4662]  & \all_features[4663]  & (\all_features[4661]  | (\all_features[4660]  & (\all_features[4659]  | \all_features[4658] )));
  assign new_n26169_ = new_n21483_ & new_n21451_ & new_n21478_;
  assign new_n26170_ = ~new_n18110_ & new_n19836_;
  assign new_n26171_ = ~new_n26163_ & new_n14923_;
  assign new_n26172_ = ~new_n10728_ & new_n16526_;
  assign new_n26173_ = new_n26174_ & (~new_n26171_ | (~new_n18887_ & new_n26170_) | (~new_n26172_ & ~new_n26170_));
  assign new_n26174_ = new_n26175_ & (~new_n26162_ | (~new_n26161_ & new_n26164_) | (~new_n15364_ & ~new_n26164_));
  assign new_n26175_ = ~new_n26163_ | ((~new_n6884_ | ~new_n13516_ | new_n15549_) & (~new_n15549_ | (new_n26177_ & ~new_n26176_)));
  assign new_n26176_ = ~new_n16890_ & (~new_n16887_ | ~new_n16879_);
  assign new_n26177_ = ~new_n26203_ & ~new_n26178_ & ~new_n26201_;
  assign new_n26178_ = new_n26188_ & (~new_n26191_ | (new_n26194_ & (new_n26179_ | new_n26198_ | new_n26199_)));
  assign new_n26179_ = new_n26180_ & (~new_n26183_ | (~new_n26187_ & \all_features[1653]  & \all_features[1654]  & \all_features[1655] ));
  assign new_n26180_ = \all_features[1655]  & (\all_features[1654]  | (~new_n26181_ & \all_features[1653] ));
  assign new_n26181_ = new_n26182_ & ~\all_features[1652]  & ~\all_features[1650]  & ~\all_features[1651] ;
  assign new_n26182_ = ~\all_features[1648]  & ~\all_features[1649] ;
  assign new_n26183_ = \all_features[1655]  & \all_features[1654]  & ~new_n26186_ & new_n26184_;
  assign new_n26184_ = \all_features[1655]  & (\all_features[1654]  | (new_n26185_ & (\all_features[1650]  | \all_features[1651]  | \all_features[1649] )));
  assign new_n26185_ = \all_features[1652]  & \all_features[1653] ;
  assign new_n26186_ = ~\all_features[1650]  & ~\all_features[1651]  & ~\all_features[1652]  & ~\all_features[1653]  & (~\all_features[1649]  | ~\all_features[1648] );
  assign new_n26187_ = ~\all_features[1651]  & ~\all_features[1652]  & (~\all_features[1650]  | new_n26182_);
  assign new_n26188_ = ~new_n26189_ & (\all_features[1651]  | \all_features[1652]  | \all_features[1653]  | \all_features[1654]  | \all_features[1655] );
  assign new_n26189_ = ~\all_features[1653]  & new_n26190_ & ((~\all_features[1650]  & new_n26182_) | ~\all_features[1652]  | ~\all_features[1651] );
  assign new_n26190_ = ~\all_features[1654]  & ~\all_features[1655] ;
  assign new_n26191_ = ~new_n26192_ & ~new_n26193_;
  assign new_n26192_ = new_n26190_ & (~new_n26185_ | ~\all_features[1651]  | (~\all_features[1650]  & (~\all_features[1648]  | ~\all_features[1649] )));
  assign new_n26193_ = new_n26190_ & (~\all_features[1653]  | (~\all_features[1652]  & (~\all_features[1651]  | (~\all_features[1650]  & ~\all_features[1649] ))));
  assign new_n26194_ = ~new_n26195_ & ~new_n26197_;
  assign new_n26195_ = ~\all_features[1655]  & (~\all_features[1654]  | (~\all_features[1652]  & ~\all_features[1653]  & ~new_n26196_));
  assign new_n26196_ = \all_features[1650]  & \all_features[1651] ;
  assign new_n26197_ = ~\all_features[1655]  & (~\all_features[1654]  | (~\all_features[1653]  & (new_n26182_ | ~new_n26196_ | ~\all_features[1652] )));
  assign new_n26198_ = ~\all_features[1655]  & (~new_n26196_ | ~\all_features[1648]  | ~\all_features[1649]  | ~\all_features[1654]  | ~new_n26185_);
  assign new_n26199_ = ~new_n26200_ & ~\all_features[1655] ;
  assign new_n26200_ = \all_features[1653]  & \all_features[1654]  & (\all_features[1652]  | (\all_features[1650]  & \all_features[1651]  & \all_features[1649] ));
  assign new_n26201_ = new_n26191_ & ~new_n26202_ & new_n26188_;
  assign new_n26202_ = ~new_n26195_ & ~new_n26197_ & ~new_n26198_ & ~new_n26199_ & (~new_n26183_ | ~new_n26180_);
  assign new_n26203_ = new_n26191_ & new_n26188_ & new_n26194_ & ~new_n26198_ & ~new_n26199_;
  assign new_n26204_ = new_n26205_ ? (~new_n26257_ ^ new_n26277_) : (new_n26257_ ^ new_n26277_);
  assign new_n26205_ = new_n26206_ ? (~new_n26157_ ^ new_n26250_) : (new_n26157_ ^ new_n26250_);
  assign new_n26206_ = new_n26207_ ? (~new_n26237_ ^ new_n26150_) : (new_n26237_ ^ new_n26150_);
  assign new_n26207_ = new_n26208_ ? (new_n26218_ ^ new_n26236_) : (~new_n26218_ ^ new_n26236_);
  assign new_n26208_ = ~new_n26216_ & new_n26209_;
  assign new_n26209_ = ~new_n26210_ & (~new_n11902_ | ((new_n26211_ | ~new_n26212_) & (new_n26213_ | new_n26214_ | new_n26212_)));
  assign new_n26210_ = ~new_n14388_ & ~new_n11902_ & new_n12730_ & (~new_n20483_ | new_n12627_);
  assign new_n26211_ = (~new_n16156_ & new_n25407_ & (~new_n11857_ | new_n23968_)) | (new_n23814_ & new_n24456_ & (new_n16156_ | ~new_n25407_));
  assign new_n26212_ = ~new_n15921_ & new_n19341_;
  assign new_n26213_ = ~new_n25808_ & new_n17802_;
  assign new_n26214_ = new_n23947_ & new_n26215_;
  assign new_n26215_ = new_n14495_ & new_n14499_;
  assign new_n26216_ = ~new_n11902_ & ((~new_n26217_ & ~new_n12730_) | (~new_n23220_ & new_n14388_ & new_n8161_ & new_n12730_));
  assign new_n26217_ = (~new_n13356_ & new_n20263_ & new_n20800_) | (new_n22383_ & new_n12984_ & ~new_n20800_);
  assign new_n26218_ = ~new_n26219_ & new_n26234_;
  assign new_n26219_ = (new_n26227_ & (new_n26232_ ? new_n26226_ : ~new_n26233_)) | (new_n26225_ & new_n26220_ & ~new_n26227_);
  assign new_n26220_ = (~new_n26221_ | ~new_n26224_) & (~new_n22323_ | ~new_n26223_);
  assign new_n26221_ = ~new_n21569_ & new_n26222_;
  assign new_n26222_ = ~\all_features[5783]  & ~\all_features[5782]  & ~\all_features[5781]  & ~\all_features[5779]  & ~\all_features[5780] ;
  assign new_n26223_ = ~new_n19545_ & new_n21569_;
  assign new_n26224_ = new_n6627_ & (new_n6605_ | ~new_n6629_);
  assign new_n26225_ = (new_n26222_ | new_n21569_) & (~new_n19545_ | ~new_n14782_ | ~new_n21569_);
  assign new_n26226_ = ~new_n13243_ & (~new_n17998_ | (~new_n17976_ & new_n17999_));
  assign new_n26227_ = new_n19163_ & (~new_n26228_ | ~new_n19191_);
  assign new_n26228_ = ~new_n19184_ & (new_n19183_ | new_n26229_);
  assign new_n26229_ = ~new_n19179_ & (new_n19181_ | (~new_n19174_ & (new_n19175_ | (~new_n19167_ & ~new_n26230_))));
  assign new_n26230_ = ~new_n19169_ & (~new_n19189_ | (new_n19188_ & (~new_n19185_ | (~new_n26231_ & new_n19186_))));
  assign new_n26231_ = \all_features[4438]  & \all_features[4439]  & (\all_features[4437]  | (~new_n19187_ & \all_features[4436] ));
  assign new_n26232_ = ~new_n12784_ & new_n18893_;
  assign new_n26233_ = (new_n22795_ & new_n23156_ & new_n25913_) | (~new_n14147_ & new_n25362_ & ~new_n25913_);
  assign new_n26234_ = new_n26227_ ? (new_n26232_ ? ~new_n26226_ : new_n26233_) : new_n26235_;
  assign new_n26235_ = (new_n22323_ | ~new_n26223_) & (new_n26224_ | ~new_n26221_);
  assign new_n26236_ = ~new_n25911_ & ~new_n25925_;
  assign new_n26237_ = ~new_n26238_ & new_n26247_;
  assign new_n26238_ = new_n26239_ & (~new_n10573_ | (new_n26244_ & new_n12264_) | (new_n26246_ & ~new_n12264_));
  assign new_n26239_ = new_n10573_ | (new_n25279_ ? ~new_n26240_ : (new_n24040_ ? new_n26241_ : new_n26242_));
  assign new_n26240_ = ~new_n23926_ & (new_n18631_ | (new_n18598_ & new_n18619_ & new_n18627_));
  assign new_n26241_ = ~new_n16652_ & new_n12006_;
  assign new_n26242_ = new_n10284_ & new_n26243_;
  assign new_n26243_ = ~new_n21610_ & ~new_n21606_;
  assign new_n26244_ = (new_n26245_ | new_n8093_) & (new_n26215_ | ~new_n14470_ | ~new_n8093_);
  assign new_n26245_ = new_n21559_ & (new_n21537_ | (new_n22786_ & new_n25658_));
  assign new_n26246_ = (~new_n9234_ | (~new_n9211_ & new_n9236_)) & (new_n14493_ | (~new_n14494_ & new_n14471_));
  assign new_n26247_ = ~new_n26249_ & ~new_n26248_ & (~new_n10573_ | (~new_n26244_ & new_n12264_) | (~new_n26246_ & ~new_n12264_));
  assign new_n26248_ = ~new_n10573_ & ~new_n26240_ & new_n25279_ & (~new_n23926_ | ~new_n8892_);
  assign new_n26249_ = ~new_n10573_ & ~new_n25279_ & (new_n24040_ ? new_n26241_ : new_n26242_);
  assign new_n26250_ = new_n26251_ & (new_n26256_ | new_n26253_ | new_n25771_);
  assign new_n26251_ = ~new_n26254_ & (~new_n26252_ | (new_n21048_ & (new_n21045_ | ~new_n21016_)));
  assign new_n26252_ = ~new_n25771_ & ~new_n9514_ & ~new_n9516_ & new_n26253_ & (~new_n9507_ | ~new_n9486_);
  assign new_n26253_ = new_n11672_ & (new_n11669_ | new_n11636_);
  assign new_n26254_ = new_n26255_ & (~new_n10936_ | (~new_n21199_ & ~new_n10912_));
  assign new_n26255_ = ~new_n26146_ & new_n25771_ & (new_n26228_ | ~new_n19162_);
  assign new_n26256_ = (~new_n25384_ & new_n19094_) | (new_n23608_ & new_n23632_ & new_n23630_ & ~new_n19094_);
  assign new_n26257_ = ~new_n26258_ & ~new_n26276_;
  assign new_n26258_ = new_n26259_ & (~new_n26275_ | (new_n26265_ & (new_n22374_ ? ~new_n26266_ : new_n12562_)));
  assign new_n26259_ = new_n26260_ & (~new_n26273_ | ~new_n26272_);
  assign new_n26260_ = ~new_n26267_ & new_n26261_ & ((~new_n23032_ & new_n23002_) | new_n26271_ | ~new_n26270_);
  assign new_n26261_ = (~new_n26265_ | ~new_n26266_ | ~new_n22374_) & (~new_n26264_ | ~new_n26262_);
  assign new_n26262_ = ~new_n26263_ & new_n25666_;
  assign new_n26263_ = new_n9458_ & new_n9340_;
  assign new_n26264_ = ~new_n20882_ & new_n17710_;
  assign new_n26265_ = new_n26263_ & new_n16377_;
  assign new_n26266_ = new_n22083_ & (new_n22080_ | ~new_n23870_);
  assign new_n26267_ = new_n26268_ & (new_n20800_ ? ~new_n10490_ : ~new_n26269_);
  assign new_n26268_ = ~new_n16377_ & new_n26263_;
  assign new_n26269_ = new_n13975_ & (new_n13971_ | new_n13964_);
  assign new_n26270_ = ~new_n25666_ & ~new_n26263_;
  assign new_n26271_ = ~new_n16562_ & (~new_n16559_ | new_n21391_);
  assign new_n26272_ = new_n26270_ & new_n26271_;
  assign new_n26273_ = ~new_n8132_ & (~new_n8129_ | new_n26274_);
  assign new_n26274_ = ~new_n8100_ & ~new_n8121_;
  assign new_n26275_ = (~new_n26262_ | new_n26264_) & (~new_n26268_ | (new_n20800_ ? ~new_n10490_ : ~new_n26269_));
  assign new_n26276_ = ~new_n26273_ & new_n26272_;
  assign new_n26277_ = ~new_n26278_ & ~new_n26290_;
  assign new_n26278_ = new_n26279_ & (~new_n26289_ | (~new_n16757_ & new_n25745_) | (new_n16946_ & ~new_n25745_));
  assign new_n26279_ = (~new_n26288_ & new_n26280_ & new_n8667_) | (~new_n8667_ & (new_n26287_ | (new_n24039_ & ~new_n15669_)));
  assign new_n26280_ = (~new_n26281_ & ~new_n18194_ & ~new_n18221_ & new_n25142_) | (~new_n25142_ & (new_n12685_ | new_n22877_));
  assign new_n26281_ = new_n26282_ & (new_n18216_ | (~new_n18214_ & (new_n18212_ | (~new_n18205_ & ~new_n26283_))));
  assign new_n26282_ = new_n18217_ & (\all_features[5323]  | \all_features[5324]  | \all_features[5325]  | \all_features[5326]  | \all_features[5327] );
  assign new_n26283_ = ~new_n18207_ & (new_n18208_ | (~new_n18210_ & (~new_n26286_ | new_n26284_)));
  assign new_n26284_ = \all_features[5327]  & ((~new_n26285_ & ~\all_features[5325]  & \all_features[5326] ) | (~new_n18201_ & (\all_features[5326]  | (~new_n18197_ & \all_features[5325] ))));
  assign new_n26285_ = (\all_features[5324]  & ~new_n18199_) | (~new_n18204_ & ~\all_features[5324]  & new_n18199_);
  assign new_n26286_ = \all_features[5327]  & (\all_features[5325]  | \all_features[5326]  | \all_features[5324] );
  assign new_n26287_ = new_n12595_ & ~new_n12563_ & new_n12592_;
  assign new_n26288_ = ~new_n21048_ & (~new_n21041_ | ~new_n21045_ | ~new_n21017_);
  assign new_n26289_ = ~new_n8667_ & new_n26287_;
  assign new_n26290_ = new_n25745_ & ~new_n16757_ & new_n26289_;
  assign new_n26291_ = ~new_n26173_ & new_n26158_;
  assign new_n26292_ = ~new_n26298_ & (~new_n26293_ | (~new_n26299_ & new_n26301_));
  assign new_n26293_ = ~new_n26294_ & (new_n26078_ | ((new_n26297_ | new_n22655_) & (new_n18161_ | new_n21245_ | ~new_n22655_)));
  assign new_n26294_ = new_n26295_ & new_n21689_;
  assign new_n26295_ = new_n26296_ & new_n23184_;
  assign new_n26296_ = ~new_n11725_ & new_n26078_;
  assign new_n26297_ = ~new_n26176_ & new_n8133_;
  assign new_n26298_ = ~new_n21689_ & new_n26295_;
  assign new_n26299_ = (~new_n25208_ | ~new_n26300_) & (new_n22655_ | new_n26078_ | ~new_n26297_);
  assign new_n26300_ = ~new_n23184_ & new_n26296_;
  assign new_n26301_ = new_n26302_ & (new_n25208_ | ~new_n26300_);
  assign new_n26302_ = new_n26303_ & (new_n26078_ | ~new_n22655_ | (new_n21245_ ? ~new_n26304_ : ~new_n18161_));
  assign new_n26303_ = ~new_n11725_ | ~new_n26078_;
  assign new_n26304_ = ~new_n13095_ & new_n13066_;
  assign new_n26305_ = new_n26351_ & (~new_n24810_ | ~new_n26353_ | ~new_n26306_ | ~new_n26309_);
  assign new_n26306_ = new_n26307_ & (~new_n26350_ | ~new_n26349_);
  assign new_n26307_ = ~new_n26308_ & (new_n26312_ | new_n26348_ | new_n12597_) & (~new_n23868_ | new_n26311_ | ~new_n12597_);
  assign new_n26308_ = new_n26310_ & ~new_n24810_ & new_n26309_;
  assign new_n26309_ = ~new_n23868_ & new_n12597_;
  assign new_n26310_ = ~new_n10726_ & (~new_n10703_ | new_n10728_);
  assign new_n26311_ = ~new_n13976_ & ~new_n24954_;
  assign new_n26312_ = new_n26313_ & new_n26342_;
  assign new_n26313_ = ~new_n26314_ & ~new_n26338_;
  assign new_n26314_ = new_n26329_ & (~new_n26334_ | (~new_n26332_ & ~new_n26315_ & ~new_n26337_));
  assign new_n26315_ = ~new_n26327_ & ~new_n26325_ & (~new_n26328_ | ~new_n26324_ | new_n26316_);
  assign new_n26316_ = new_n26317_ & new_n26321_ & (new_n26319_ | ~\all_features[5653]  | ~\all_features[5654]  | ~\all_features[5655] );
  assign new_n26317_ = \all_features[5655]  & (\all_features[5654]  | (new_n26318_ & (\all_features[5650]  | \all_features[5651]  | \all_features[5649] )));
  assign new_n26318_ = \all_features[5652]  & \all_features[5653] ;
  assign new_n26319_ = ~\all_features[5651]  & ~\all_features[5652]  & (~\all_features[5650]  | new_n26320_);
  assign new_n26320_ = ~\all_features[5648]  & ~\all_features[5649] ;
  assign new_n26321_ = \all_features[5654]  & \all_features[5655]  & (\all_features[5652]  | \all_features[5653]  | new_n26323_ | ~new_n26322_);
  assign new_n26322_ = ~\all_features[5650]  & ~\all_features[5651] ;
  assign new_n26323_ = \all_features[5648]  & \all_features[5649] ;
  assign new_n26324_ = \all_features[5655]  & (\all_features[5654]  | (\all_features[5653]  & (\all_features[5652]  | ~new_n26322_ | ~new_n26320_)));
  assign new_n26325_ = ~new_n26326_ & ~\all_features[5655] ;
  assign new_n26326_ = \all_features[5653]  & \all_features[5654]  & (\all_features[5652]  | (\all_features[5650]  & \all_features[5651]  & \all_features[5649] ));
  assign new_n26327_ = ~\all_features[5655]  & (~new_n26323_ | ~\all_features[5650]  | ~\all_features[5651]  | ~\all_features[5654]  | ~new_n26318_);
  assign new_n26328_ = \all_features[5655]  & (\all_features[5653]  | \all_features[5654]  | \all_features[5652] );
  assign new_n26329_ = ~new_n26330_ & (\all_features[5651]  | \all_features[5652]  | \all_features[5653]  | \all_features[5654]  | \all_features[5655] );
  assign new_n26330_ = ~\all_features[5653]  & new_n26331_ & ((~\all_features[5650]  & new_n26320_) | ~\all_features[5652]  | ~\all_features[5651] );
  assign new_n26331_ = ~\all_features[5654]  & ~\all_features[5655] ;
  assign new_n26332_ = ~\all_features[5655]  & (~\all_features[5654]  | new_n26333_);
  assign new_n26333_ = ~\all_features[5653]  & (new_n26320_ | ~\all_features[5651]  | ~\all_features[5652]  | ~\all_features[5650] );
  assign new_n26334_ = ~new_n26335_ & ~new_n26336_;
  assign new_n26335_ = new_n26331_ & (~\all_features[5653]  | (~\all_features[5652]  & (~\all_features[5651]  | (~\all_features[5650]  & ~\all_features[5649] ))));
  assign new_n26336_ = new_n26331_ & (~\all_features[5651]  | ~new_n26318_ | (~new_n26323_ & ~\all_features[5650] ));
  assign new_n26337_ = ~\all_features[5655]  & (~\all_features[5654]  | (~\all_features[5653]  & ~\all_features[5652]  & (~\all_features[5651]  | ~\all_features[5650] )));
  assign new_n26338_ = ~new_n26339_ & (\all_features[5651]  | \all_features[5652]  | \all_features[5653]  | \all_features[5654]  | \all_features[5655] );
  assign new_n26339_ = ~new_n26330_ & (new_n26335_ | (~new_n26336_ & (new_n26337_ | (~new_n26332_ & ~new_n26340_))));
  assign new_n26340_ = ~new_n26325_ & (new_n26327_ | (new_n26328_ & (~new_n26324_ | (~new_n26341_ & new_n26317_))));
  assign new_n26341_ = ~\all_features[5653]  & \all_features[5654]  & \all_features[5655]  & (\all_features[5652]  ? new_n26322_ : (new_n26323_ | ~new_n26322_));
  assign new_n26342_ = ~new_n26343_ & ~new_n26346_;
  assign new_n26343_ = new_n26334_ & ~new_n26344_ & new_n26329_;
  assign new_n26344_ = ~new_n26337_ & ~new_n26327_ & ~new_n26325_ & ~new_n26332_ & ~new_n26345_;
  assign new_n26345_ = new_n26328_ & new_n26324_ & new_n26317_ & new_n26321_;
  assign new_n26346_ = new_n26329_ & new_n26347_ & ~new_n26325_ & ~new_n26335_;
  assign new_n26347_ = ~new_n26337_ & ~new_n26336_ & ~new_n26332_ & ~new_n26327_;
  assign new_n26348_ = ~new_n6879_ & (~new_n19096_ | ~new_n19125_ | ~new_n19127_);
  assign new_n26349_ = ~new_n12597_ & new_n26312_;
  assign new_n26350_ = (new_n10910_ | new_n25708_) & (new_n20077_ | new_n20080_ | ~new_n26086_ | ~new_n25708_);
  assign new_n26351_ = new_n26352_ & (new_n26350_ | ~new_n26349_);
  assign new_n26352_ = ~new_n12597_ | (new_n23868_ ? ~new_n26311_ : (new_n24810_ ? new_n26353_ : new_n26310_));
  assign new_n26353_ = ~new_n26361_ & new_n26364_ & ((~new_n26365_ & ~\all_features[5911]  & new_n26367_) | (~new_n26354_ & (\all_features[5911]  | new_n26367_)));
  assign new_n26354_ = (new_n26355_ | \all_features[5911] ) & (new_n26360_ | ~\all_features[5910]  | ~\all_features[5911] );
  assign new_n26355_ = \all_features[5905]  & \all_features[5904]  & new_n26358_ & new_n26356_ & new_n26357_;
  assign new_n26356_ = \all_features[5906]  & \all_features[5907] ;
  assign new_n26357_ = \all_features[5909]  & \all_features[5910]  & (\all_features[5908]  | (\all_features[5906]  & \all_features[5907]  & \all_features[5905] ));
  assign new_n26358_ = \all_features[5908]  & \all_features[5910]  & ~\all_features[5911]  & \all_features[5909] ;
  assign new_n26360_ = ~\all_features[5906]  & ~\all_features[5907]  & ~\all_features[5908]  & ~\all_features[5909]  & (~\all_features[5905]  | ~\all_features[5904] );
  assign new_n26361_ = ~\all_features[5911]  & ~new_n26362_ & ~\all_features[5910] ;
  assign new_n26362_ = new_n26363_ & (\all_features[5907]  | \all_features[5908] ) & (\all_features[5906]  | (\all_features[5904]  & \all_features[5905] ));
  assign new_n26363_ = \all_features[5907]  & \all_features[5909]  & ~\all_features[5910]  & \all_features[5908] ;
  assign new_n26364_ = \all_features[5911]  | (new_n26366_ & new_n26357_ & new_n26365_);
  assign new_n26365_ = \all_features[5910]  & (\all_features[5908]  | \all_features[5909]  | new_n26356_);
  assign new_n26366_ = \all_features[5910]  & \all_features[5909]  & \all_features[5908]  & \all_features[5905]  & new_n26356_ & \all_features[5904] ;
  assign new_n26367_ = \all_features[5910]  & (\all_features[5909]  | (\all_features[5908]  & new_n26356_ & (\all_features[5905]  | \all_features[5904] )));
  assign new_n26368_ = ~new_n26382_ & new_n26369_;
  assign new_n26369_ = ~new_n26378_ & new_n26370_ & (~new_n26379_ | (~new_n22050_ & new_n26380_) | (new_n26381_ & ~new_n26380_));
  assign new_n26370_ = new_n26371_ & (~new_n26374_ | (new_n24041_ & new_n26376_) | (new_n26377_ & ~new_n26376_));
  assign new_n26371_ = new_n18578_ | ((new_n19340_ | ~new_n26372_ | ~new_n25549_) & (new_n26373_ | new_n25549_));
  assign new_n26372_ = new_n13012_ & (new_n13009_ | ~new_n22355_);
  assign new_n26373_ = new_n19497_ & (new_n19494_ | (new_n19470_ & new_n21717_));
  assign new_n26374_ = ~new_n26375_ & new_n18578_;
  assign new_n26375_ = ~new_n24180_ & ~new_n10682_;
  assign new_n26376_ = ~new_n6495_ & (~new_n6491_ | new_n20242_);
  assign new_n26377_ = ~new_n15198_ & new_n19380_;
  assign new_n26378_ = new_n25549_ & ~new_n21605_ & ~new_n26372_ & ~new_n18578_;
  assign new_n26379_ = new_n18578_ & new_n26375_;
  assign new_n26380_ = ~new_n26346_ & (~new_n26343_ | new_n26313_);
  assign new_n26381_ = ~new_n9634_ & (~new_n9612_ | new_n9635_);
  assign new_n26382_ = new_n26383_ & (~new_n26374_ | (~new_n24041_ & new_n26376_) | (~new_n26377_ & ~new_n26376_));
  assign new_n26383_ = ~new_n26385_ & (new_n18578_ | (new_n26384_ & new_n25549_) | (~new_n26373_ & ~new_n25549_));
  assign new_n26384_ = new_n26372_ ? ~new_n19340_ : ~new_n21605_;
  assign new_n26385_ = new_n26380_ & ~new_n22050_ & new_n26379_;
  assign new_n26386_ = new_n18582_ & (new_n26387_ | (new_n26388_ & (new_n26390_ | new_n16267_)));
  assign new_n26387_ = ~new_n26388_ & ((~new_n12936_ & new_n12909_) ? (~new_n14530_ & new_n26135_) : new_n21854_);
  assign new_n26388_ = new_n26389_ & new_n12115_;
  assign new_n26389_ = new_n12084_ & new_n12112_;
  assign new_n26390_ = new_n15147_ & new_n15115_ & new_n15144_;
  assign new_n26391_ = new_n26392_ & (new_n26449_ | ~new_n26446_);
  assign new_n26392_ = new_n26401_ & new_n26393_ & (~new_n26426_ | (~new_n26427_ & new_n12686_) | (new_n26431_ & ~new_n12686_));
  assign new_n26393_ = (~new_n26399_ | ~new_n26394_) & (~new_n26398_ | (new_n6919_ ? new_n26400_ : new_n25208_));
  assign new_n26394_ = ~new_n14349_ & new_n26395_;
  assign new_n26395_ = ~new_n26397_ & new_n26396_;
  assign new_n26396_ = new_n14919_ & new_n12253_;
  assign new_n26397_ = new_n25199_ & new_n22702_;
  assign new_n26398_ = new_n26396_ & new_n26397_;
  assign new_n26399_ = ~new_n20533_ & (~new_n20531_ | ~new_n20500_);
  assign new_n26400_ = new_n22443_ & new_n25766_;
  assign new_n26401_ = (~new_n26395_ | ~new_n14349_) & (new_n13887_ | new_n14388_ | ~new_n26402_);
  assign new_n26402_ = ~new_n26396_ & ~new_n26403_;
  assign new_n26403_ = ~new_n26424_ & ~new_n26404_ & ~new_n26422_;
  assign new_n26404_ = ~new_n26416_ & (new_n26418_ | (new_n26405_ & (new_n26410_ | new_n26419_ | new_n26420_)));
  assign new_n26405_ = ~new_n26406_ & ~new_n26408_;
  assign new_n26406_ = ~\all_features[2503]  & (~\all_features[2502]  | (~\all_features[2500]  & ~\all_features[2501]  & ~new_n26407_));
  assign new_n26407_ = \all_features[2498]  & \all_features[2499] ;
  assign new_n26408_ = ~\all_features[2503]  & (~\all_features[2502]  | (~\all_features[2501]  & (new_n26409_ | ~new_n26407_ | ~\all_features[2500] )));
  assign new_n26409_ = ~\all_features[2496]  & ~\all_features[2497] ;
  assign new_n26410_ = new_n26411_ & (~new_n26414_ | (~new_n26413_ & \all_features[2501]  & \all_features[2502]  & \all_features[2503] ));
  assign new_n26411_ = \all_features[2503]  & (\all_features[2502]  | (\all_features[2501]  & (\all_features[2500]  | ~new_n26412_ | ~new_n26409_)));
  assign new_n26412_ = ~\all_features[2498]  & ~\all_features[2499] ;
  assign new_n26413_ = ~\all_features[2499]  & ~\all_features[2500]  & (~\all_features[2498]  | new_n26409_);
  assign new_n26414_ = \all_features[2502]  & \all_features[2503]  & (\all_features[2500]  | \all_features[2501]  | new_n26415_ | ~new_n26412_);
  assign new_n26415_ = \all_features[2496]  & \all_features[2497] ;
  assign new_n26416_ = ~\all_features[2501]  & ~\all_features[2502]  & ~\all_features[2503]  & (~new_n26417_ | (~\all_features[2498]  & new_n26409_));
  assign new_n26417_ = \all_features[2499]  & \all_features[2500] ;
  assign new_n26418_ = ~\all_features[2502]  & ~\all_features[2503]  & (~\all_features[2501]  | ~new_n26417_ | (~\all_features[2498]  & ~new_n26415_));
  assign new_n26419_ = ~\all_features[2503]  & (~new_n26407_ | ~\all_features[2500]  | ~\all_features[2501]  | ~\all_features[2502]  | ~new_n26415_);
  assign new_n26420_ = ~new_n26421_ & ~\all_features[2503] ;
  assign new_n26421_ = \all_features[2501]  & \all_features[2502]  & (\all_features[2500]  | (\all_features[2498]  & \all_features[2499]  & \all_features[2497] ));
  assign new_n26422_ = new_n26405_ & new_n26423_ & ~new_n26420_ & ~new_n26416_ & ~new_n26419_;
  assign new_n26423_ = ~new_n26418_ & (\all_features[2499]  | \all_features[2500]  | \all_features[2501]  | \all_features[2502]  | \all_features[2503] );
  assign new_n26424_ = ~new_n26416_ & ~new_n26418_ & (~new_n26425_ | (new_n26411_ & new_n26414_));
  assign new_n26425_ = ~new_n26420_ & ~new_n26419_ & ~new_n26406_ & ~new_n26408_;
  assign new_n26426_ = ~new_n26396_ & new_n26403_;
  assign new_n26427_ = new_n24498_ & (new_n20659_ | (~new_n20658_ & (new_n20660_ | new_n26428_)));
  assign new_n26428_ = ~new_n20655_ & (new_n20647_ | (~new_n20653_ & (new_n20651_ | (~new_n20645_ & ~new_n26429_))));
  assign new_n26429_ = new_n20643_ & (~new_n20648_ | (new_n20641_ & (new_n26430_ | ~new_n20638_)));
  assign new_n26430_ = \all_features[5702]  & \all_features[5703]  & (\all_features[5701]  | (\all_features[5700]  & (\all_features[5699]  | \all_features[5698] )));
  assign new_n26431_ = ~new_n26439_ & new_n26442_ & ((~new_n26443_ & ~\all_features[3391]  & new_n26445_) | (~new_n26432_ & (\all_features[3391]  | new_n26445_)));
  assign new_n26432_ = (new_n26433_ | \all_features[3391] ) & (new_n26438_ | ~\all_features[3390]  | ~\all_features[3391] );
  assign new_n26433_ = \all_features[3385]  & \all_features[3384]  & new_n26436_ & new_n26434_ & new_n26435_;
  assign new_n26434_ = \all_features[3386]  & \all_features[3387] ;
  assign new_n26435_ = \all_features[3389]  & \all_features[3390]  & (\all_features[3388]  | (\all_features[3386]  & \all_features[3387]  & \all_features[3385] ));
  assign new_n26436_ = \all_features[3388]  & \all_features[3390]  & ~\all_features[3391]  & \all_features[3389] ;
  assign new_n26438_ = ~\all_features[3386]  & ~\all_features[3387]  & ~\all_features[3388]  & ~\all_features[3389]  & (~\all_features[3385]  | ~\all_features[3384] );
  assign new_n26439_ = ~\all_features[3391]  & ~new_n26440_ & ~\all_features[3390] ;
  assign new_n26440_ = new_n26441_ & (\all_features[3387]  | \all_features[3388] ) & (\all_features[3386]  | (\all_features[3384]  & \all_features[3385] ));
  assign new_n26441_ = \all_features[3387]  & \all_features[3389]  & ~\all_features[3390]  & \all_features[3388] ;
  assign new_n26442_ = \all_features[3391]  | (new_n26444_ & new_n26435_ & new_n26443_);
  assign new_n26443_ = \all_features[3390]  & (\all_features[3388]  | \all_features[3389]  | new_n26434_);
  assign new_n26444_ = \all_features[3390]  & \all_features[3389]  & \all_features[3388]  & \all_features[3385]  & new_n26434_ & \all_features[3384] ;
  assign new_n26445_ = \all_features[3390]  & (\all_features[3389]  | (\all_features[3388]  & new_n26434_ & (\all_features[3385]  | \all_features[3384] )));
  assign new_n26446_ = ~new_n26447_ & new_n26448_ & (new_n26399_ | ~new_n26394_);
  assign new_n26447_ = new_n26402_ & (new_n13887_ ? ~new_n13806_ : new_n14388_);
  assign new_n26448_ = (new_n6919_ | ~new_n26398_ | ~new_n25208_) & (new_n26427_ | ~new_n26426_ | ~new_n12686_);
  assign new_n26449_ = (~new_n26398_ | ~new_n26400_ | ~new_n6919_) & (new_n12686_ | ~new_n26426_ | ~new_n26431_);
  assign \o[50]  = new_n26451_ ? (new_n26452_ ^ new_n26511_) : (~new_n26452_ ^ new_n26511_);
  assign new_n26451_ = new_n25538_ & new_n26391_;
  assign new_n26452_ = new_n26453_ ? (~new_n26509_ ^ new_n26510_) : (new_n26509_ ^ new_n26510_);
  assign new_n26453_ = new_n26454_ ? (~new_n26507_ ^ new_n26508_) : (new_n26507_ ^ new_n26508_);
  assign new_n26454_ = new_n26455_ ? (new_n26493_ ^ new_n26494_) : (~new_n26493_ ^ new_n26494_);
  assign new_n26455_ = new_n26456_ ? (new_n26479_ ^ new_n26480_) : (~new_n26479_ ^ new_n26480_);
  assign new_n26456_ = new_n26457_ ? (new_n26466_ ^ new_n26478_) : (~new_n26466_ ^ new_n26478_);
  assign new_n26457_ = new_n26458_ ? (~new_n26464_ ^ new_n26465_) : (new_n26464_ ^ new_n26465_);
  assign new_n26458_ = new_n26459_ ? (new_n26462_ ^ new_n26463_) : (~new_n26462_ ^ new_n26463_);
  assign new_n26459_ = ~new_n26461_ & new_n26460_;
  assign new_n26460_ = ~new_n26298_ & new_n26293_;
  assign new_n26461_ = new_n26299_ & new_n26301_;
  assign new_n26462_ = new_n26306_ & new_n26351_;
  assign new_n26463_ = ~new_n25909_ & new_n25907_;
  assign new_n26464_ = (new_n25952_ & new_n25970_) | (new_n25928_ & (new_n25952_ | new_n25970_));
  assign new_n26465_ = (new_n25812_ & new_n25906_) | (new_n25760_ & (new_n25812_ | new_n25906_));
  assign new_n26466_ = new_n26467_ ? (new_n26471_ ^ new_n26472_) : (~new_n26471_ ^ new_n26472_);
  assign new_n26467_ = new_n26468_ ? (new_n26469_ ^ new_n26470_) : (~new_n26469_ ^ new_n26470_);
  assign new_n26468_ = new_n26369_ & new_n26382_;
  assign new_n26469_ = new_n25649_ & new_n25702_;
  assign new_n26470_ = new_n25813_ & new_n25901_;
  assign new_n26471_ = (new_n25648_ & new_n25703_) | (new_n25545_ & (new_n25648_ | new_n25703_));
  assign new_n26472_ = new_n26473_ ? (new_n26474_ ^ new_n26475_) : (~new_n26474_ ^ new_n26475_);
  assign new_n26473_ = new_n25623_ & new_n25546_ & (new_n25611_ | ~new_n25609_ | ~new_n25624_);
  assign new_n26474_ = new_n26392_ & new_n26446_;
  assign new_n26475_ = new_n26476_ & (~new_n26477_ | (~new_n25755_ & ~new_n25756_));
  assign new_n26476_ = new_n25704_ & new_n25748_;
  assign new_n26477_ = ~new_n25758_ & new_n25757_;
  assign new_n26478_ = (~new_n25759_ & new_n25910_) | (~new_n25544_ & (~new_n25759_ | new_n25910_));
  assign new_n26479_ = (~new_n25926_ & new_n26045_) | (~new_n25543_ & (~new_n25926_ | new_n26045_));
  assign new_n26480_ = new_n26481_ ? (~new_n26482_ ^ new_n26492_) : (new_n26482_ ^ new_n26492_);
  assign new_n26481_ = (~new_n26081_ & new_n26150_) | (~new_n26048_ & (~new_n26081_ | new_n26150_));
  assign new_n26482_ = new_n26483_ ? (new_n26487_ ^ new_n26491_) : (~new_n26487_ ^ new_n26491_);
  assign new_n26483_ = new_n26484_ ? (new_n26485_ ^ new_n26486_) : (~new_n26485_ ^ new_n26486_);
  assign new_n26484_ = ~new_n26276_ & new_n26259_;
  assign new_n26485_ = new_n25929_ & new_n25948_;
  assign new_n26486_ = new_n25761_ & new_n25809_;
  assign new_n26487_ = new_n26488_ ? (new_n26489_ ^ new_n26490_) : (~new_n26489_ ^ new_n26490_);
  assign new_n26488_ = ~new_n26290_ & new_n26278_;
  assign new_n26489_ = ~new_n26143_ & new_n26149_;
  assign new_n26490_ = ~new_n25971_ & new_n25998_;
  assign new_n26491_ = (new_n26129_ & new_n26142_) | (new_n26082_ & (new_n26129_ | new_n26142_));
  assign new_n26492_ = (new_n25999_ & new_n25910_) | (~new_n25927_ & (new_n25999_ | new_n25910_));
  assign new_n26493_ = (~new_n26046_ & new_n26157_) | (~new_n25542_ & (~new_n26046_ | new_n26157_));
  assign new_n26494_ = new_n26495_ ? (~new_n26505_ ^ new_n26506_) : (new_n26505_ ^ new_n26506_);
  assign new_n26495_ = new_n26496_ ? (~new_n26503_ ^ new_n26504_) : (new_n26503_ ^ new_n26504_);
  assign new_n26496_ = new_n26497_ ? (~new_n26498_ ^ new_n26502_) : (new_n26498_ ^ new_n26502_);
  assign new_n26497_ = (new_n26057_ & new_n26076_) | (new_n26049_ & (new_n26057_ | new_n26076_));
  assign new_n26498_ = new_n26499_ ? (new_n26500_ ^ new_n26501_) : (~new_n26500_ ^ new_n26501_);
  assign new_n26499_ = ~new_n26075_ & new_n26058_;
  assign new_n26500_ = new_n26219_ & new_n26234_;
  assign new_n26501_ = new_n26083_ & new_n26127_;
  assign new_n26502_ = (new_n26218_ & new_n26236_) | (new_n26208_ & (new_n26218_ | new_n26236_));
  assign new_n26503_ = (new_n26237_ & new_n26150_) | (~new_n26207_ & (new_n26237_ | new_n26150_));
  assign new_n26504_ = new_n26238_ & new_n26247_;
  assign new_n26505_ = (new_n26045_ & new_n26156_) | (~new_n26047_ & (new_n26045_ | new_n26156_));
  assign new_n26506_ = (new_n26157_ & new_n26250_) | (~new_n26206_ & (new_n26157_ | new_n26250_));
  assign new_n26507_ = (~new_n26204_ & new_n26291_) | (~new_n25541_ & (~new_n26204_ | new_n26291_));
  assign new_n26508_ = (new_n26257_ & new_n26277_) | (~new_n26205_ & (new_n26257_ | new_n26277_));
  assign new_n26509_ = (new_n26292_ & new_n26305_) | (~new_n25540_ & (new_n26292_ | new_n26305_));
  assign new_n26510_ = new_n26000_ & new_n26043_;
  assign new_n26511_ = (new_n26368_ & new_n26386_) | (~new_n25539_ & (new_n26368_ | new_n26386_));
  assign \o[51]  = ~new_n26513_ ^ new_n26514_;
  assign new_n26513_ = (~new_n26452_ & new_n26511_) | (new_n26451_ & (~new_n26452_ | new_n26511_));
  assign new_n26514_ = new_n26515_ ^ new_n26516_;
  assign new_n26515_ = (new_n26509_ & new_n26510_) | (~new_n26453_ & (new_n26509_ | new_n26510_));
  assign new_n26516_ = ~new_n26517_ ^ new_n26518_;
  assign new_n26517_ = (new_n26507_ & new_n26508_) | (~new_n26454_ & (new_n26507_ | new_n26508_));
  assign new_n26518_ = new_n26519_ ? (new_n26520_ ^ new_n26547_) : (~new_n26520_ ^ new_n26547_);
  assign new_n26519_ = (~new_n26494_ & new_n26493_) | (~new_n26455_ & (~new_n26494_ | new_n26493_));
  assign new_n26520_ = new_n26521_ ? (new_n26522_ ^ new_n26539_) : (~new_n26522_ ^ new_n26539_);
  assign new_n26521_ = (~new_n26480_ & new_n26479_) | (~new_n26456_ & (~new_n26480_ | new_n26479_));
  assign new_n26522_ = new_n26523_ ? (new_n26527_ ^ new_n26528_) : (~new_n26527_ ^ new_n26528_);
  assign new_n26523_ = new_n26524_ ? (new_n26525_ ^ new_n26526_) : (~new_n26525_ ^ new_n26526_);
  assign new_n26524_ = (new_n26464_ & new_n26465_) | (~new_n26458_ & (new_n26464_ | new_n26465_));
  assign new_n26525_ = (~new_n26487_ & new_n26491_) | (~new_n26483_ & (~new_n26487_ | new_n26491_));
  assign new_n26526_ = (new_n26485_ & new_n26486_) | (new_n26484_ & (new_n26485_ | new_n26486_));
  assign new_n26527_ = (~new_n26466_ & new_n26478_) | (~new_n26457_ & (~new_n26466_ | new_n26478_));
  assign new_n26528_ = new_n26529_ ? (new_n26532_ ^ new_n26538_) : (~new_n26532_ ^ new_n26538_);
  assign new_n26529_ = ~new_n26530_ ^ new_n26531_;
  assign new_n26530_ = (new_n26462_ & new_n26463_) | (new_n26459_ & (new_n26462_ | new_n26463_));
  assign new_n26531_ = (new_n26469_ & new_n26470_) | (new_n26468_ & (new_n26469_ | new_n26470_));
  assign new_n26532_ = new_n26533_ ^ new_n26537_;
  assign new_n26533_ = new_n26534_ ? (new_n26535_ ^ new_n26536_) : (~new_n26535_ ^ new_n26536_);
  assign new_n26534_ = new_n26460_ & new_n26461_;
  assign new_n26535_ = new_n25624_ & new_n25546_ & new_n25623_;
  assign new_n26536_ = new_n26476_ & new_n26477_;
  assign new_n26537_ = (new_n26474_ & new_n26475_) | (new_n26473_ & (new_n26474_ | new_n26475_));
  assign new_n26538_ = (~new_n26472_ & new_n26471_) | (~new_n26467_ & (~new_n26472_ | new_n26471_));
  assign new_n26539_ = new_n26540_ ? (~new_n26541_ ^ new_n26546_) : (new_n26541_ ^ new_n26546_);
  assign new_n26540_ = (new_n26503_ & new_n26504_) | (~new_n26496_ & (new_n26503_ | new_n26504_));
  assign new_n26541_ = ~new_n26542_ ^ new_n26543_;
  assign new_n26542_ = (~new_n26498_ & new_n26502_) | (new_n26497_ & (~new_n26498_ | new_n26502_));
  assign new_n26543_ = new_n26544_ ^ new_n26545_;
  assign new_n26544_ = (new_n26500_ & new_n26501_) | (new_n26499_ & (new_n26500_ | new_n26501_));
  assign new_n26545_ = (new_n26489_ & new_n26490_) | (new_n26488_ & (new_n26489_ | new_n26490_));
  assign new_n26546_ = (~new_n26482_ & new_n26492_) | (new_n26481_ & (~new_n26482_ | new_n26492_));
  assign new_n26547_ = (new_n26505_ & new_n26506_) | (~new_n26495_ & (new_n26505_ | new_n26506_));
  assign \o[52]  = ((new_n26549_ | new_n26550_) & (new_n26551_ ^ new_n26552_)) | (~new_n26549_ & ~new_n26550_ & (~new_n26551_ ^ new_n26552_));
  assign new_n26549_ = ~new_n26514_ & new_n26513_;
  assign new_n26550_ = ~new_n26516_ & new_n26515_;
  assign new_n26551_ = new_n26517_ & new_n26518_;
  assign new_n26552_ = ~new_n26553_ ^ new_n26554_;
  assign new_n26553_ = (~new_n26520_ & new_n26547_) | (new_n26519_ & (~new_n26520_ | new_n26547_));
  assign new_n26554_ = new_n26555_ ? (new_n26556_ ^ new_n26568_) : (~new_n26556_ ^ new_n26568_);
  assign new_n26555_ = (~new_n26522_ & ~new_n26539_) | (new_n26521_ & (~new_n26522_ | ~new_n26539_));
  assign new_n26556_ = new_n26557_ ? (new_n26561_ ^ new_n26562_) : (~new_n26561_ ^ new_n26562_);
  assign new_n26557_ = new_n26558_ ? (new_n26559_ ^ new_n26560_) : (~new_n26559_ ^ new_n26560_);
  assign new_n26558_ = (new_n26525_ & new_n26526_) | (new_n26524_ & (new_n26525_ | new_n26526_));
  assign new_n26559_ = new_n26542_ & new_n26543_;
  assign new_n26560_ = new_n26544_ & new_n26545_;
  assign new_n26561_ = (~new_n26528_ & new_n26527_) | (~new_n26523_ & (~new_n26528_ | new_n26527_));
  assign new_n26562_ = new_n26563_ ? (~new_n26564_ ^ new_n26567_) : (new_n26564_ ^ new_n26567_);
  assign new_n26563_ = (~new_n26532_ & new_n26538_) | (~new_n26529_ & (~new_n26532_ | new_n26538_));
  assign new_n26564_ = ~new_n26565_ ^ new_n26566_;
  assign new_n26565_ = ~new_n26533_ & new_n26537_;
  assign new_n26566_ = (new_n26535_ & new_n26536_) | (new_n26534_ & (new_n26535_ | new_n26536_));
  assign new_n26567_ = new_n26530_ & new_n26531_;
  assign new_n26568_ = (~new_n26541_ & new_n26546_) | (new_n26540_ & (~new_n26541_ | new_n26546_));
  assign \o[53]  = ~new_n26570_ ^ new_n26571_;
  assign new_n26570_ = (new_n26551_ | (~new_n26552_ & (new_n26550_ | new_n26549_))) & (new_n26550_ | new_n26549_ | ~new_n26552_);
  assign new_n26571_ = new_n26572_ ^ new_n26573_;
  assign new_n26572_ = new_n26553_ & new_n26554_;
  assign new_n26573_ = ~new_n26574_ ^ new_n26575_;
  assign new_n26574_ = (~new_n26556_ & new_n26568_) | (new_n26555_ & (~new_n26556_ | new_n26568_));
  assign new_n26575_ = new_n26576_ ? (new_n26577_ ^ new_n26580_) : (~new_n26577_ ^ new_n26580_);
  assign new_n26576_ = (~new_n26562_ & new_n26561_) | (~new_n26557_ & (~new_n26562_ | new_n26561_));
  assign new_n26577_ = ~new_n26578_ ^ new_n26579_;
  assign new_n26578_ = (~new_n26564_ & new_n26567_) | (new_n26563_ & (~new_n26564_ | new_n26567_));
  assign new_n26579_ = new_n26565_ & new_n26566_;
  assign new_n26580_ = (new_n26559_ & new_n26560_) | (new_n26558_ & (new_n26559_ | new_n26560_));
  assign \o[54]  = ((new_n26585_ ^ new_n26586_) & ((~new_n26582_ & ~new_n26583_ & ~new_n26584_) | (new_n26584_ & (new_n26582_ | new_n26583_)))) | (((~new_n26584_ & (new_n26582_ | new_n26583_)) | (~new_n26582_ & ~new_n26583_ & new_n26584_)) & (new_n26585_ ^ ~new_n26586_));
  assign new_n26582_ = ~new_n26571_ & new_n26570_;
  assign new_n26583_ = ~new_n26573_ & new_n26572_;
  assign new_n26584_ = new_n26574_ & new_n26575_;
  assign new_n26585_ = (~new_n26577_ & new_n26580_) | (new_n26576_ & (~new_n26577_ | new_n26580_));
  assign new_n26586_ = new_n26578_ & new_n26579_;
  assign \o[55]  = (~new_n26584_ | ~new_n26585_ | ~new_n26586_ | (~new_n26582_ & ~new_n26583_)) & (new_n26584_ | new_n26585_ | new_n26586_) & (new_n26582_ | new_n26583_ | ((new_n26585_ | new_n26586_) & (new_n26584_ | (new_n26585_ & new_n26586_))));
  assign \o[56]  = new_n26589_ ? (new_n27000_ ^ new_n27020_) : (~new_n27000_ ^ new_n27020_);
  assign new_n26589_ = new_n26590_ ? (~new_n26957_ ^ new_n26979_) : (new_n26957_ ^ new_n26979_);
  assign new_n26590_ = new_n26591_ ? (new_n26880_ ^ new_n26940_) : (~new_n26880_ ^ new_n26940_);
  assign new_n26591_ = new_n26592_ ? (new_n26694_ ^ new_n26861_) : (~new_n26694_ ^ new_n26861_);
  assign new_n26592_ = new_n26593_ ? (new_n26681_ ^ new_n26693_) : (~new_n26681_ ^ new_n26693_);
  assign new_n26593_ = new_n26594_ ? (new_n26631_ ^ new_n26680_) : (~new_n26631_ ^ new_n26680_);
  assign new_n26594_ = new_n26595_ ? (new_n26614_ ^ new_n26620_) : (~new_n26614_ ^ new_n26620_);
  assign new_n26595_ = ~new_n26596_ & new_n26612_;
  assign new_n26596_ = new_n26610_ & new_n26598_ & (~new_n26611_ | new_n26597_);
  assign new_n26597_ = new_n16278_ ? new_n20441_ : new_n15143_;
  assign new_n26598_ = (~new_n24023_ | ~new_n26603_) & (~new_n26606_ | ~new_n26608_) & (new_n26609_ | ~new_n26599_);
  assign new_n26599_ = ~new_n10242_ & new_n26600_;
  assign new_n26600_ = ~new_n26601_ & ~new_n26602_;
  assign new_n26601_ = ~new_n6734_ & (~new_n6732_ | ~new_n15166_);
  assign new_n26602_ = new_n9935_ & new_n9932_;
  assign new_n26603_ = new_n26604_ & new_n10645_;
  assign new_n26604_ = ~new_n26605_ & new_n26601_;
  assign new_n26605_ = ~new_n6737_ & ~new_n6766_;
  assign new_n26606_ = new_n22283_ ? new_n7374_ : ~new_n26607_;
  assign new_n26607_ = new_n24388_ & new_n18581_;
  assign new_n26608_ = new_n26601_ & new_n26605_;
  assign new_n26609_ = ~new_n24035_ & new_n22419_;
  assign new_n26610_ = (~new_n10242_ | ~new_n26600_) & (new_n10645_ | new_n13850_ | ~new_n26604_);
  assign new_n26611_ = ~new_n26601_ & new_n26602_;
  assign new_n26612_ = new_n26613_ & (new_n26606_ | ~new_n26608_) & (~new_n26611_ | ~new_n26597_);
  assign new_n26613_ = (new_n24023_ | ~new_n26603_) & (~new_n26599_ | ~new_n26609_);
  assign new_n26614_ = ~new_n26616_ & ~new_n26618_ & (new_n26617_ | (new_n26615_ & ~new_n16192_) | (new_n26619_ & new_n16192_));
  assign new_n26615_ = new_n16956_ ? ~new_n25903_ : ~new_n17898_;
  assign new_n26616_ = new_n26617_ & new_n18385_ & (new_n24905_ ? new_n8985_ : new_n8200_);
  assign new_n26617_ = new_n25920_ & new_n8915_;
  assign new_n26618_ = ~new_n18385_ & new_n18887_ & new_n26617_ & new_n6841_ & (new_n6838_ | new_n6805_);
  assign new_n26619_ = ~new_n8133_ & (new_n20447_ | ~new_n18961_);
  assign new_n26620_ = ~new_n26625_ & new_n26627_ & (new_n10539_ | (new_n26621_ & ~new_n26630_) | (new_n26623_ & new_n26630_));
  assign new_n26621_ = (new_n26622_ & new_n8292_ & (new_n16411_ | new_n8269_)) | (~new_n25934_ & new_n25771_ & (~new_n8292_ | (~new_n16411_ & ~new_n8269_)));
  assign new_n26622_ = ~new_n14913_ & (~new_n14906_ | ~new_n14885_ | ~new_n14915_);
  assign new_n26623_ = (new_n26624_ & (new_n16101_ | new_n16098_)) | (new_n17330_ & new_n17357_ & ~new_n26624_);
  assign new_n26624_ = ~new_n12354_ & (~new_n14164_ | new_n14172_);
  assign new_n26625_ = ~new_n9457_ & new_n10539_ & (new_n15716_ ? new_n10936_ : (new_n19125_ | new_n26626_));
  assign new_n26626_ = new_n19127_ & (new_n19118_ | new_n19097_);
  assign new_n26627_ = ~new_n9457_ | ~new_n10539_ | ((new_n26629_ | ~new_n26628_) & (new_n23081_ | ~new_n21487_ | new_n26628_));
  assign new_n26628_ = ~new_n10526_ & new_n9583_;
  assign new_n26629_ = ~new_n19592_ & new_n18705_;
  assign new_n26630_ = ~new_n15788_ & new_n23964_;
  assign new_n26631_ = new_n26632_ ? (new_n26657_ ^ new_n26672_) : (~new_n26657_ ^ new_n26672_);
  assign new_n26632_ = ~new_n26633_ & new_n26654_;
  assign new_n26633_ = ~new_n26650_ & new_n26634_ & (~new_n26651_ | (new_n24023_ & new_n26653_) | (new_n26652_ & ~new_n26653_));
  assign new_n26634_ = ~new_n26635_ & (~new_n26640_ | (~new_n26641_ & new_n26648_) | (~new_n26649_ & ~new_n26648_));
  assign new_n26635_ = new_n26636_ & ((new_n26638_ & new_n13014_ & new_n8703_) | (~new_n26639_ & new_n24007_ & ~new_n8703_));
  assign new_n26636_ = new_n12537_ & new_n26637_;
  assign new_n26637_ = ~new_n24186_ & ~new_n24190_;
  assign new_n26638_ = ~new_n25924_ & new_n6908_;
  assign new_n26639_ = new_n26274_ & new_n8128_;
  assign new_n26640_ = ~new_n16749_ & ~new_n26636_;
  assign new_n26641_ = new_n20405_ & (new_n20402_ | new_n26642_);
  assign new_n26642_ = new_n26643_ & new_n20377_;
  assign new_n26643_ = (new_n26644_ | (new_n20401_ & (~\all_features[1851]  | ~\all_features[1852]  | (~\all_features[1850]  & new_n20381_)))) & (~new_n20401_ | \all_features[1851]  | \all_features[1852] );
  assign new_n26644_ = ~new_n20390_ & (new_n20389_ | (~new_n20393_ & (new_n20395_ | (~new_n26645_ & ~new_n20398_))));
  assign new_n26645_ = ~new_n20397_ & (~\all_features[1855]  | new_n26646_ | (~\all_features[1852]  & ~\all_features[1853]  & ~\all_features[1854] ));
  assign new_n26646_ = \all_features[1855]  & ((~new_n26647_ & ~\all_features[1853]  & \all_features[1854] ) | (~new_n20383_ & (\all_features[1854]  | (~new_n20380_ & \all_features[1853] ))));
  assign new_n26647_ = (\all_features[1852]  & (\all_features[1850]  | \all_features[1851] )) | (~new_n20386_ & ~\all_features[1850]  & ~\all_features[1851]  & ~\all_features[1852] );
  assign new_n26648_ = ~new_n9234_ & (~new_n9211_ | new_n9236_);
  assign new_n26649_ = new_n20086_ & new_n22838_;
  assign new_n26650_ = new_n26636_ & (new_n8703_ ? ~new_n13014_ : ~new_n24007_);
  assign new_n26651_ = ~new_n26636_ & new_n16749_;
  assign new_n26652_ = ~new_n19083_ & (~new_n19060_ | new_n25958_);
  assign new_n26653_ = ~new_n9930_ & ~new_n9932_;
  assign new_n26654_ = new_n26655_ & (new_n26653_ | ~new_n26652_ | ~new_n26651_);
  assign new_n26655_ = new_n26656_ & (~new_n26640_ | (new_n26641_ & new_n26648_) | (new_n26649_ & ~new_n26648_));
  assign new_n26656_ = ~new_n26636_ | ((new_n26638_ | ~new_n13014_ | ~new_n8703_) & (~new_n26639_ | ~new_n24007_ | new_n8703_));
  assign new_n26657_ = ~new_n26658_ & new_n26669_;
  assign new_n26658_ = new_n26659_ & new_n26666_;
  assign new_n26659_ = (~new_n26664_ | new_n26665_) & (~new_n26660_ | (new_n26663_ ? ~new_n22546_ : new_n14436_));
  assign new_n26660_ = new_n26661_ & new_n26662_;
  assign new_n26661_ = new_n10310_ & (~new_n10339_ | ~new_n10335_);
  assign new_n26662_ = new_n20201_ & new_n20173_ & new_n20194_;
  assign new_n26663_ = new_n10168_ & new_n13098_;
  assign new_n26664_ = ~new_n26662_ & new_n26661_;
  assign new_n26665_ = new_n18578_ & new_n25366_;
  assign new_n26666_ = new_n26661_ | (new_n20845_ ? (new_n11171_ ? ~new_n26668_ : new_n26232_) : ~new_n26667_);
  assign new_n26667_ = (~new_n19821_ & new_n16946_) | (new_n9999_ & new_n7501_ & ~new_n16946_);
  assign new_n26668_ = ~new_n16759_ & new_n10833_;
  assign new_n26669_ = new_n26670_ & (new_n26661_ | ((~new_n26671_ | ~new_n20845_) & (~new_n16946_ | ~new_n19821_ | new_n20845_)));
  assign new_n26670_ = (~new_n26665_ | ~new_n26664_) & (~new_n26660_ | (new_n26663_ ? new_n22546_ : ~new_n14436_));
  assign new_n26671_ = new_n11171_ ? ~new_n26668_ : new_n26232_;
  assign new_n26672_ = new_n26673_ & (~new_n15494_ | ~new_n14469_ | new_n25035_ | new_n26676_);
  assign new_n26673_ = ~new_n26674_ & (~new_n26679_ | ~new_n26676_ | new_n26677_ | new_n26678_);
  assign new_n26674_ = new_n21616_ & new_n26675_ & ~new_n14469_ & ~new_n26676_;
  assign new_n26675_ = ~new_n14422_ & new_n14393_;
  assign new_n26676_ = new_n9411_ & (new_n9414_ | new_n9418_ | new_n9389_);
  assign new_n26677_ = new_n16263_ & (new_n16261_ | ~new_n18386_);
  assign new_n26678_ = new_n17802_ & (new_n17800_ | ~new_n18043_);
  assign new_n26679_ = new_n16334_ & new_n10637_;
  assign new_n26680_ = new_n26633_ & new_n26654_;
  assign new_n26681_ = ~new_n26682_ & new_n26691_;
  assign new_n26682_ = new_n26683_ & (~new_n23666_ | (~new_n26688_ & new_n26690_) | (new_n26689_ & ~new_n26690_));
  assign new_n26683_ = new_n23666_ | (~new_n21527_ & new_n22932_ & ~new_n17709_) | (new_n26684_ & new_n17709_);
  assign new_n26684_ = new_n26687_ ? new_n26685_ : new_n26686_;
  assign new_n26685_ = ~new_n8544_ & ~new_n6955_;
  assign new_n26686_ = ~new_n7367_ & new_n7340_;
  assign new_n26687_ = new_n18444_ & (new_n18451_ | new_n18422_);
  assign new_n26688_ = (~new_n22998_ & ~new_n21529_) | (new_n23737_ & new_n25359_ & new_n21529_);
  assign new_n26689_ = new_n9457_ & new_n12560_ & (new_n12538_ | ~new_n26637_);
  assign new_n26690_ = new_n9996_ & new_n16348_;
  assign new_n26691_ = (new_n26692_ | ~new_n17709_ | new_n23666_) & (~new_n23666_ | (new_n26690_ ? new_n26688_ : ~new_n26689_));
  assign new_n26692_ = new_n26687_ ? ~new_n26685_ : ~new_n26686_;
  assign new_n26693_ = new_n16890_ & ~new_n22389_ & new_n16887_;
  assign new_n26694_ = new_n26695_ ? (new_n26736_ ^ new_n26854_) : (~new_n26736_ ^ new_n26854_);
  assign new_n26695_ = new_n26696_ ? (~new_n26726_ ^ new_n26727_) : (new_n26726_ ^ new_n26727_);
  assign new_n26696_ = new_n26697_ ? (new_n26711_ ^ new_n26720_) : (~new_n26711_ ^ new_n26720_);
  assign new_n26697_ = ~new_n26698_ & new_n26708_;
  assign new_n26698_ = new_n26699_ & (~new_n26701_ | ((new_n26706_ | new_n26707_ | ~new_n24452_) & (new_n18754_ | new_n24452_)));
  assign new_n26699_ = (~new_n26700_ | new_n26705_) & (new_n26701_ | (new_n10241_ ? new_n26704_ : ~new_n26702_));
  assign new_n26700_ = new_n26701_ & ~new_n24452_ & new_n18754_;
  assign new_n26701_ = ~new_n12490_ & (~new_n12487_ | new_n15714_);
  assign new_n26702_ = new_n26703_ ? ~new_n12117_ : ~new_n7635_;
  assign new_n26703_ = new_n22083_ & (new_n22080_ | new_n22053_);
  assign new_n26704_ = new_n9725_ & (new_n25032_ | ~new_n23834_);
  assign new_n26705_ = ~new_n9544_ & new_n9518_;
  assign new_n26706_ = ~new_n26389_ & ~new_n12115_;
  assign new_n26707_ = ~new_n17320_ & ~new_n17322_ & (~new_n17313_ | ~new_n17292_);
  assign new_n26708_ = new_n26709_ & (new_n10241_ | new_n26701_ | (new_n26703_ ? ~new_n12117_ : ~new_n7635_));
  assign new_n26709_ = (~new_n26705_ | ~new_n26700_) & (~new_n26710_ | (new_n26706_ ? new_n19889_ : ~new_n26707_));
  assign new_n26710_ = new_n26701_ & new_n24452_;
  assign new_n26711_ = new_n26712_ & (new_n21250_ ? new_n26719_ : new_n26717_);
  assign new_n26712_ = new_n26713_ & (~new_n26716_ | ~new_n20483_ | ~new_n19717_ | ~new_n21250_);
  assign new_n26713_ = (~new_n26715_ | new_n26714_ | ~new_n21250_) & (new_n22048_ | new_n26607_ | ~new_n19244_ | new_n21250_);
  assign new_n26714_ = ~new_n23063_ & new_n7863_;
  assign new_n26715_ = ~new_n7866_ & ~new_n7942_ & ~new_n20483_;
  assign new_n26716_ = ~new_n10024_ & (~new_n10002_ | ~new_n16345_);
  assign new_n26717_ = (~new_n26718_ | ~new_n26607_) & (new_n25415_ | ~new_n22048_ | ~new_n24565_ | new_n26607_);
  assign new_n26718_ = new_n24496_ & new_n17152_ & new_n25409_;
  assign new_n26719_ = (new_n26716_ | ~new_n19773_ | ~new_n20483_) & (~new_n20262_ | ~new_n7942_ | new_n20483_);
  assign new_n26720_ = new_n26721_ & (new_n26722_ | ((new_n26724_ | ~new_n6354_) & (~new_n16946_ | ~new_n20589_ | new_n6354_)));
  assign new_n26721_ = ~new_n26722_ | ((~new_n15592_ | ~new_n22036_ | new_n16376_) & (~new_n16376_ | (new_n26723_ & ~new_n15588_)));
  assign new_n26722_ = new_n22276_ & new_n8854_;
  assign new_n26723_ = ~new_n22608_ & new_n6662_;
  assign new_n26724_ = (~new_n25663_ & ~new_n8132_) ? (new_n12141_ | ~new_n24346_) : new_n26725_;
  assign new_n26725_ = new_n6566_ & (new_n6563_ | new_n6556_);
  assign new_n26726_ = new_n26596_ & new_n26612_;
  assign new_n26727_ = new_n26734_ & (new_n25957_ ? new_n26731_ : new_n26728_);
  assign new_n26728_ = (new_n20048_ | ~new_n26729_ | ~new_n26134_) & (~new_n20582_ | ~new_n26730_ | new_n26134_);
  assign new_n26729_ = ~new_n8879_ & (~new_n8885_ | ~new_n8857_);
  assign new_n26730_ = ~new_n19017_ & (~new_n18991_ | ~new_n19018_);
  assign new_n26731_ = (~new_n11373_ | new_n26732_ | ~new_n12737_) & (new_n26733_ | new_n19813_ | ~new_n14690_ | new_n12737_);
  assign new_n26732_ = new_n7772_ & new_n7798_;
  assign new_n26733_ = new_n19802_ & new_n19811_;
  assign new_n26734_ = (~new_n26735_ | new_n26266_ | ~new_n25957_) & (new_n26729_ | ~new_n14336_ | ~new_n26134_ | new_n25957_);
  assign new_n26735_ = new_n12737_ & new_n26732_;
  assign new_n26736_ = new_n26737_ ? (new_n26786_ ^ new_n26726_) : (~new_n26786_ ^ new_n26726_);
  assign new_n26737_ = new_n26738_ ? (new_n26752_ ^ new_n26771_) : (~new_n26752_ ^ new_n26771_);
  assign new_n26738_ = ~new_n26739_ & new_n26750_;
  assign new_n26739_ = new_n26740_ & (new_n26749_ | ~new_n26745_ | ~new_n26746_ | (~new_n20262_ & ~new_n12562_));
  assign new_n26740_ = (new_n26746_ | new_n26747_ | ~new_n26745_) & (new_n26745_ | (new_n26748_ ? new_n26743_ : ~new_n26741_));
  assign new_n26741_ = new_n14159_ & ~new_n21602_ & new_n26742_;
  assign new_n26742_ = new_n24009_ & (~new_n25937_ | ~new_n24019_);
  assign new_n26743_ = new_n23926_ ? new_n26744_ : ~new_n24185_;
  assign new_n26744_ = ~new_n21793_ & new_n21800_;
  assign new_n26745_ = ~new_n17612_ & new_n24118_;
  assign new_n26746_ = new_n10282_ & new_n24156_;
  assign new_n26747_ = new_n9749_ & new_n9727_ & ~new_n9750_ & new_n18581_;
  assign new_n26748_ = ~new_n11672_ & (~new_n11669_ | ~new_n11658_);
  assign new_n26749_ = new_n12562_ & ~new_n23190_ & new_n8742_;
  assign new_n26750_ = new_n26751_ & (new_n26745_ | ~new_n26748_ | (new_n23926_ ? ~new_n26744_ : new_n24185_));
  assign new_n26751_ = (new_n26748_ | new_n26741_ | new_n26745_) & (~new_n26745_ | (new_n26746_ ? ~new_n26749_ : ~new_n26747_));
  assign new_n26752_ = ~new_n26769_ & new_n26753_;
  assign new_n26753_ = ~new_n26763_ & new_n26754_ & (new_n23649_ ? (new_n11622_ | ~new_n26766_) : new_n26767_);
  assign new_n26754_ = (new_n26755_ | ~new_n11622_ | ~new_n23649_) & (~new_n26762_ | ~new_n26761_);
  assign new_n26755_ = ~new_n26756_ & (new_n19017_ | new_n26757_);
  assign new_n26756_ = ~new_n6424_ & (~new_n6421_ | new_n6390_);
  assign new_n26757_ = new_n18991_ & (new_n19018_ | (~new_n19011_ & (new_n19010_ | (~new_n26758_ & ~new_n19006_))));
  assign new_n26758_ = ~new_n19008_ & (new_n19001_ | (~new_n19002_ & (new_n18994_ | new_n26759_)));
  assign new_n26759_ = ~new_n18996_ & (~new_n19016_ | (new_n19015_ & (~new_n19012_ | (~new_n26760_ & new_n19013_))));
  assign new_n26760_ = \all_features[2526]  & \all_features[2527]  & (\all_features[2525]  | (~new_n19014_ & \all_features[2524] ));
  assign new_n26761_ = new_n24200_ & ~new_n23217_ & ~new_n23649_;
  assign new_n26762_ = ~new_n7089_ & new_n7097_;
  assign new_n26763_ = new_n26764_ & new_n26765_;
  assign new_n26764_ = new_n23217_ & ~new_n11337_ & ~new_n23649_;
  assign new_n26765_ = new_n14784_ & new_n25362_;
  assign new_n26766_ = new_n18578_ & new_n24514_;
  assign new_n26767_ = (~new_n11337_ | ~new_n24564_ | ~new_n23217_) & (new_n24200_ | new_n26768_ | new_n23217_);
  assign new_n26768_ = ~new_n22689_ & ~new_n22685_ & ~new_n22658_;
  assign new_n26769_ = new_n26770_ & (~new_n23649_ | (~new_n26755_ & new_n11622_) | (new_n26766_ & ~new_n11622_));
  assign new_n26770_ = (new_n26765_ | ~new_n26764_) & (new_n26762_ | ~new_n26761_);
  assign new_n26771_ = ~new_n26772_ & new_n26783_;
  assign new_n26772_ = new_n26773_ & (new_n25077_ ? (new_n26607_ | (new_n22283_ & new_n26782_) | (~new_n22283_ & ~new_n26782_)) : new_n26780_);
  assign new_n26773_ = ~new_n26774_ & (~new_n25077_ | ~new_n26607_ | (new_n26779_ ? ~new_n9514_ : ~new_n26778_));
  assign new_n26774_ = new_n26776_ & new_n26775_ & ~new_n26777_ & ~new_n25077_;
  assign new_n26775_ = new_n22553_ & new_n25229_;
  assign new_n26776_ = new_n23823_ & new_n23584_;
  assign new_n26777_ = ~new_n12410_ & new_n15330_;
  assign new_n26778_ = ~new_n12624_ & (~new_n12601_ | ~new_n18164_);
  assign new_n26779_ = ~new_n19027_ & new_n18912_;
  assign new_n26780_ = (new_n26776_ | ~new_n26775_) & (~new_n26781_ | new_n26775_ | (new_n22610_ & (~new_n22635_ | ~new_n22639_)));
  assign new_n26781_ = new_n16023_ & new_n26165_ & new_n15993_;
  assign new_n26782_ = new_n19059_ & new_n25958_;
  assign new_n26783_ = new_n26785_ & ((~new_n26607_ & (new_n22283_ ^ new_n26782_)) | ~new_n25077_ | (new_n26784_ & new_n26607_));
  assign new_n26784_ = new_n26779_ ? new_n9514_ : new_n26778_;
  assign new_n26785_ = new_n25077_ | ((new_n26781_ | new_n26775_) & (~new_n26776_ | ~new_n26777_ | ~new_n26775_));
  assign new_n26786_ = new_n26787_ ^ new_n26840_;
  assign new_n26787_ = new_n26788_ & (~new_n26833_ | (new_n26836_ & (new_n26839_ | ~new_n26837_)));
  assign new_n26788_ = new_n26789_ & (~new_n26831_ | (~new_n18576_ & new_n26832_));
  assign new_n26789_ = new_n26790_ & (~new_n26795_ | ~new_n26797_) & (~new_n26793_ | new_n25377_);
  assign new_n26790_ = ~new_n26791_ | (new_n17936_ ? ~new_n23700_ : ~new_n18892_);
  assign new_n26791_ = ~new_n14084_ & ~new_n26792_;
  assign new_n26792_ = ~new_n20234_ & new_n20535_;
  assign new_n26793_ = ~new_n22710_ & new_n26794_;
  assign new_n26794_ = new_n23598_ & new_n26792_;
  assign new_n26795_ = new_n26796_ & new_n19885_;
  assign new_n26796_ = ~new_n23598_ & new_n26792_;
  assign new_n26797_ = new_n26821_ & (new_n26827_ | (~new_n26828_ & new_n26798_));
  assign new_n26798_ = ~new_n26817_ & ~new_n26819_ & ~new_n26820_ & (new_n26816_ | new_n26815_ | new_n26799_);
  assign new_n26799_ = ~new_n26809_ & ~new_n26811_ & (~new_n26814_ | ~new_n26813_ | new_n26800_);
  assign new_n26800_ = new_n26801_ & ~new_n26807_ & new_n26803_;
  assign new_n26801_ = \all_features[2207]  & (\all_features[2206]  | (new_n26802_ & (\all_features[2202]  | \all_features[2203]  | \all_features[2201] )));
  assign new_n26802_ = \all_features[2204]  & \all_features[2205] ;
  assign new_n26803_ = new_n26806_ & (new_n26804_ | \all_features[2204]  | \all_features[2205]  | ~new_n26805_);
  assign new_n26804_ = \all_features[2200]  & \all_features[2201] ;
  assign new_n26805_ = ~\all_features[2202]  & ~\all_features[2203] ;
  assign new_n26806_ = \all_features[2206]  & \all_features[2207] ;
  assign new_n26807_ = new_n26806_ & \all_features[2205]  & ((~new_n26808_ & \all_features[2202] ) | \all_features[2204]  | \all_features[2203] );
  assign new_n26808_ = ~\all_features[2200]  & ~\all_features[2201] ;
  assign new_n26809_ = ~new_n26810_ & ~\all_features[2207] ;
  assign new_n26810_ = \all_features[2205]  & \all_features[2206]  & (\all_features[2204]  | (\all_features[2202]  & \all_features[2203]  & \all_features[2201] ));
  assign new_n26811_ = ~\all_features[2207]  & (~\all_features[2206]  | ~new_n26812_ | ~new_n26804_ | ~new_n26802_);
  assign new_n26812_ = \all_features[2202]  & \all_features[2203] ;
  assign new_n26813_ = \all_features[2207]  & (\all_features[2206]  | (\all_features[2205]  & (\all_features[2204]  | ~new_n26805_ | ~new_n26808_)));
  assign new_n26814_ = \all_features[2207]  & (\all_features[2205]  | \all_features[2206]  | \all_features[2204] );
  assign new_n26815_ = ~\all_features[2207]  & (~\all_features[2206]  | (~\all_features[2204]  & ~\all_features[2205]  & ~new_n26812_));
  assign new_n26816_ = ~\all_features[2207]  & (~\all_features[2206]  | (~\all_features[2205]  & (new_n26808_ | ~\all_features[2204]  | ~new_n26812_)));
  assign new_n26817_ = new_n26818_ & (~\all_features[2205]  | (~\all_features[2204]  & (~\all_features[2203]  | (~\all_features[2202]  & ~\all_features[2201] ))));
  assign new_n26818_ = ~\all_features[2206]  & ~\all_features[2207] ;
  assign new_n26819_ = new_n26818_ & (~\all_features[2203]  | ~new_n26802_ | (~\all_features[2202]  & ~new_n26804_));
  assign new_n26820_ = ~\all_features[2205]  & new_n26818_ & ((~\all_features[2202]  & new_n26808_) | ~\all_features[2204]  | ~\all_features[2203] );
  assign new_n26821_ = new_n26817_ | ~new_n26826_ | ((new_n26824_ | new_n26820_) & (new_n26809_ | ~new_n26822_));
  assign new_n26822_ = new_n26823_ & ~new_n26816_ & ~new_n26820_;
  assign new_n26823_ = ~new_n26815_ & ~new_n26811_;
  assign new_n26824_ = ~new_n26816_ & ~new_n26809_ & new_n26823_ & (~new_n26813_ | ~new_n26825_);
  assign new_n26825_ = new_n26814_ & new_n26801_ & new_n26803_;
  assign new_n26826_ = ~new_n26819_ & ~new_n26827_;
  assign new_n26827_ = ~\all_features[2207]  & ~\all_features[2206]  & ~\all_features[2205]  & ~\all_features[2203]  & ~\all_features[2204] ;
  assign new_n26828_ = ~new_n26815_ & (new_n26816_ | (~new_n26809_ & (new_n26811_ | new_n26829_)));
  assign new_n26829_ = new_n26814_ & (~new_n26813_ | (new_n26801_ & (new_n26830_ | ~new_n26803_)));
  assign new_n26830_ = new_n26806_ & (\all_features[2205]  | (~new_n26805_ & \all_features[2204] ));
  assign new_n26831_ = ~new_n26792_ & new_n14084_;
  assign new_n26832_ = new_n12933_ & (new_n12910_ | ~new_n12935_);
  assign new_n26833_ = new_n26835_ & (~new_n19339_ | ~new_n26834_);
  assign new_n26834_ = new_n26794_ & new_n22710_;
  assign new_n26835_ = (new_n18576_ | ~new_n26831_ | ~new_n26832_) & (new_n23700_ | ~new_n26791_ | ~new_n17936_);
  assign new_n26836_ = (new_n26797_ | ~new_n26795_) & (~new_n26793_ | ~new_n25377_);
  assign new_n26837_ = ~new_n26838_ & (new_n18892_ | new_n17936_ | ~new_n26791_);
  assign new_n26838_ = new_n14038_ & new_n20114_ & ~new_n19885_ & new_n26796_;
  assign new_n26839_ = ~new_n19339_ & new_n26834_;
  assign new_n26840_ = ~new_n26841_ & new_n26850_;
  assign new_n26841_ = ~new_n26847_ & ~new_n26842_ & (~new_n26845_ | (new_n19508_ & new_n26849_) | (~new_n19159_ & ~new_n26849_));
  assign new_n26842_ = ~new_n18576_ & new_n26843_;
  assign new_n26843_ = ~new_n13405_ & new_n26844_;
  assign new_n26844_ = new_n11337_ & new_n12870_;
  assign new_n26845_ = ~new_n12870_ & new_n26846_;
  assign new_n26846_ = ~new_n11672_ & ~new_n11669_ & ~new_n11637_ & ~new_n11658_;
  assign new_n26847_ = ~new_n11337_ & new_n12870_ & (new_n26848_ | new_n10701_);
  assign new_n26848_ = ~new_n11886_ & new_n18752_;
  assign new_n26849_ = new_n23475_ & (~new_n24528_ | ~new_n23451_);
  assign new_n26850_ = ~new_n26852_ & new_n26851_ & (~new_n26853_ | (~new_n23701_ & new_n11614_));
  assign new_n26851_ = (~new_n26845_ | ~new_n19508_ | ~new_n26849_) & (~new_n18576_ | ~new_n26843_);
  assign new_n26852_ = new_n13405_ & new_n26844_ & (~new_n19412_ | (~new_n19383_ & ~new_n19414_));
  assign new_n26853_ = ~new_n12870_ & ~new_n26846_;
  assign new_n26854_ = ~new_n26858_ & ~new_n26860_ & (new_n26859_ ? (new_n15873_ | ~new_n24810_) : new_n26855_);
  assign new_n26855_ = (new_n7444_ | new_n26857_ | new_n6662_ | new_n26856_) & (~new_n21484_ | new_n24892_ | ~new_n26856_);
  assign new_n26856_ = ~new_n11576_ & new_n11904_;
  assign new_n26857_ = new_n14955_ & new_n14985_;
  assign new_n26858_ = new_n15479_ & new_n26856_ & ~new_n21484_ & ~new_n26859_;
  assign new_n26859_ = new_n24110_ & (new_n24107_ | new_n24099_);
  assign new_n26860_ = ~new_n26859_ & ~new_n26856_ & new_n26857_ & new_n18701_ & (~new_n18691_ | ~new_n18671_);
  assign new_n26861_ = ~new_n26877_ & new_n26862_;
  assign new_n26862_ = new_n26863_ & (new_n19506_ | ~new_n26875_) & (~new_n26874_ | ~new_n22365_ | ~new_n26876_);
  assign new_n26863_ = ~new_n26864_ & (~new_n26867_ | (~new_n20489_ & new_n26868_) | (~new_n26873_ & ~new_n26868_));
  assign new_n26864_ = new_n26865_ & (new_n20738_ ? ~new_n25614_ : new_n18751_);
  assign new_n26865_ = ~new_n23556_ & ~new_n26866_;
  assign new_n26866_ = new_n15042_ & new_n24002_;
  assign new_n26867_ = new_n23556_ & new_n23450_;
  assign new_n26868_ = ~new_n26869_ & ~new_n18510_;
  assign new_n26869_ = ~new_n18503_ & new_n18507_ & new_n18481_ & (new_n18502_ | new_n26870_);
  assign new_n26870_ = ~new_n18498_ & (new_n18500_ | (~new_n18494_ & (new_n18496_ | (~new_n26871_ & ~new_n18504_))));
  assign new_n26871_ = ~new_n18506_ & (~new_n18492_ | (new_n18491_ & (~new_n18486_ | (~new_n26872_ & new_n18488_))));
  assign new_n26872_ = \all_features[5102]  & \all_features[5103]  & (\all_features[5101]  | (~new_n18490_ & \all_features[5100] ));
  assign new_n26873_ = ~new_n22893_ & ~new_n19318_;
  assign new_n26874_ = ~new_n23556_ & new_n26866_;
  assign new_n26875_ = ~new_n23450_ & new_n23556_;
  assign new_n26876_ = new_n25207_ & new_n20957_;
  assign new_n26877_ = ~new_n26878_ & new_n26879_ & (~new_n26867_ | (new_n20489_ & new_n26868_) | (new_n26873_ & ~new_n26868_));
  assign new_n26878_ = new_n26865_ & (new_n20738_ ? new_n25614_ : ~new_n18751_);
  assign new_n26879_ = (~new_n26875_ | ~new_n19506_ | ~new_n26765_) & (~new_n26874_ | (new_n26876_ & new_n22365_));
  assign new_n26880_ = new_n26881_ ? (~new_n26906_ ^ new_n26924_) : (new_n26906_ ^ new_n26924_);
  assign new_n26881_ = new_n26680_ ? (~new_n26882_ ^ new_n26898_) : (new_n26882_ ^ new_n26898_);
  assign new_n26882_ = new_n26883_ ? (new_n26888_ ^ new_n26893_) : (~new_n26888_ ^ new_n26893_);
  assign new_n26883_ = new_n26886_ & ((~new_n12409_ & new_n18039_ & (new_n6734_ | new_n26885_)) | (~new_n26884_ & (new_n12409_ | ~new_n18039_)));
  assign new_n26884_ = new_n25549_ & ~new_n6734_ & new_n11897_;
  assign new_n26885_ = (new_n20043_ & new_n25804_) ? (~new_n8890_ | ~new_n22457_) : ~new_n24452_;
  assign new_n26886_ = (~new_n26887_ | ~new_n22532_) & (new_n9996_ | ~new_n9611_ | ~new_n26388_ | ~new_n6734_ | new_n22532_);
  assign new_n26887_ = ~new_n18444_ & new_n6734_ & new_n13350_ & (~new_n18451_ | ~new_n18422_);
  assign new_n26888_ = ~new_n26889_ & (~new_n26213_ | ((~new_n19433_ | ~new_n20786_ | new_n26892_) & (new_n19773_ | ~new_n26892_)));
  assign new_n26889_ = new_n26890_ & (new_n17675_ ? new_n20155_ : new_n26891_);
  assign new_n26890_ = ~new_n26213_ & ~new_n24784_ & (~new_n25066_ | ~new_n24760_);
  assign new_n26891_ = new_n21856_ & new_n21880_;
  assign new_n26892_ = new_n21804_ & new_n21771_ & new_n21801_;
  assign new_n26893_ = (new_n26897_ | ~new_n20923_ | new_n26756_) & (~new_n26756_ | (~new_n26896_ & (~new_n24512_ | new_n26894_)));
  assign new_n26894_ = new_n12408_ ? new_n11674_ : ~new_n26895_;
  assign new_n26895_ = ~new_n15793_ & new_n23964_;
  assign new_n26896_ = ~new_n24512_ & new_n18420_ & (new_n14374_ | (new_n14352_ & new_n14376_));
  assign new_n26897_ = (new_n12141_ & (~new_n12142_ | new_n12119_)) ? new_n24112_ : new_n23779_;
  assign new_n26898_ = ~new_n26903_ & (new_n12864_ ? (new_n26904_ ? new_n26901_ : new_n26905_) : new_n26899_);
  assign new_n26899_ = (new_n26900_ | ~new_n25277_ | ~new_n21589_) & (new_n15745_ | ~new_n6497_ | new_n21589_);
  assign new_n26900_ = new_n11269_ & ~new_n18903_ & new_n11267_;
  assign new_n26901_ = (~new_n14044_ & new_n7228_ & ~new_n26902_) | (~new_n23781_ & new_n10562_ & (~new_n7228_ | new_n26902_));
  assign new_n26902_ = new_n7257_ & new_n7253_;
  assign new_n26903_ = ~new_n25277_ & ~new_n12864_ & new_n21589_ & (~new_n24008_ | new_n11616_);
  assign new_n26904_ = ~new_n22932_ & (~new_n22934_ | ~new_n22145_);
  assign new_n26905_ = (~new_n22772_ & new_n12525_ & new_n12600_) | (~new_n12600_ & (new_n16058_ | ~new_n25214_));
  assign new_n26906_ = ~new_n26907_ & new_n26922_;
  assign new_n26907_ = ~new_n26919_ & new_n26908_;
  assign new_n26908_ = new_n26914_ & (~new_n26913_ | new_n26917_) & (~new_n26909_ | (~new_n26916_ & ~new_n26918_));
  assign new_n26909_ = new_n26910_ & new_n26912_;
  assign new_n26910_ = ~new_n20925_ & new_n26911_;
  assign new_n26911_ = ~new_n20945_ & new_n24144_;
  assign new_n26912_ = new_n21411_ & new_n22994_;
  assign new_n26913_ = ~new_n26910_ & new_n26912_;
  assign new_n26914_ = new_n26912_ | ((new_n22771_ | ~new_n26607_ | ~new_n26765_) & (~new_n26915_ | new_n26765_));
  assign new_n26915_ = ~new_n18705_ & (~new_n18702_ | new_n18670_);
  assign new_n26916_ = ~new_n26706_ & ~new_n26895_;
  assign new_n26917_ = (~new_n13556_ & (~new_n13545_ | ~new_n13553_)) ? new_n12977_ : new_n17709_;
  assign new_n26918_ = new_n26706_ & new_n23134_;
  assign new_n26919_ = ~new_n26912_ & ((~new_n26915_ & new_n24145_ & ~new_n26765_) | (~new_n26607_ & ~new_n26920_ & new_n26765_));
  assign new_n26920_ = new_n25905_ & new_n26921_;
  assign new_n26921_ = new_n14760_ & new_n14782_;
  assign new_n26922_ = ~new_n26923_ & (~new_n26913_ | ~new_n26917_) & (new_n26916_ | new_n26918_ | ~new_n26909_);
  assign new_n26923_ = ~new_n26912_ & new_n26765_ & (new_n26607_ ? new_n22771_ : new_n26920_);
  assign new_n26924_ = ~new_n26925_ & new_n26938_;
  assign new_n26925_ = ~new_n26936_ & new_n26926_ & (~new_n26935_ | (~new_n16524_ & new_n26937_));
  assign new_n26926_ = (~new_n26927_ | new_n26931_) & (~new_n26929_ | (new_n26933_ ? ~new_n13318_ : ~new_n26934_));
  assign new_n26927_ = new_n26636_ & new_n26928_;
  assign new_n26928_ = ~new_n16400_ & (~new_n16378_ | ~new_n21891_);
  assign new_n26929_ = ~new_n26636_ & new_n26930_;
  assign new_n26930_ = ~new_n20252_ & new_n9893_;
  assign new_n26931_ = new_n26932_ & new_n12154_ & (~new_n18890_ | (~new_n18858_ & ~new_n18888_));
  assign new_n26932_ = new_n12185_ & new_n12187_;
  assign new_n26933_ = new_n8879_ & new_n16811_ & new_n8857_;
  assign new_n26934_ = new_n26869_ & new_n18510_;
  assign new_n26935_ = ~new_n26636_ & ~new_n26930_;
  assign new_n26936_ = ~new_n26928_ & new_n26636_ & (new_n10525_ | (~new_n14876_ & new_n11726_));
  assign new_n26937_ = ~new_n12081_ & (~new_n12074_ | new_n15168_);
  assign new_n26938_ = new_n26939_ & (~new_n26929_ | (new_n13318_ & new_n26933_) | (new_n26934_ & ~new_n26933_));
  assign new_n26939_ = (new_n16524_ | ~new_n26937_ | ~new_n26935_) & (~new_n26931_ | ~new_n26927_);
  assign new_n26940_ = ~new_n26941_ & new_n26954_;
  assign new_n26941_ = new_n26942_ & (new_n26953_ | ~new_n26950_) & (new_n26952_ | new_n26948_ | ~new_n26951_);
  assign new_n26942_ = (new_n26947_ | ~new_n26946_) & (new_n21250_ | ~new_n26943_);
  assign new_n26943_ = new_n26944_ & new_n16348_;
  assign new_n26944_ = ~new_n26945_ & new_n26742_;
  assign new_n26945_ = ~new_n24324_ & ~new_n24315_ & ~new_n24322_;
  assign new_n26946_ = new_n26742_ & new_n26945_;
  assign new_n26947_ = new_n14384_ & new_n17247_;
  assign new_n26948_ = ~new_n26949_ & new_n16956_;
  assign new_n26949_ = new_n10129_ & (~new_n10159_ | ~new_n10155_);
  assign new_n26950_ = ~new_n24375_ & ~new_n26742_;
  assign new_n26951_ = ~new_n26742_ & new_n24375_;
  assign new_n26952_ = new_n16277_ & new_n26949_;
  assign new_n26953_ = (~new_n13038_ | (~new_n23769_ & (new_n23736_ | ~new_n23766_))) & (new_n15992_ | ~new_n16023_ | new_n23769_ | (~new_n23736_ & new_n23766_));
  assign new_n26954_ = new_n26955_ & (~new_n21250_ | ~new_n26943_) & (~new_n26950_ | ~new_n26953_);
  assign new_n26955_ = ~new_n26956_ & (~new_n26946_ | ~new_n26947_) & (~new_n26951_ | (~new_n26952_ & ~new_n26948_));
  assign new_n26956_ = new_n20436_ & new_n20407_ & ~new_n16348_ & new_n26944_;
  assign new_n26957_ = ~new_n26958_ & new_n26976_;
  assign new_n26958_ = new_n26959_ & ((new_n26971_ & ~new_n26974_) | (new_n26969_ & new_n26975_ & new_n25105_));
  assign new_n26959_ = new_n26968_ & new_n26960_ & (~new_n26970_ | new_n25105_ | ~new_n26969_);
  assign new_n26960_ = (~new_n26964_ | ~new_n22437_) & (new_n18750_ | ~new_n26961_);
  assign new_n26961_ = new_n26962_ & new_n14276_;
  assign new_n26962_ = ~new_n26963_ & ~new_n12908_;
  assign new_n26963_ = new_n13675_ & new_n13707_;
  assign new_n26964_ = ~new_n26967_ & new_n26965_;
  assign new_n26965_ = new_n12908_ & new_n26966_;
  assign new_n26966_ = ~new_n19345_ & new_n14070_;
  assign new_n26967_ = ~new_n24973_ & new_n16101_;
  assign new_n26968_ = (new_n15830_ | ~new_n26965_ | ~new_n26967_) & (~new_n26962_ | new_n14276_);
  assign new_n26969_ = ~new_n12908_ & new_n26963_;
  assign new_n26970_ = ~new_n13040_ & ~new_n10438_;
  assign new_n26971_ = ~new_n26973_ & new_n26972_;
  assign new_n26972_ = ~new_n26966_ & new_n12908_;
  assign new_n26973_ = ~new_n23271_ & (~new_n23273_ | new_n23330_);
  assign new_n26974_ = ~new_n20811_ & ~new_n20842_;
  assign new_n26975_ = new_n10204_ & (new_n10201_ | new_n13097_);
  assign new_n26976_ = new_n26977_ & (~new_n26973_ | ~new_n26972_) & (~new_n26964_ | new_n22437_);
  assign new_n26977_ = new_n26978_ & (~new_n18750_ | ~new_n26961_) & (~new_n26974_ | ~new_n26971_);
  assign new_n26978_ = ~new_n26969_ | (new_n25105_ ? new_n26975_ : new_n26970_);
  assign new_n26979_ = ~new_n26995_ & new_n26980_;
  assign new_n26980_ = new_n26981_ & (new_n26994_ | ~new_n26993_);
  assign new_n26981_ = new_n26982_ & (~new_n26991_ | (~new_n7732_ & new_n26848_) | (~new_n26992_ & ~new_n26848_));
  assign new_n26982_ = (~new_n12528_ | ~new_n26990_ | ~new_n26053_) & (~new_n23337_ | ~new_n26983_);
  assign new_n26983_ = new_n20968_ & new_n26984_;
  assign new_n26984_ = ~new_n14384_ & ~new_n26985_;
  assign new_n26985_ = new_n18190_ & (~new_n26986_ | (~new_n17231_ & (new_n17235_ | (~new_n26987_ & ~new_n17234_))));
  assign new_n26986_ = new_n17218_ & (\all_features[2315]  | \all_features[2316]  | \all_features[2317]  | \all_features[2318]  | \all_features[2319] );
  assign new_n26987_ = ~new_n17237_ & (new_n17239_ | (~new_n17242_ & (new_n17241_ | new_n26988_)));
  assign new_n26988_ = \all_features[2319]  & ((~new_n26989_ & \all_features[2318]  & new_n17226_) | (~new_n17224_ & ((~new_n26989_ & new_n17226_) | (~new_n17221_ & ~\all_features[2318] ))));
  assign new_n26989_ = ~\all_features[2317]  & \all_features[2318]  & \all_features[2319]  & (\all_features[2316]  ? new_n17223_ : (new_n17228_ | ~new_n17223_));
  assign new_n26990_ = ~new_n24023_ & new_n26985_;
  assign new_n26991_ = new_n24023_ & new_n26985_;
  assign new_n26992_ = ~new_n24324_ & (~new_n24322_ | (~new_n24315_ & ~new_n24293_));
  assign new_n26993_ = ~new_n26985_ & new_n14384_;
  assign new_n26994_ = (~new_n6591_ & (new_n11061_ | ~new_n6569_)) ? new_n7832_ : ~new_n12908_;
  assign new_n26995_ = new_n26998_ & new_n26996_ & (new_n26992_ | new_n26848_ | ~new_n26991_);
  assign new_n26996_ = (~new_n26983_ | new_n23337_) & (~new_n26990_ | (new_n26053_ ? new_n12528_ : ~new_n26997_));
  assign new_n26997_ = new_n21406_ & ~new_n19673_ & ~new_n21402_;
  assign new_n26998_ = new_n26999_ & (~new_n26993_ | ~new_n26994_) & (new_n26053_ | new_n26997_ | ~new_n26990_);
  assign new_n26999_ = (new_n7732_ | ~new_n26991_ | ~new_n26848_) & (new_n20968_ | ~new_n26984_ | ~new_n7558_);
  assign new_n27000_ = new_n27015_ & (~new_n27001_ | (new_n27018_ & new_n27019_));
  assign new_n27001_ = new_n27002_ & (new_n27013_ | new_n27014_ | ~new_n27012_);
  assign new_n27002_ = new_n27003_ & (~new_n23084_ | ~new_n27009_) & (new_n27011_ | new_n7581_ | ~new_n27010_);
  assign new_n27003_ = (~new_n8666_ | ~new_n27005_) & (new_n17973_ | new_n23649_ | ~new_n27004_);
  assign new_n27004_ = ~new_n24334_ & new_n7600_;
  assign new_n27005_ = ~new_n27008_ & new_n27006_;
  assign new_n27006_ = ~new_n27007_ & new_n24334_;
  assign new_n27007_ = ~new_n17414_ & (~new_n19644_ | ~new_n17392_);
  assign new_n27008_ = ~new_n14291_ & new_n11232_;
  assign new_n27009_ = new_n27006_ & new_n27008_;
  assign new_n27010_ = new_n24334_ & new_n27007_;
  assign new_n27011_ = ~new_n25379_ & ~new_n10677_;
  assign new_n27012_ = ~new_n7600_ & ~new_n24334_;
  assign new_n27013_ = new_n22998_ & (new_n14786_ | (new_n19774_ & new_n25278_));
  assign new_n27014_ = ~new_n22998_ & new_n25327_;
  assign new_n27015_ = new_n27016_ & (new_n24334_ | ((new_n27017_ | ~new_n23649_ | ~new_n7600_) & (~new_n27013_ | new_n7600_)));
  assign new_n27016_ = (~new_n27009_ | new_n23084_) & (~new_n27010_ | (new_n7581_ ? ~new_n11756_ : ~new_n27011_));
  assign new_n27017_ = new_n10308_ & (new_n10285_ | ~new_n26243_);
  assign new_n27018_ = new_n27004_ & (new_n23649_ ? new_n27017_ : new_n17973_);
  assign new_n27019_ = (new_n8666_ | ~new_n27005_) & (~new_n27012_ | ~new_n27014_);
  assign new_n27020_ = ~new_n27021_ & new_n27029_;
  assign new_n27021_ = ~new_n27022_ & new_n27026_ & (new_n27028_ | ~new_n27027_);
  assign new_n27022_ = ~new_n21535_ & ((~new_n27024_ & ~new_n19245_ & ~new_n12980_ & ~new_n27025_) | (~new_n27023_ & new_n27025_));
  assign new_n27023_ = ~new_n23606_ & (new_n24813_ | ~new_n24002_);
  assign new_n27024_ = ~new_n19541_ & (~new_n19538_ | new_n19509_);
  assign new_n27025_ = ~new_n13441_ & (~new_n13438_ | new_n13408_);
  assign new_n27026_ = ~new_n21535_ | ((new_n18754_ | ~new_n21350_ | ~new_n14292_) & (new_n13806_ | ~new_n26846_ | new_n14292_));
  assign new_n27027_ = new_n27024_ & ~new_n27025_ & ~new_n21535_;
  assign new_n27028_ = ~new_n17176_ & (~new_n17154_ | new_n17177_);
  assign new_n27029_ = (~new_n27028_ | ~new_n27027_) & (~new_n21535_ | (new_n14292_ ? new_n27030_ : new_n27031_));
  assign new_n27030_ = new_n18754_ ? ~new_n15917_ : new_n21350_;
  assign new_n27031_ = ~new_n13806_ & new_n26846_;
  assign \o[57]  = new_n27033_ ? (new_n27092_ ^ new_n27093_) : (~new_n27092_ ^ new_n27093_);
  assign new_n27033_ = new_n27034_ ? (~new_n27090_ ^ new_n27091_) : (new_n27090_ ^ new_n27091_);
  assign new_n27034_ = new_n27035_ ? (new_n27070_ ^ new_n27089_) : (~new_n27070_ ^ new_n27089_);
  assign new_n27035_ = new_n27036_ ? (new_n27055_ ^ new_n27069_) : (~new_n27055_ ^ new_n27069_);
  assign new_n27036_ = new_n27037_ ? (new_n27044_ ^ new_n27054_) : (~new_n27044_ ^ new_n27054_);
  assign new_n27037_ = new_n27038_ ? (~new_n27042_ ^ new_n27043_) : (new_n27042_ ^ new_n27043_);
  assign new_n27038_ = new_n27039_ ? (new_n27040_ ^ new_n27041_) : (~new_n27040_ ^ new_n27041_);
  assign new_n27039_ = new_n26976_ & new_n26959_;
  assign new_n27040_ = new_n26980_ & new_n26995_;
  assign new_n27041_ = new_n26772_ & new_n26783_;
  assign new_n27042_ = (new_n26752_ & new_n26771_) | (new_n26738_ & (new_n26752_ | new_n26771_));
  assign new_n27043_ = (new_n26711_ & new_n26720_) | (new_n26697_ & (new_n26711_ | new_n26720_));
  assign new_n27044_ = new_n27045_ ? (~new_n27049_ ^ new_n27050_) : (new_n27049_ ^ new_n27050_);
  assign new_n27045_ = new_n27046_ ^ new_n27048_;
  assign new_n27046_ = new_n27001_ & ~new_n27047_ & new_n27015_;
  assign new_n27047_ = ~new_n27018_ & new_n27019_;
  assign new_n27048_ = new_n26833_ & new_n26788_ & (~new_n26839_ | ~new_n26837_ | ~new_n26836_);
  assign new_n27049_ = ~new_n26787_ & ~new_n26840_;
  assign new_n27050_ = new_n27051_ ? (new_n27052_ ^ new_n27053_) : (~new_n27052_ ^ new_n27053_);
  assign new_n27051_ = new_n26739_ & new_n26750_;
  assign new_n27052_ = new_n26841_ & new_n26850_;
  assign new_n27053_ = new_n27021_ & new_n27029_;
  assign new_n27054_ = (~new_n26786_ & new_n26726_) | (~new_n26737_ & (~new_n26786_ | new_n26726_));
  assign new_n27055_ = new_n27056_ ? (~new_n27057_ ^ new_n27068_) : (new_n27057_ ^ new_n27068_);
  assign new_n27056_ = (~new_n26631_ & new_n26680_) | (~new_n26594_ & (~new_n26631_ | new_n26680_));
  assign new_n27057_ = new_n27058_ ? (new_n27063_ ^ new_n27064_) : (~new_n27063_ ^ new_n27064_);
  assign new_n27058_ = new_n27059_ ? (new_n27060_ ^ new_n27061_) : (~new_n27060_ ^ new_n27061_);
  assign new_n27059_ = new_n26862_ & new_n26877_;
  assign new_n27060_ = new_n26907_ & new_n26922_;
  assign new_n27061_ = new_n27062_ & new_n26698_ & new_n26708_;
  assign new_n27062_ = new_n19889_ & new_n26710_ & new_n26706_;
  assign new_n27063_ = (new_n26657_ & new_n26672_) | (new_n26632_ & (new_n26657_ | new_n26672_));
  assign new_n27064_ = new_n27065_ ? (new_n27066_ ^ new_n27067_) : (~new_n27066_ ^ new_n27067_);
  assign new_n27065_ = new_n26941_ & new_n26954_;
  assign new_n27066_ = new_n26753_ & new_n26769_;
  assign new_n27067_ = new_n26925_ & new_n26938_;
  assign new_n27068_ = (new_n26726_ & new_n26727_) | (~new_n26696_ & (new_n26726_ | new_n26727_));
  assign new_n27069_ = (~new_n26736_ & new_n26854_) | (~new_n26695_ & (~new_n26736_ | new_n26854_));
  assign new_n27070_ = new_n27071_ ? (~new_n27072_ ^ new_n27088_) : (new_n27072_ ^ new_n27088_);
  assign new_n27071_ = (~new_n26693_ & new_n26681_) | (~new_n26593_ & (~new_n26693_ | new_n26681_));
  assign new_n27072_ = new_n27073_ ? (~new_n27074_ ^ new_n27087_) : (new_n27074_ ^ new_n27087_);
  assign new_n27073_ = (new_n26614_ & new_n26620_) | (new_n26595_ & (new_n26614_ | new_n26620_));
  assign new_n27074_ = new_n27075_ ? (new_n27076_ ^ new_n27077_) : (~new_n27076_ ^ new_n27077_);
  assign new_n27075_ = new_n26682_ & new_n26691_;
  assign new_n27076_ = new_n26658_ & new_n26669_;
  assign new_n27077_ = new_n26672_ & new_n27078_ & (~new_n26676_ | new_n27080_);
  assign new_n27078_ = new_n27079_ & (new_n26676_ | (~new_n25035_ & new_n15494_ & new_n14469_) | (new_n21616_ & ~new_n14469_));
  assign new_n27079_ = (~new_n26678_ | new_n14782_ | ~new_n26676_) & (new_n26675_ | new_n14469_ | ~new_n21616_ | new_n26676_);
  assign new_n27080_ = (new_n27081_ | ~new_n14782_ | ~new_n26203_ | ~new_n26678_) & (new_n26678_ | (new_n26679_ & ~new_n26677_));
  assign new_n27081_ = ~new_n26201_ & (~new_n27082_ | (~new_n27083_ & ~new_n26189_));
  assign new_n27082_ = new_n26178_ & (\all_features[1651]  | \all_features[1652]  | \all_features[1653]  | \all_features[1654]  | \all_features[1655] );
  assign new_n27083_ = ~new_n26193_ & (new_n26192_ | (~new_n26195_ & (new_n26197_ | (~new_n27084_ & ~new_n26199_))));
  assign new_n27084_ = ~new_n26198_ & (~\all_features[1655]  | new_n27085_ | (~\all_features[1652]  & ~\all_features[1653]  & ~\all_features[1654] ));
  assign new_n27085_ = \all_features[1655]  & ((~new_n27086_ & ~\all_features[1653]  & \all_features[1654] ) | (~new_n26184_ & (\all_features[1654]  | (~new_n26181_ & \all_features[1653] ))));
  assign new_n27086_ = (~\all_features[1650]  & ~\all_features[1651]  & ~\all_features[1652]  & (~\all_features[1649]  | ~\all_features[1648] )) | (\all_features[1652]  & (\all_features[1650]  | \all_features[1651] ));
  assign new_n27087_ = (new_n26888_ & new_n26893_) | (new_n26883_ & (new_n26888_ | new_n26893_));
  assign new_n27088_ = (~new_n26882_ & new_n26898_) | (new_n26680_ & (~new_n26882_ | new_n26898_));
  assign new_n27089_ = (~new_n26694_ & new_n26861_) | (~new_n26592_ & (~new_n26694_ | new_n26861_));
  assign new_n27090_ = (~new_n26880_ & new_n26940_) | (~new_n26591_ & (~new_n26880_ | new_n26940_));
  assign new_n27091_ = (new_n26906_ & new_n26924_) | (~new_n26881_ & (new_n26906_ | new_n26924_));
  assign new_n27092_ = (new_n27000_ & new_n27020_) | (~new_n26589_ & (new_n27000_ | new_n27020_));
  assign new_n27093_ = (new_n26957_ & new_n26979_) | (~new_n26590_ & (new_n26957_ | new_n26979_));
  assign \o[58]  = ~new_n27095_ ^ new_n27096_;
  assign new_n27095_ = (new_n27092_ & new_n27093_) | (~new_n27033_ & (new_n27092_ | new_n27093_));
  assign new_n27096_ = new_n27097_ ^ new_n27098_;
  assign new_n27097_ = (new_n27090_ & new_n27091_) | (~new_n27034_ & (new_n27090_ | new_n27091_));
  assign new_n27098_ = new_n27099_ ? (~new_n27100_ ^ new_n27125_) : (new_n27100_ ^ new_n27125_);
  assign new_n27099_ = (~new_n27070_ & new_n27089_) | (~new_n27035_ & (~new_n27070_ | new_n27089_));
  assign new_n27100_ = new_n27101_ ? (new_n27102_ ^ new_n27119_) : (~new_n27102_ ^ new_n27119_);
  assign new_n27101_ = (~new_n27055_ & new_n27069_) | (~new_n27036_ & (~new_n27055_ | new_n27069_));
  assign new_n27102_ = new_n27103_ ? (new_n27104_ ^ new_n27115_) : (~new_n27104_ ^ new_n27115_);
  assign new_n27103_ = (~new_n27044_ & new_n27054_) | (~new_n27037_ & (~new_n27044_ | new_n27054_));
  assign new_n27104_ = new_n27105_ ? (new_n27108_ ^ new_n27109_) : (~new_n27108_ ^ new_n27109_);
  assign new_n27105_ = ~new_n27106_ ^ new_n27107_;
  assign new_n27106_ = (new_n27040_ & new_n27041_) | (new_n27039_ & (new_n27040_ | new_n27041_));
  assign new_n27107_ = (new_n27052_ & new_n27053_) | (new_n27051_ & (new_n27052_ | new_n27053_));
  assign new_n27108_ = (~new_n27049_ & ~new_n27050_) | (~new_n27045_ & (~new_n27049_ | ~new_n27050_));
  assign new_n27109_ = new_n27110_ ? (new_n27111_ ^ new_n27114_) : (~new_n27111_ ^ new_n27114_);
  assign new_n27110_ = ~new_n27046_ & ~new_n27048_;
  assign new_n27111_ = new_n27112_ ^ new_n27113_;
  assign new_n27112_ = new_n27047_ & new_n27001_ & new_n27015_;
  assign new_n27113_ = new_n26837_ & new_n26836_ & new_n26788_ & new_n26833_;
  assign new_n27114_ = new_n26698_ & ~new_n27062_ & new_n26708_;
  assign new_n27115_ = new_n27116_ ? (new_n27117_ ^ new_n27118_) : (~new_n27117_ ^ new_n27118_);
  assign new_n27116_ = (new_n27042_ & new_n27043_) | (~new_n27038_ & (new_n27042_ | new_n27043_));
  assign new_n27117_ = (~new_n27064_ & new_n27063_) | (~new_n27058_ & (~new_n27064_ | new_n27063_));
  assign new_n27118_ = (new_n27066_ & new_n27067_) | (new_n27065_ & (new_n27066_ | new_n27067_));
  assign new_n27119_ = new_n27120_ ? (~new_n27121_ ^ new_n27122_) : (new_n27121_ ^ new_n27122_);
  assign new_n27120_ = (~new_n27057_ & new_n27068_) | (new_n27056_ & (~new_n27057_ | new_n27068_));
  assign new_n27121_ = (~new_n27074_ & new_n27087_) | (new_n27073_ & (~new_n27074_ | new_n27087_));
  assign new_n27122_ = ~new_n27123_ ^ new_n27124_;
  assign new_n27123_ = (new_n27060_ & new_n27061_) | (new_n27059_ & (new_n27060_ | new_n27061_));
  assign new_n27124_ = (new_n27076_ & new_n27077_) | (new_n27075_ & (new_n27076_ | new_n27077_));
  assign new_n27125_ = (~new_n27072_ & new_n27088_) | (new_n27071_ & (~new_n27072_ | new_n27088_));
  assign \o[59]  = ((new_n27127_ | new_n27128_) & (new_n27129_ ^ new_n27130_)) | (~new_n27127_ & ~new_n27128_ & (~new_n27129_ ^ new_n27130_));
  assign new_n27127_ = ~new_n27096_ & new_n27095_;
  assign new_n27128_ = ~new_n27098_ & new_n27097_;
  assign new_n27129_ = (~new_n27100_ & new_n27125_) | (new_n27099_ & (~new_n27100_ | new_n27125_));
  assign new_n27130_ = new_n27131_ ? (~new_n27132_ ^ new_n27143_) : (new_n27132_ ^ new_n27143_);
  assign new_n27131_ = (~new_n27102_ & ~new_n27119_) | (new_n27101_ & (~new_n27102_ | ~new_n27119_));
  assign new_n27132_ = new_n27133_ ? (new_n27134_ ^ new_n27140_) : (~new_n27134_ ^ new_n27140_);
  assign new_n27133_ = (~new_n27104_ & ~new_n27115_) | (new_n27103_ & (~new_n27104_ | ~new_n27115_));
  assign new_n27134_ = new_n27135_ ? (~new_n27136_ ^ new_n27139_) : (new_n27136_ ^ new_n27139_);
  assign new_n27135_ = (~new_n27109_ & new_n27108_) | (~new_n27105_ & (~new_n27109_ | new_n27108_));
  assign new_n27136_ = new_n27137_ ^ new_n27138_;
  assign new_n27137_ = (~new_n27111_ & new_n27114_) | (~new_n27110_ & (~new_n27111_ | new_n27114_));
  assign new_n27138_ = ~new_n27112_ & ~new_n27113_;
  assign new_n27139_ = new_n27106_ & new_n27107_;
  assign new_n27140_ = ~new_n27141_ ^ new_n27142_;
  assign new_n27141_ = (new_n27117_ & new_n27118_) | (new_n27116_ & (new_n27117_ | new_n27118_));
  assign new_n27142_ = new_n27123_ & new_n27124_;
  assign new_n27143_ = (~new_n27122_ & new_n27121_) | (new_n27120_ & (~new_n27122_ | new_n27121_));
  assign \o[60]  = ~new_n27145_ ^ new_n27146_;
  assign new_n27145_ = (new_n27129_ | (~new_n27130_ & (new_n27128_ | new_n27127_))) & (new_n27128_ | new_n27127_ | ~new_n27130_);
  assign new_n27146_ = new_n27147_ ^ new_n27148_;
  assign new_n27147_ = (~new_n27132_ & new_n27143_) | (new_n27131_ & (~new_n27132_ | new_n27143_));
  assign new_n27148_ = new_n27149_ ? (~new_n27150_ ^ new_n27153_) : (new_n27150_ ^ new_n27153_);
  assign new_n27149_ = (~new_n27134_ & ~new_n27140_) | (new_n27133_ & (~new_n27134_ | ~new_n27140_));
  assign new_n27150_ = ~new_n27151_ ^ new_n27152_;
  assign new_n27151_ = (~new_n27136_ & new_n27139_) | (new_n27135_ & (~new_n27136_ | new_n27139_));
  assign new_n27152_ = ~new_n27138_ & new_n27137_;
  assign new_n27153_ = new_n27141_ & new_n27142_;
  assign \o[61]  = ((new_n27155_ | new_n27156_) & (~new_n27157_ ^ new_n27158_)) | (~new_n27155_ & ~new_n27156_ & (new_n27157_ ^ new_n27158_));
  assign new_n27155_ = ~new_n27146_ & new_n27145_;
  assign new_n27156_ = ~new_n27148_ & new_n27147_;
  assign new_n27157_ = (~new_n27150_ & new_n27153_) | (new_n27149_ & (~new_n27150_ | new_n27153_));
  assign new_n27158_ = new_n27151_ & new_n27152_;
  assign \o[62]  = (new_n27158_ | new_n27155_ | new_n27156_) & (new_n27157_ | (new_n27158_ & (new_n27155_ | new_n27156_)));
  assign \o[63]  = new_n27161_ ^ new_n27714_;
  assign new_n27161_ = new_n27162_ ? (new_n27687_ ^ new_n27701_) : (~new_n27687_ ^ new_n27701_);
  assign new_n27162_ = new_n27163_ ? (new_n27581_ ^ new_n27676_) : (~new_n27581_ ^ new_n27676_);
  assign new_n27163_ = new_n27164_ ? (new_n27343_ ^ new_n27578_) : (~new_n27343_ ^ new_n27578_);
  assign new_n27164_ = new_n27165_ ? (~new_n27303_ ^ new_n27311_) : (new_n27303_ ^ new_n27311_);
  assign new_n27165_ = new_n27166_ ? (new_n27196_ ^ new_n27302_) : (~new_n27196_ ^ new_n27302_);
  assign new_n27166_ = new_n27167_ ? (new_n27181_ ^ new_n27191_) : (~new_n27181_ ^ new_n27191_);
  assign new_n27167_ = ~new_n27168_ & new_n27178_;
  assign new_n27168_ = new_n27169_ & (~new_n19546_ | ((new_n13405_ | ~new_n13807_ | ~new_n27173_) & (~new_n25711_ | new_n27173_)));
  assign new_n27169_ = new_n27170_ & ((~new_n26932_ & ~new_n27177_) | ~new_n26921_ | new_n19546_);
  assign new_n27170_ = new_n27171_ & (new_n18916_ | ~new_n27176_);
  assign new_n27171_ = (~new_n27172_ | new_n21961_) & (~new_n27174_ | (new_n27175_ ? ~new_n15550_ : new_n16758_));
  assign new_n27172_ = new_n19546_ & ~new_n27173_ & ~new_n25711_;
  assign new_n27173_ = new_n22986_ & (new_n22982_ | new_n22956_);
  assign new_n27174_ = ~new_n19546_ & ~new_n26921_;
  assign new_n27175_ = ~new_n9414_ & new_n9388_;
  assign new_n27176_ = new_n19546_ & new_n13405_ & new_n27173_;
  assign new_n27177_ = new_n21804_ & (new_n21793_ | new_n21801_ | new_n21772_);
  assign new_n27178_ = ~new_n27180_ & new_n27179_ & (~new_n18916_ | ~new_n27176_);
  assign new_n27179_ = (new_n15550_ | ~new_n27175_ | ~new_n27174_) & (~new_n21961_ | ~new_n27172_);
  assign new_n27180_ = ~new_n19546_ & ((~new_n26932_ & ~new_n27177_ & new_n26921_) | (~new_n27175_ & new_n16758_ & ~new_n26921_));
  assign new_n27181_ = ~new_n27189_ & new_n27182_;
  assign new_n27182_ = new_n27188_ ? (new_n27184_ & (new_n23966_ | ~new_n27186_ | ~new_n12486_)) : new_n27183_;
  assign new_n27183_ = new_n25158_ & new_n24380_;
  assign new_n27184_ = (new_n8889_ | new_n12486_ | ~new_n27186_) & (new_n21768_ | ~new_n27185_ | new_n27186_);
  assign new_n27185_ = new_n10455_ & new_n20041_;
  assign new_n27186_ = new_n27187_ & new_n15477_;
  assign new_n27187_ = new_n15473_ & new_n15445_;
  assign new_n27188_ = ~new_n18321_ & new_n18290_;
  assign new_n27189_ = ~new_n27188_ | (new_n27186_ ? (new_n12486_ ? ~new_n23966_ : ~new_n8889_) : new_n27190_);
  assign new_n27190_ = ~new_n21768_ & new_n27185_;
  assign new_n27191_ = ~new_n27192_ & (new_n27193_ | ((new_n25662_ | ~new_n23607_ | ~new_n12264_) & (new_n27194_ | new_n12264_)));
  assign new_n27192_ = new_n27193_ & new_n19850_ & new_n19873_ & new_n19874_ & (~new_n7040_ | ~new_n15039_);
  assign new_n27193_ = ~new_n19318_ & (~new_n22893_ | ~new_n22880_);
  assign new_n27194_ = (~new_n11407_ & (new_n13844_ | ~new_n11409_)) ? ~new_n7269_ : new_n27195_;
  assign new_n27195_ = ~new_n24290_ & ~new_n24288_ & ~new_n24260_ & ~new_n24281_;
  assign new_n27196_ = new_n27197_ ? (new_n27242_ ^ new_n27254_) : (~new_n27242_ ^ new_n27254_);
  assign new_n27197_ = ~new_n27198_ & new_n27238_;
  assign new_n27198_ = new_n27199_ & (~new_n27236_ | ~new_n26342_ | ~new_n27202_);
  assign new_n27199_ = ~new_n27200_ | ((~new_n22363_ | ~new_n27203_) & (~new_n15284_ | ~new_n15308_ | new_n27203_));
  assign new_n27200_ = ~new_n27202_ & new_n27201_;
  assign new_n27201_ = new_n9893_ & (new_n9870_ | new_n20776_);
  assign new_n27202_ = ~new_n14749_ & (~new_n14727_ | (~new_n14751_ & ~new_n14755_));
  assign new_n27203_ = ~new_n27204_ & new_n27231_;
  assign new_n27204_ = ~new_n27230_ & (~new_n27223_ | (~new_n27228_ & (new_n27221_ | new_n27229_ | ~new_n27205_)));
  assign new_n27205_ = ~new_n27217_ & ~new_n27215_ & ((~new_n27212_ & new_n27206_) | ~new_n27220_ | ~new_n27219_);
  assign new_n27206_ = \all_features[5511]  & \all_features[5510]  & ~new_n27209_ & new_n27207_;
  assign new_n27207_ = \all_features[5511]  & (\all_features[5510]  | (new_n27208_ & (\all_features[5506]  | \all_features[5507]  | \all_features[5505] )));
  assign new_n27208_ = \all_features[5508]  & \all_features[5509] ;
  assign new_n27209_ = new_n27211_ & ~\all_features[5509]  & ~new_n27210_ & ~\all_features[5508] ;
  assign new_n27210_ = \all_features[5504]  & \all_features[5505] ;
  assign new_n27211_ = ~\all_features[5506]  & ~\all_features[5507] ;
  assign new_n27212_ = \all_features[5511]  & \all_features[5510]  & ~new_n27213_ & \all_features[5509] ;
  assign new_n27213_ = ~\all_features[5507]  & ~\all_features[5508]  & (~\all_features[5506]  | new_n27214_);
  assign new_n27214_ = ~\all_features[5504]  & ~\all_features[5505] ;
  assign new_n27215_ = ~new_n27216_ & ~\all_features[5511] ;
  assign new_n27216_ = \all_features[5509]  & \all_features[5510]  & (\all_features[5508]  | (\all_features[5506]  & \all_features[5507]  & \all_features[5505] ));
  assign new_n27217_ = ~\all_features[5511]  & (~\all_features[5510]  | ~new_n27218_ | ~new_n27210_ | ~new_n27208_);
  assign new_n27218_ = \all_features[5506]  & \all_features[5507] ;
  assign new_n27219_ = \all_features[5511]  & (\all_features[5510]  | (\all_features[5509]  & (\all_features[5508]  | ~new_n27211_ | ~new_n27214_)));
  assign new_n27220_ = \all_features[5511]  & (\all_features[5509]  | \all_features[5510]  | \all_features[5508] );
  assign new_n27221_ = ~new_n27215_ & (new_n27217_ | (new_n27220_ & (~new_n27219_ | (~new_n27222_ & new_n27207_))));
  assign new_n27222_ = ~\all_features[5509]  & \all_features[5510]  & \all_features[5511]  & (\all_features[5508]  ? new_n27211_ : (new_n27210_ | ~new_n27211_));
  assign new_n27223_ = ~new_n27227_ & ~new_n27224_ & ~new_n27226_;
  assign new_n27224_ = new_n27225_ & (~\all_features[5509]  | (~\all_features[5508]  & (~\all_features[5507]  | (~\all_features[5506]  & ~\all_features[5505] ))));
  assign new_n27225_ = ~\all_features[5510]  & ~\all_features[5511] ;
  assign new_n27226_ = ~\all_features[5509]  & new_n27225_ & ((~\all_features[5506]  & new_n27214_) | ~\all_features[5508]  | ~\all_features[5507] );
  assign new_n27227_ = new_n27225_ & (~\all_features[5507]  | ~new_n27208_ | (~\all_features[5506]  & ~new_n27210_));
  assign new_n27228_ = ~\all_features[5511]  & (~\all_features[5510]  | (~\all_features[5508]  & ~\all_features[5509]  & ~new_n27218_));
  assign new_n27229_ = ~\all_features[5511]  & (~\all_features[5510]  | (~\all_features[5509]  & (new_n27214_ | ~\all_features[5508]  | ~new_n27218_)));
  assign new_n27230_ = ~\all_features[5511]  & ~\all_features[5510]  & ~\all_features[5509]  & ~\all_features[5507]  & ~\all_features[5508] ;
  assign new_n27231_ = new_n27224_ | ~new_n27234_ | ((new_n27215_ | ~new_n27235_) & (new_n27232_ | new_n27227_));
  assign new_n27232_ = new_n27233_ & (~new_n27206_ | ~new_n27219_ | ~new_n27220_);
  assign new_n27233_ = ~new_n27217_ & ~new_n27215_ & ~new_n27228_ & ~new_n27229_;
  assign new_n27234_ = ~new_n27226_ & ~new_n27230_;
  assign new_n27235_ = ~new_n27227_ & ~new_n27217_ & ~new_n27228_ & ~new_n27229_;
  assign new_n27236_ = (new_n8666_ & (~new_n10876_ | new_n8663_)) ? new_n27237_ : new_n14181_;
  assign new_n27237_ = new_n7432_ & (new_n7438_ | new_n7410_);
  assign new_n27238_ = ~new_n27239_ & (new_n27202_ ? (new_n26342_ ? new_n27236_ : ~new_n27240_) : new_n27201_);
  assign new_n27239_ = new_n27200_ & ~new_n22363_ & new_n27203_;
  assign new_n27240_ = (~new_n27241_ | new_n13806_) & (~new_n26733_ | ~new_n19813_ | ~new_n13806_);
  assign new_n27241_ = new_n26065_ & ~new_n13127_ & ~new_n13130_;
  assign new_n27242_ = ~new_n27243_ & new_n27251_;
  assign new_n27243_ = ~new_n27244_ & (new_n27246_ ? ~new_n25915_ : (new_n27247_ ? ~new_n27249_ : new_n27248_));
  assign new_n27244_ = new_n27245_ & new_n14293_;
  assign new_n27245_ = new_n26849_ & ~new_n25915_ & new_n27246_;
  assign new_n27246_ = ~new_n17840_ & (~new_n20164_ | ~new_n25110_);
  assign new_n27247_ = ~new_n15215_ & new_n16764_;
  assign new_n27248_ = ~new_n26891_ & (new_n15082_ | (~new_n25357_ & new_n15079_));
  assign new_n27249_ = new_n10871_ & ~new_n17932_ & ~new_n27250_;
  assign new_n27250_ = ~new_n21387_ & (~new_n21382_ | ~new_n21357_);
  assign new_n27251_ = new_n27252_ & (new_n14293_ | ~new_n27245_);
  assign new_n27252_ = (new_n27246_ | (new_n27247_ ? ~new_n27250_ : ~new_n27248_)) & (~new_n27253_ | new_n25915_ | ~new_n27246_);
  assign new_n27253_ = ~new_n18174_ & ~new_n26849_;
  assign new_n27254_ = ~new_n27255_ & new_n27300_;
  assign new_n27255_ = new_n27261_ & (~new_n27262_ | ((new_n27256_ | ~new_n27297_) & (new_n27264_ | ~new_n27298_ | new_n27297_)));
  assign new_n27256_ = new_n18563_ & new_n10838_ & new_n10871_ & ~new_n27257_ & new_n18547_;
  assign new_n27257_ = new_n18569_ & (new_n18553_ | new_n18561_ | (~new_n18551_ & ~new_n27258_ & ~new_n18555_));
  assign new_n27258_ = \all_features[2959]  & (new_n27259_ | ~new_n18559_ | ~new_n18558_) & (new_n27260_ | \all_features[2958] );
  assign new_n27259_ = new_n18560_ & \all_features[2957]  & ((~new_n18562_ & \all_features[2954] ) | \all_features[2956]  | \all_features[2955] );
  assign new_n27260_ = \all_features[2957]  & (\all_features[2954]  | \all_features[2955]  | \all_features[2956]  | ~new_n18562_);
  assign new_n27261_ = new_n27262_ | ~new_n27263_ | (new_n13098_ & ~new_n9027_);
  assign new_n27262_ = ~new_n8956_ & (~new_n8930_ | new_n15868_);
  assign new_n27263_ = new_n21591_ & (~new_n21592_ | ~new_n13758_);
  assign new_n27264_ = ~new_n27265_ & new_n27293_;
  assign new_n27265_ = ~new_n27292_ & (new_n27285_ | new_n27288_ | new_n27290_ | new_n27291_ | new_n27266_);
  assign new_n27266_ = ~new_n27279_ & ~new_n27284_ & ((~new_n27267_ & new_n27276_) | new_n27283_ | new_n27281_);
  assign new_n27267_ = new_n27268_ & (new_n27274_ | ~\all_features[2949]  | ~\all_features[2950]  | ~\all_features[2951] );
  assign new_n27268_ = \all_features[2951]  & \all_features[2950]  & ~new_n27269_ & new_n27272_;
  assign new_n27269_ = new_n27270_ & ~\all_features[2949]  & ~new_n27271_ & ~\all_features[2948] ;
  assign new_n27270_ = ~\all_features[2946]  & ~\all_features[2947] ;
  assign new_n27271_ = \all_features[2944]  & \all_features[2945] ;
  assign new_n27272_ = \all_features[2951]  & (\all_features[2950]  | (new_n27273_ & (\all_features[2946]  | \all_features[2947]  | \all_features[2945] )));
  assign new_n27273_ = \all_features[2948]  & \all_features[2949] ;
  assign new_n27274_ = ~\all_features[2947]  & ~\all_features[2948]  & (~\all_features[2946]  | new_n27275_);
  assign new_n27275_ = ~\all_features[2944]  & ~\all_features[2945] ;
  assign new_n27276_ = new_n27277_ & new_n27278_;
  assign new_n27277_ = \all_features[2951]  & (\all_features[2950]  | (\all_features[2949]  & (\all_features[2948]  | ~new_n27275_ | ~new_n27270_)));
  assign new_n27278_ = \all_features[2951]  & (\all_features[2949]  | \all_features[2950]  | \all_features[2948] );
  assign new_n27279_ = ~\all_features[2951]  & (~\all_features[2950]  | (~\all_features[2949]  & (new_n27275_ | ~new_n27280_ | ~\all_features[2948] )));
  assign new_n27280_ = \all_features[2946]  & \all_features[2947] ;
  assign new_n27281_ = ~new_n27282_ & ~\all_features[2951] ;
  assign new_n27282_ = \all_features[2949]  & \all_features[2950]  & (\all_features[2948]  | (\all_features[2946]  & \all_features[2947]  & \all_features[2945] ));
  assign new_n27283_ = ~\all_features[2951]  & (~\all_features[2950]  | ~new_n27271_ | ~new_n27273_ | ~new_n27280_);
  assign new_n27284_ = ~\all_features[2951]  & (~\all_features[2950]  | (~\all_features[2948]  & ~\all_features[2949]  & ~new_n27280_));
  assign new_n27285_ = ~new_n27284_ & (new_n27279_ | (~new_n27281_ & (new_n27283_ | new_n27286_)));
  assign new_n27286_ = new_n27278_ & (~new_n27277_ | (~new_n27287_ & new_n27272_));
  assign new_n27287_ = ~\all_features[2949]  & \all_features[2950]  & \all_features[2951]  & (\all_features[2948]  ? new_n27270_ : (new_n27271_ | ~new_n27270_));
  assign new_n27288_ = new_n27289_ & (~\all_features[2949]  | (~\all_features[2948]  & (~\all_features[2947]  | (~\all_features[2946]  & ~\all_features[2945] ))));
  assign new_n27289_ = ~\all_features[2950]  & ~\all_features[2951] ;
  assign new_n27290_ = new_n27289_ & (~\all_features[2947]  | ~new_n27273_ | (~\all_features[2946]  & ~new_n27271_));
  assign new_n27291_ = ~\all_features[2949]  & new_n27289_ & ((~\all_features[2946]  & new_n27275_) | ~\all_features[2948]  | ~\all_features[2947] );
  assign new_n27292_ = ~\all_features[2951]  & ~\all_features[2950]  & ~\all_features[2949]  & ~\all_features[2947]  & ~\all_features[2948] ;
  assign new_n27293_ = new_n27288_ | ~new_n27295_ | ((new_n27281_ | ~new_n27296_) & (new_n27294_ | new_n27290_));
  assign new_n27294_ = ~new_n27279_ & ~new_n27281_ & ~new_n27283_ & ~new_n27284_ & (~new_n27276_ | ~new_n27268_);
  assign new_n27295_ = ~new_n27291_ & ~new_n27292_;
  assign new_n27296_ = ~new_n27290_ & ~new_n27284_ & ~new_n27279_ & ~new_n27283_;
  assign new_n27297_ = ~new_n20623_ & (~new_n20620_ | ~new_n20612_);
  assign new_n27298_ = new_n27299_ & new_n25868_ & new_n25892_;
  assign new_n27299_ = new_n25896_ & new_n25899_;
  assign new_n27300_ = new_n27262_ ? ((~new_n27256_ & new_n27297_) | (~new_n27264_ & new_n27298_ & ~new_n27297_)) : new_n27301_;
  assign new_n27301_ = (~new_n22175_ | new_n27263_) & (new_n9027_ | ~new_n13098_ | ~new_n27263_);
  assign new_n27302_ = new_n27243_ & new_n27251_;
  assign new_n27303_ = new_n27304_ & new_n27308_;
  assign new_n27304_ = new_n22036_ ? new_n27305_ : ((~new_n27307_ | new_n24179_) & (new_n14654_ | new_n20852_ | ~new_n24179_));
  assign new_n27305_ = (~new_n27306_ | ~new_n24395_) & (new_n24359_ | ~new_n25011_ | new_n24395_);
  assign new_n27306_ = new_n12908_ & new_n21693_;
  assign new_n27307_ = new_n13806_ ? (~new_n14947_ | (~new_n20730_ & ~new_n14924_)) : ~new_n19349_;
  assign new_n27308_ = new_n27309_ & (new_n22036_ | (new_n27307_ & ~new_n24179_) | (new_n27310_ & new_n24179_));
  assign new_n27309_ = ~new_n22036_ | (~new_n24359_ & new_n25011_ & ~new_n24395_) | (new_n27306_ & new_n24395_);
  assign new_n27310_ = new_n20852_ ? new_n24752_ : ~new_n14654_;
  assign new_n27311_ = ~new_n27312_ & new_n27341_;
  assign new_n27312_ = new_n27313_ & new_n27318_;
  assign new_n27313_ = (~new_n23592_ | (new_n27316_ ? ~new_n27317_ : ~new_n27314_)) & (new_n27315_ | new_n24033_ | new_n23592_);
  assign new_n27314_ = ~new_n24373_ & new_n14416_ & (new_n14394_ | ~new_n14417_);
  assign new_n27315_ = new_n13063_ & (~new_n7991_ | (~new_n7958_ & ~new_n7988_));
  assign new_n27316_ = ~new_n15264_ & (~new_n15244_ | new_n16763_);
  assign new_n27317_ = ~new_n23147_ & ~new_n13038_;
  assign new_n27318_ = ~new_n27321_ & (~new_n27319_ | ~new_n27320_) & (~new_n27322_ | (~new_n27323_ & ~new_n27324_));
  assign new_n27319_ = new_n24373_ & new_n15906_ & (new_n15904_ | ~new_n23075_);
  assign new_n27320_ = ~new_n27316_ & new_n23592_;
  assign new_n27321_ = new_n23592_ & new_n27316_ & ~new_n7445_ & ~new_n27317_;
  assign new_n27322_ = ~new_n23592_ & new_n24033_;
  assign new_n27323_ = ~new_n9193_ & new_n19507_;
  assign new_n27324_ = ~new_n27336_ & new_n27337_;
  assign new_n27336_ = ~\all_features[4895]  & ~\all_features[4894]  & ~\all_features[4893]  & ~\all_features[4891]  & ~\all_features[4892] ;
  assign new_n27337_ = \all_features[4894]  | \all_features[4895]  | (~new_n27338_ & \all_features[4893]  & new_n27340_);
  assign new_n27338_ = ~\all_features[4892]  & (~\all_features[4891]  | (~\all_features[4890]  & ~\all_features[4889] ));
  assign new_n27340_ = \all_features[4891]  & \all_features[4892]  & \all_features[4893]  & (\all_features[4890]  | (\all_features[4889]  & \all_features[4888] ));
  assign new_n27341_ = new_n27342_ & (new_n27319_ | new_n27314_ | ~new_n27320_);
  assign new_n27342_ = new_n23592_ | ((~new_n27315_ | new_n24033_) & (new_n27323_ | new_n27324_ | ~new_n24033_));
  assign new_n27343_ = new_n27344_ ? (new_n27428_ ^ new_n27303_) : (~new_n27428_ ^ new_n27303_);
  assign new_n27344_ = new_n27345_ ? (~new_n27386_ ^ new_n27427_) : (new_n27386_ ^ new_n27427_);
  assign new_n27345_ = new_n27346_ ? (~new_n27371_ ^ new_n27378_) : (new_n27371_ ^ new_n27378_);
  assign new_n27346_ = ~new_n27347_ & new_n27367_;
  assign new_n27347_ = ~new_n27366_ & new_n27354_ & new_n27348_ & (new_n27358_ | ~new_n16026_ | ~new_n27356_);
  assign new_n27348_ = (~new_n27351_ | ~new_n27352_ | ~new_n27353_) & (~new_n14918_ | ~new_n27349_);
  assign new_n27349_ = ~new_n6532_ & new_n27350_;
  assign new_n27350_ = new_n19544_ & new_n27293_;
  assign new_n27351_ = ~new_n19544_ & new_n27293_;
  assign new_n27352_ = new_n11407_ & (new_n11409_ | ~new_n13844_);
  assign new_n27353_ = ~\all_features[5351]  & ~\all_features[5350]  & ~\all_features[5349]  & ~\all_features[5347]  & ~\all_features[5348] ;
  assign new_n27354_ = (~new_n27360_ | ~new_n27355_) & (~new_n27359_ | (new_n8164_ ? ~new_n27361_ : new_n16758_));
  assign new_n27355_ = new_n27356_ & new_n27358_;
  assign new_n27356_ = ~new_n27293_ & new_n27357_;
  assign new_n27357_ = ~new_n16354_ & ~new_n9995_;
  assign new_n27358_ = ~new_n19509_ & new_n21562_;
  assign new_n27359_ = ~new_n27357_ & ~new_n27293_;
  assign new_n27360_ = ~new_n13203_ & new_n11674_;
  assign new_n27361_ = ~new_n25096_ & (~new_n25101_ | (~new_n27362_ & new_n25103_ & new_n25083_));
  assign new_n27362_ = ~new_n25090_ & ~new_n25095_ & ((~new_n27363_ & new_n27365_) | new_n25094_ | new_n25092_);
  assign new_n27363_ = ~new_n25087_ & new_n25085_ & \all_features[2070]  & \all_features[2071]  & (~\all_features[2069]  | new_n27364_);
  assign new_n27364_ = ~\all_features[2067]  & ~\all_features[2068]  & (~\all_features[2066]  | (~\all_features[2065]  & ~\all_features[2064] ));
  assign new_n27365_ = \all_features[2071]  & (\all_features[2070]  | new_n25089_);
  assign new_n27366_ = new_n27350_ & new_n6532_ & (new_n8225_ | (new_n24524_ & new_n8202_));
  assign new_n27367_ = new_n27368_ & new_n27370_;
  assign new_n27368_ = (new_n14918_ | ~new_n27349_) & (~new_n27351_ | (~new_n27369_ & (new_n27352_ | ~new_n27353_)));
  assign new_n27369_ = ~new_n7192_ & ~new_n27353_ & (~new_n7164_ | ~new_n22779_);
  assign new_n27370_ = (~new_n27355_ | new_n27360_) & (~new_n27359_ | (new_n8164_ ? new_n27361_ : ~new_n16758_));
  assign new_n27371_ = ~new_n27372_ & new_n27377_;
  assign new_n27372_ = new_n27375_ & (new_n25711_ | (new_n27373_ & (new_n23337_ | ~new_n18797_ | ~new_n24395_)));
  assign new_n27373_ = (new_n11633_ | new_n18797_ | ~new_n24395_) & (new_n21355_ | ~new_n27374_ | new_n24395_);
  assign new_n27374_ = ~new_n12872_ & new_n12900_;
  assign new_n27375_ = ~new_n25711_ & (new_n24395_ | new_n27374_ | new_n25711_ | new_n7942_);
  assign new_n27377_ = new_n25711_ | ((new_n27374_ | ~new_n7942_ | new_n24395_) & (~new_n18797_ | ~new_n23337_ | ~new_n24395_));
  assign new_n27378_ = (new_n27379_ & (new_n19147_ | ~new_n16026_ | ~new_n24023_)) | (new_n27385_ & ~new_n19147_ & new_n16026_ & new_n24023_);
  assign new_n27379_ = ~new_n27380_ & ((~new_n27383_ & (~new_n24077_ | new_n24023_)) | (~new_n24023_ & (new_n27384_ | (~new_n27382_ & ~new_n24077_))));
  assign new_n27380_ = new_n24023_ & new_n19147_ & ~new_n27381_ & ~new_n14206_;
  assign new_n27381_ = new_n6799_ & (new_n6801_ | new_n25349_);
  assign new_n27382_ = ~new_n7039_ & (~new_n7036_ | ~new_n7003_);
  assign new_n27383_ = ~new_n24023_ | (new_n19147_ ? (new_n27381_ ? new_n8992_ : ~new_n14206_) : new_n16026_);
  assign new_n27384_ = new_n17813_ & ~new_n11517_ & ~new_n11541_;
  assign new_n27385_ = new_n21166_ & (new_n21422_ | new_n21414_ | new_n21431_);
  assign new_n27386_ = ~new_n27387_ & new_n27426_;
  assign new_n27387_ = new_n27388_ & ~new_n27425_ & (new_n24812_ | new_n26911_ | new_n27391_ | ~new_n7556_);
  assign new_n27388_ = (~new_n27424_ & new_n27423_ & new_n27391_) | (~new_n27391_ & (new_n24812_ | ~new_n27389_));
  assign new_n27389_ = ~new_n7556_ & new_n20406_ & (new_n20365_ | new_n20371_);
  assign new_n27391_ = ~new_n27392_ & (new_n27407_ | new_n27409_ | new_n27401_ | new_n27418_ | ~new_n27422_);
  assign new_n27392_ = new_n27414_ & (new_n27393_ | new_n27417_) & (new_n27407_ | new_n27401_ | new_n27419_);
  assign new_n27393_ = ~new_n27409_ & (new_n27412_ | (~new_n27413_ & (new_n27411_ | (~new_n27407_ & ~new_n27394_))));
  assign new_n27394_ = ~new_n27401_ & (~new_n27405_ | (new_n27395_ & (~new_n27404_ | (~new_n27406_ & new_n27398_))));
  assign new_n27395_ = \all_features[5959]  & (\all_features[5958]  | new_n27396_);
  assign new_n27396_ = \all_features[5957]  & (\all_features[5954]  | \all_features[5955]  | \all_features[5956]  | ~new_n27397_);
  assign new_n27397_ = ~\all_features[5952]  & ~\all_features[5953] ;
  assign new_n27398_ = \all_features[5959]  & ~new_n27399_ & \all_features[5958] ;
  assign new_n27399_ = ~\all_features[5957]  & ~\all_features[5956]  & ~\all_features[5955]  & ~new_n27400_ & ~\all_features[5954] ;
  assign new_n27400_ = \all_features[5952]  & \all_features[5953] ;
  assign new_n27401_ = ~\all_features[5959]  & (~\all_features[5958]  | ~new_n27400_ | ~new_n27402_ | ~new_n27403_);
  assign new_n27402_ = \all_features[5954]  & \all_features[5955] ;
  assign new_n27403_ = \all_features[5956]  & \all_features[5957] ;
  assign new_n27404_ = \all_features[5959]  & (\all_features[5958]  | (new_n27403_ & (\all_features[5954]  | \all_features[5955]  | \all_features[5953] )));
  assign new_n27405_ = \all_features[5959]  & (\all_features[5957]  | \all_features[5958]  | \all_features[5956] );
  assign new_n27406_ = \all_features[5958]  & \all_features[5959]  & (\all_features[5957]  | (\all_features[5956]  & (\all_features[5955]  | \all_features[5954] )));
  assign new_n27407_ = ~new_n27408_ & ~\all_features[5959] ;
  assign new_n27408_ = \all_features[5957]  & \all_features[5958]  & (\all_features[5956]  | (\all_features[5954]  & \all_features[5955]  & \all_features[5953] ));
  assign new_n27409_ = new_n27410_ & (~\all_features[5957]  | (~\all_features[5956]  & (~\all_features[5955]  | (~\all_features[5954]  & ~\all_features[5953] ))));
  assign new_n27410_ = ~\all_features[5958]  & ~\all_features[5959] ;
  assign new_n27411_ = ~\all_features[5959]  & (~\all_features[5958]  | (~\all_features[5957]  & (new_n27397_ | ~\all_features[5956]  | ~new_n27402_)));
  assign new_n27412_ = new_n27410_ & (~\all_features[5955]  | ~new_n27403_ | (~\all_features[5954]  & ~new_n27400_));
  assign new_n27413_ = ~\all_features[5959]  & (~\all_features[5958]  | (~\all_features[5956]  & ~\all_features[5957]  & ~new_n27402_));
  assign new_n27414_ = new_n27416_ & ~new_n27411_ & (new_n27407_ | new_n27401_ | new_n27415_ | new_n27413_);
  assign new_n27415_ = new_n27405_ & new_n27404_ & new_n27395_ & new_n27398_;
  assign new_n27416_ = ~new_n27418_ & ~new_n27413_ & ~new_n27417_ & ~new_n27409_ & ~new_n27412_;
  assign new_n27417_ = ~\all_features[5957]  & new_n27410_ & ((~\all_features[5954]  & new_n27397_) | ~\all_features[5956]  | ~\all_features[5955] );
  assign new_n27418_ = ~\all_features[5959]  & ~\all_features[5958]  & ~\all_features[5957]  & ~\all_features[5955]  & ~\all_features[5956] ;
  assign new_n27419_ = new_n27405_ & ~new_n27420_ & new_n27395_;
  assign new_n27420_ = ~new_n27399_ & new_n27404_ & \all_features[5958]  & \all_features[5959]  & (~\all_features[5957]  | new_n27421_);
  assign new_n27421_ = ~\all_features[5955]  & ~\all_features[5956]  & (~\all_features[5954]  | new_n27397_);
  assign new_n27422_ = ~new_n27413_ & ~new_n27417_ & ~new_n27411_ & ~new_n27412_;
  assign new_n27423_ = ~new_n13707_ & (~new_n7736_ | new_n22708_);
  assign new_n27424_ = ~new_n19630_ & (~new_n19606_ | ~new_n19632_);
  assign new_n27425_ = ~new_n27391_ & new_n24812_ & (new_n18594_ ? new_n14278_ : new_n22998_);
  assign new_n27426_ = (~new_n27423_ | new_n27424_ | ~new_n27391_) & (new_n24812_ | ~new_n26911_ | ~new_n7556_ | new_n27391_);
  assign new_n27427_ = new_n27182_ & new_n27189_;
  assign new_n27428_ = new_n27429_ ? (new_n27544_ ^ new_n27427_) : (~new_n27544_ ^ new_n27427_);
  assign new_n27429_ = new_n27430_ ? (new_n27453_ ^ new_n27533_) : (~new_n27453_ ^ new_n27533_);
  assign new_n27430_ = ~new_n27431_ & new_n27451_;
  assign new_n27431_ = ~new_n27432_ & new_n27448_;
  assign new_n27432_ = new_n27433_ & (new_n24007_ | ~new_n27444_) & (new_n16570_ | new_n23319_ | ~new_n27447_);
  assign new_n27433_ = (~new_n27434_ | new_n27438_) & (~new_n27437_ | (new_n27443_ ? new_n27439_ : new_n26768_));
  assign new_n27434_ = new_n27435_ & new_n27436_;
  assign new_n27435_ = ~new_n24564_ & ~new_n17975_;
  assign new_n27436_ = ~new_n12257_ & (~new_n12254_ | ~new_n12229_);
  assign new_n27437_ = ~new_n24564_ & new_n17975_;
  assign new_n27438_ = ~new_n23132_ & ~new_n12398_;
  assign new_n27439_ = new_n17359_ & (new_n17387_ | (~new_n27440_ & ~new_n17386_));
  assign new_n27440_ = ~new_n17375_ & (new_n17377_ | (~new_n17381_ & (new_n17372_ | (~new_n17378_ & ~new_n27441_))));
  assign new_n27441_ = ~new_n17380_ & (~new_n17371_ | (new_n17370_ & (~new_n17365_ | (~new_n27442_ & new_n17367_))));
  assign new_n27442_ = \all_features[3862]  & \all_features[3863]  & (\all_features[3861]  | (~new_n17368_ & \all_features[3860] ));
  assign new_n27443_ = new_n17517_ & new_n17518_;
  assign new_n27444_ = ~new_n27446_ & new_n27445_;
  assign new_n27445_ = ~new_n18574_ & new_n24564_;
  assign new_n27446_ = ~new_n20205_ & new_n23078_;
  assign new_n27447_ = new_n18574_ & new_n24564_;
  assign new_n27448_ = new_n27449_ & (new_n27436_ | ~new_n16761_ | ~new_n27435_) & (new_n8060_ | ~new_n27450_);
  assign new_n27449_ = (~new_n24007_ | ~new_n27444_) & (~new_n27447_ | (new_n23319_ ? new_n19160_ : ~new_n16570_));
  assign new_n27450_ = new_n27445_ & new_n27446_;
  assign new_n27451_ = new_n27452_ & (~new_n27447_ | ~new_n23319_ | ~new_n19160_) & (~new_n27450_ | ~new_n8060_);
  assign new_n27452_ = (~new_n27438_ | ~new_n27434_) & (~new_n27437_ | (new_n27443_ ? ~new_n27439_ : ~new_n26768_));
  assign new_n27453_ = new_n27454_ & (~new_n27500_ | new_n27493_);
  assign new_n27454_ = new_n27455_ & (~new_n27491_ | (~new_n19717_ & new_n27492_) | (~new_n22361_ & ~new_n27492_));
  assign new_n27455_ = ~new_n27460_ & (~new_n27458_ | ~new_n27490_) & (~new_n27456_ | new_n27489_);
  assign new_n27456_ = ~new_n24922_ & new_n27457_;
  assign new_n27457_ = ~new_n23184_ & ~new_n25918_;
  assign new_n27458_ = new_n27459_ & new_n16899_;
  assign new_n27459_ = ~new_n11824_ & new_n23184_;
  assign new_n27460_ = new_n27461_ & new_n27241_ & (new_n27488_ | ~new_n27478_) & (new_n27462_ | new_n27488_);
  assign new_n27461_ = new_n23184_ & new_n11824_;
  assign new_n27462_ = new_n27478_ & (new_n27485_ | (~new_n27484_ & new_n27463_ & (new_n27472_ | new_n27482_)));
  assign new_n27463_ = ~new_n27472_ & ~new_n27474_ & (~new_n27477_ | ~new_n27476_ | new_n27464_);
  assign new_n27464_ = new_n27465_ & ~new_n27470_ & new_n27467_;
  assign new_n27465_ = \all_features[5767]  & (\all_features[5766]  | (new_n27466_ & (\all_features[5762]  | \all_features[5763]  | \all_features[5761] )));
  assign new_n27466_ = \all_features[5764]  & \all_features[5765] ;
  assign new_n27467_ = new_n27469_ & (\all_features[5764]  | \all_features[5765]  | ~new_n27468_ | (\all_features[5761]  & \all_features[5760] ));
  assign new_n27468_ = ~\all_features[5762]  & ~\all_features[5763] ;
  assign new_n27469_ = \all_features[5766]  & \all_features[5767] ;
  assign new_n27470_ = new_n27469_ & \all_features[5765]  & ((~new_n27471_ & \all_features[5762] ) | \all_features[5764]  | \all_features[5763] );
  assign new_n27471_ = ~\all_features[5760]  & ~\all_features[5761] ;
  assign new_n27472_ = ~new_n27473_ & ~\all_features[5767] ;
  assign new_n27473_ = \all_features[5765]  & \all_features[5766]  & (\all_features[5764]  | (\all_features[5762]  & \all_features[5763]  & \all_features[5761] ));
  assign new_n27474_ = ~\all_features[5767]  & (~new_n27466_ | ~\all_features[5760]  | ~\all_features[5761]  | ~\all_features[5766]  | ~new_n27475_);
  assign new_n27475_ = \all_features[5762]  & \all_features[5763] ;
  assign new_n27476_ = \all_features[5767]  & (\all_features[5766]  | (\all_features[5765]  & (\all_features[5764]  | ~new_n27468_ | ~new_n27471_)));
  assign new_n27477_ = \all_features[5767]  & (\all_features[5765]  | \all_features[5766]  | \all_features[5764] );
  assign new_n27478_ = \all_features[5766]  | \all_features[5767]  | (~new_n27481_ & new_n27480_ & \all_features[5765] );
  assign new_n27480_ = new_n27466_ & \all_features[5763]  & (\all_features[5762]  | (\all_features[5760]  & \all_features[5761] ));
  assign new_n27481_ = ~\all_features[5764]  & (~\all_features[5763]  | (~\all_features[5762]  & ~\all_features[5761] ));
  assign new_n27482_ = ~new_n27474_ & (~new_n27477_ | (new_n27476_ & (~new_n27465_ | (~new_n27483_ & new_n27467_))));
  assign new_n27483_ = new_n27469_ & (\all_features[5765]  | (~new_n27468_ & \all_features[5764] ));
  assign new_n27484_ = ~\all_features[5767]  & (~\all_features[5766]  | (~\all_features[5765]  & (new_n27471_ | ~\all_features[5764]  | ~new_n27475_)));
  assign new_n27485_ = ~\all_features[5767]  & (~\all_features[5766]  | (~\all_features[5764]  & ~\all_features[5765]  & ~new_n27475_));
  assign new_n27488_ = ~\all_features[5767]  & ~\all_features[5766]  & ~\all_features[5765]  & ~\all_features[5763]  & ~\all_features[5764] ;
  assign new_n27489_ = ~new_n26642_ & new_n25709_;
  assign new_n27490_ = ~new_n9275_ & (~new_n9249_ | ~new_n12529_);
  assign new_n27491_ = ~new_n23184_ & new_n25918_;
  assign new_n27492_ = new_n14317_ & (new_n14295_ | ~new_n14320_);
  assign new_n27493_ = ~new_n27494_ & (~new_n27495_ | (new_n27496_ & (new_n27492_ | new_n22361_ | ~new_n27491_)));
  assign new_n27494_ = new_n27456_ & new_n27489_;
  assign new_n27495_ = (new_n19717_ | ~new_n27492_ | ~new_n27491_) & (~new_n27458_ | new_n27490_);
  assign new_n27496_ = (new_n22543_ | ~new_n27498_) & (new_n27499_ | ~new_n27497_);
  assign new_n27497_ = ~new_n27241_ & new_n27461_;
  assign new_n27498_ = ~new_n16899_ & new_n27459_;
  assign new_n27499_ = ~new_n10516_ & new_n10490_;
  assign new_n27500_ = (~new_n27498_ | ~new_n22543_) & (~new_n27457_ | ~new_n27501_) & (~new_n27497_ | ~new_n27499_);
  assign new_n27501_ = ~new_n27502_ & new_n24922_;
  assign new_n27502_ = new_n27527_ & (~new_n27503_ | (~new_n27522_ & (new_n27523_ | (~new_n27531_ & ~new_n27524_))));
  assign new_n27503_ = ~new_n27525_ & new_n27520_ & (new_n27522_ | (~new_n27504_ & ~new_n27523_ & ~new_n27524_));
  assign new_n27504_ = ~new_n27516_ & ~new_n27514_ & ((~new_n27511_ & new_n27505_) | ~new_n27519_ | ~new_n27518_);
  assign new_n27505_ = \all_features[1847]  & \all_features[1846]  & ~new_n27508_ & new_n27506_;
  assign new_n27506_ = \all_features[1847]  & (\all_features[1846]  | (new_n27507_ & (\all_features[1842]  | \all_features[1843]  | \all_features[1841] )));
  assign new_n27507_ = \all_features[1844]  & \all_features[1845] ;
  assign new_n27508_ = new_n27510_ & ~\all_features[1845]  & ~new_n27509_ & ~\all_features[1844] ;
  assign new_n27509_ = \all_features[1840]  & \all_features[1841] ;
  assign new_n27510_ = ~\all_features[1842]  & ~\all_features[1843] ;
  assign new_n27511_ = \all_features[1847]  & \all_features[1846]  & ~new_n27512_ & \all_features[1845] ;
  assign new_n27512_ = ~\all_features[1843]  & ~\all_features[1844]  & (~\all_features[1842]  | new_n27513_);
  assign new_n27513_ = ~\all_features[1840]  & ~\all_features[1841] ;
  assign new_n27514_ = ~new_n27515_ & ~\all_features[1847] ;
  assign new_n27515_ = \all_features[1845]  & \all_features[1846]  & (\all_features[1844]  | (\all_features[1842]  & \all_features[1843]  & \all_features[1841] ));
  assign new_n27516_ = ~\all_features[1847]  & (~\all_features[1846]  | ~new_n27509_ | ~new_n27507_ | ~new_n27517_);
  assign new_n27517_ = \all_features[1842]  & \all_features[1843] ;
  assign new_n27518_ = \all_features[1847]  & (\all_features[1846]  | (\all_features[1845]  & (\all_features[1844]  | ~new_n27510_ | ~new_n27513_)));
  assign new_n27519_ = \all_features[1847]  & (\all_features[1845]  | \all_features[1846]  | \all_features[1844] );
  assign new_n27520_ = \all_features[1845]  | \all_features[1846]  | \all_features[1847]  | (\all_features[1844]  & \all_features[1843]  & ~new_n27521_);
  assign new_n27521_ = ~\all_features[1842]  & new_n27513_;
  assign new_n27522_ = ~\all_features[1846]  & ~\all_features[1847]  & (~\all_features[1843]  | ~new_n27507_ | (~\all_features[1842]  & ~new_n27509_));
  assign new_n27523_ = ~\all_features[1847]  & (~\all_features[1846]  | (~\all_features[1844]  & ~\all_features[1845]  & ~new_n27517_));
  assign new_n27524_ = ~\all_features[1847]  & (~\all_features[1846]  | (~\all_features[1845]  & (new_n27513_ | ~\all_features[1844]  | ~new_n27517_)));
  assign new_n27525_ = ~\all_features[1847]  & ~new_n27526_ & ~\all_features[1846] ;
  assign new_n27526_ = \all_features[1845]  & (\all_features[1844]  | (\all_features[1843]  & (\all_features[1842]  | \all_features[1841] )));
  assign new_n27527_ = new_n27525_ | ~new_n27520_ | ((new_n27522_ | new_n27530_) & (new_n27514_ | ~new_n27528_));
  assign new_n27528_ = new_n27529_ & ~new_n27522_ & ~new_n27524_;
  assign new_n27529_ = ~new_n27523_ & ~new_n27516_;
  assign new_n27530_ = ~new_n27514_ & ~new_n27524_ & new_n27529_ & (~new_n27519_ | ~new_n27518_ | ~new_n27505_);
  assign new_n27531_ = ~new_n27514_ & (new_n27516_ | (new_n27519_ & (~new_n27518_ | (~new_n27532_ & new_n27506_))));
  assign new_n27532_ = ~\all_features[1845]  & \all_features[1846]  & \all_features[1847]  & (\all_features[1844]  ? new_n27510_ : (new_n27509_ | ~new_n27510_));
  assign new_n27533_ = ~new_n27534_ & new_n27541_;
  assign new_n27534_ = new_n27535_ & (new_n27539_ | ~new_n27538_);
  assign new_n27535_ = (new_n13168_ | new_n27537_ | new_n18420_) & (~new_n18420_ | (new_n22928_ ? new_n22545_ : ~new_n27536_));
  assign new_n27536_ = (new_n26213_ & new_n18989_) | (~new_n14787_ & ~new_n14810_ & new_n18081_ & ~new_n18989_);
  assign new_n27537_ = (~new_n26343_ | ~new_n26346_ | ~new_n26314_ | ~new_n26338_) & (~new_n21056_ | ~new_n9445_);
  assign new_n27538_ = ~new_n18420_ & new_n13168_;
  assign new_n27539_ = new_n27540_ ? ~new_n26141_ : (new_n17176_ | (new_n17154_ & new_n19313_));
  assign new_n27540_ = ~new_n10240_ & (~new_n10208_ | ~new_n10229_ | ~new_n10238_);
  assign new_n27541_ = new_n27542_ & (~new_n27539_ | ~new_n27538_);
  assign new_n27542_ = (new_n13168_ | ~new_n27537_ | new_n18420_) & (~new_n18420_ | (new_n22928_ ? ~new_n27543_ : new_n27536_));
  assign new_n27543_ = new_n22545_ & new_n25711_;
  assign new_n27544_ = new_n27545_ ? (new_n27557_ ^ new_n27567_) : (~new_n27557_ ^ new_n27567_);
  assign new_n27545_ = ~new_n27546_ & new_n27555_;
  assign new_n27546_ = new_n27547_ & new_n27550_ & (new_n16276_ | ~new_n27554_) & (~new_n27553_ | ~new_n23967_);
  assign new_n27547_ = ~new_n15757_ | (new_n18961_ ? (new_n27549_ ? ~new_n20463_ : ~new_n19605_) : ~new_n27548_);
  assign new_n27548_ = new_n12047_ & new_n22546_ & (~new_n22494_ | ~new_n22467_);
  assign new_n27549_ = ~new_n27187_ & ~new_n15477_;
  assign new_n27550_ = new_n15757_ | (~new_n27551_ & new_n27552_);
  assign new_n27551_ = ~new_n12190_ & new_n14528_ & (new_n14505_ | new_n14530_);
  assign new_n27552_ = new_n20956_ & (new_n20954_ | new_n20924_);
  assign new_n27553_ = new_n15757_ & ~new_n12047_ & ~new_n18961_;
  assign new_n27554_ = new_n27552_ & ~new_n15757_ & new_n12190_;
  assign new_n27555_ = new_n27556_ & (~new_n27554_ | ~new_n16276_);
  assign new_n27556_ = ~new_n15757_ | ((new_n12047_ | new_n23967_ | new_n18961_) & (new_n27549_ | new_n19605_ | ~new_n18961_));
  assign new_n27557_ = ~new_n27558_ & ~new_n27566_;
  assign new_n27558_ = ~new_n27559_ & new_n27562_ & (~new_n14390_ | (new_n27563_ & ~new_n17934_) | (new_n27564_ & new_n17934_));
  assign new_n27559_ = ~new_n14390_ & ~new_n27560_ & (~new_n27561_ | (~new_n18797_ & ~new_n26396_));
  assign new_n27560_ = ~new_n17554_ & ~new_n21692_ & ~new_n27561_;
  assign new_n27561_ = ~new_n6883_ & new_n7950_;
  assign new_n27562_ = new_n14390_ | (~new_n27560_ & (~new_n18797_ | ~new_n27561_ | ~new_n18893_));
  assign new_n27563_ = ~new_n23967_ & new_n24352_;
  assign new_n27564_ = new_n27565_ ? (new_n20436_ | (~new_n24403_ & new_n20408_)) : new_n12798_;
  assign new_n27565_ = new_n12119_ & new_n12141_;
  assign new_n27566_ = new_n27563_ & ~new_n17934_ & new_n14390_;
  assign new_n27567_ = ~new_n27568_ & new_n27576_;
  assign new_n27568_ = (new_n27572_ | new_n27574_ | new_n18582_) & (~new_n18582_ | (new_n27575_ ? new_n27571_ : new_n27569_));
  assign new_n27569_ = (~new_n27570_ | ~new_n17998_ | new_n7126_ | (new_n23081_ & new_n7104_)) & (~new_n11303_ | (~new_n7126_ & (~new_n23081_ | ~new_n7104_)));
  assign new_n27570_ = new_n17976_ & new_n18000_;
  assign new_n27571_ = ~new_n21015_ & (new_n25856_ | ~new_n26092_);
  assign new_n27572_ = new_n20365_ & new_n27573_ & new_n20343_;
  assign new_n27573_ = new_n20371_ & new_n20406_;
  assign new_n27574_ = ~new_n18108_ & ~new_n9163_;
  assign new_n27575_ = new_n23887_ & ~new_n23911_ & ~new_n23915_;
  assign new_n27576_ = ~new_n27577_ & (~new_n18582_ | (~new_n27569_ & ~new_n27575_) | (~new_n27571_ & new_n27575_));
  assign new_n27577_ = ~new_n18582_ & (new_n27574_ | new_n27572_) & (~new_n18739_ | ~new_n17590_ | ~new_n17612_ | ~new_n27572_);
  assign new_n27578_ = ~new_n27579_ & new_n25060_;
  assign new_n27579_ = (~new_n24514_ & ~new_n23184_ & new_n27580_) | (~new_n27580_ & (new_n19766_ ? new_n24401_ : ~new_n25356_));
  assign new_n27580_ = ~new_n14070_ & (~new_n14047_ | new_n15164_);
  assign new_n27581_ = new_n27582_ ? (~new_n27659_ ^ new_n27675_) : (new_n27659_ ^ new_n27675_);
  assign new_n27582_ = new_n27583_ ? (~new_n27647_ ^ new_n27654_) : (new_n27647_ ^ new_n27654_);
  assign new_n27583_ = new_n27584_ ? (~new_n27302_ ^ new_n27640_) : (new_n27302_ ^ new_n27640_);
  assign new_n27584_ = new_n27585_ ? (new_n27596_ ^ new_n27633_) : (~new_n27596_ ^ new_n27633_);
  assign new_n27585_ = ~new_n27586_ & new_n27594_;
  assign new_n27586_ = new_n27587_ & (~new_n27593_ | (~new_n27591_ & new_n27592_) | (~new_n7601_ & ~new_n27592_));
  assign new_n27587_ = new_n27589_ ? ~new_n27590_ : (new_n19046_ ? new_n27588_ : new_n26304_);
  assign new_n27588_ = (new_n12870_ & new_n20233_) | (~new_n6532_ & ~new_n20233_ & (~new_n6529_ | new_n21602_));
  assign new_n27589_ = ~new_n26346_ & (~new_n26343_ | ~new_n26314_);
  assign new_n27590_ = ~new_n17888_ & (~new_n17886_ | ~new_n17877_);
  assign new_n27591_ = ~new_n24388_ & new_n16304_;
  assign new_n27592_ = ~new_n23769_ & (~new_n23766_ | ~new_n24336_);
  assign new_n27593_ = ~new_n27590_ & new_n27589_;
  assign new_n27594_ = ~new_n27595_ & (~new_n27593_ | (new_n27591_ & new_n27592_) | (new_n7601_ & ~new_n27592_));
  assign new_n27595_ = ~new_n27589_ & ((new_n26304_ & ~new_n19046_) | (new_n20233_ & new_n12870_ & new_n19046_));
  assign new_n27596_ = ~new_n27630_ & (new_n10681_ | (new_n27597_ & (new_n11726_ | ~new_n11575_ | ~new_n27598_)));
  assign new_n27597_ = (new_n11575_ | new_n27600_ | ~new_n27598_) & (new_n27599_ | new_n25147_ | new_n27598_);
  assign new_n27598_ = new_n8391_ & (new_n10395_ | new_n10380_);
  assign new_n27599_ = ~new_n21559_ & (~new_n21537_ | new_n25657_);
  assign new_n27600_ = ~new_n27601_ & new_n27628_ & new_n27626_ & (~new_n27629_ | (new_n27622_ & new_n27624_));
  assign new_n27601_ = ~new_n27616_ & (new_n27618_ | (~new_n27619_ & (new_n27620_ | (~new_n27602_ & ~new_n27621_))));
  assign new_n27602_ = ~new_n27606_ & (new_n27608_ | (new_n27615_ & (~new_n27603_ | (~new_n27612_ & new_n27611_))));
  assign new_n27603_ = \all_features[5527]  & (\all_features[5526]  | new_n27604_);
  assign new_n27604_ = \all_features[5525]  & (\all_features[5522]  | \all_features[5523]  | \all_features[5524]  | ~new_n27605_);
  assign new_n27605_ = ~\all_features[5520]  & ~\all_features[5521] ;
  assign new_n27606_ = ~new_n27607_ & ~\all_features[5527] ;
  assign new_n27607_ = \all_features[5525]  & \all_features[5526]  & (\all_features[5524]  | (\all_features[5522]  & \all_features[5523]  & \all_features[5521] ));
  assign new_n27608_ = ~\all_features[5527]  & (~new_n27610_ | ~\all_features[5520]  | ~\all_features[5521]  | ~\all_features[5526]  | ~new_n27609_);
  assign new_n27609_ = \all_features[5524]  & \all_features[5525] ;
  assign new_n27610_ = \all_features[5522]  & \all_features[5523] ;
  assign new_n27611_ = \all_features[5527]  & (\all_features[5526]  | (new_n27609_ & (\all_features[5522]  | \all_features[5523]  | \all_features[5521] )));
  assign new_n27612_ = ~new_n27614_ & ~\all_features[5525]  & new_n27613_ & (~\all_features[5524]  | (~\all_features[5522]  & ~\all_features[5523] ));
  assign new_n27613_ = \all_features[5526]  & \all_features[5527] ;
  assign new_n27614_ = ~\all_features[5522]  & ~\all_features[5523]  & ~\all_features[5524]  & ~\all_features[5525]  & (~\all_features[5521]  | ~\all_features[5520] );
  assign new_n27615_ = \all_features[5527]  & (\all_features[5525]  | \all_features[5526]  | \all_features[5524] );
  assign new_n27616_ = ~\all_features[5525]  & new_n27617_ & ((~\all_features[5522]  & new_n27605_) | ~\all_features[5524]  | ~\all_features[5523] );
  assign new_n27617_ = ~\all_features[5526]  & ~\all_features[5527] ;
  assign new_n27618_ = new_n27617_ & (~\all_features[5525]  | (~\all_features[5524]  & (~\all_features[5523]  | (~\all_features[5522]  & ~\all_features[5521] ))));
  assign new_n27619_ = new_n27617_ & (~new_n27609_ | ~\all_features[5523]  | (~\all_features[5522]  & (~\all_features[5520]  | ~\all_features[5521] )));
  assign new_n27620_ = ~\all_features[5527]  & (~\all_features[5526]  | (~\all_features[5524]  & ~\all_features[5525]  & ~new_n27610_));
  assign new_n27621_ = ~\all_features[5527]  & (~\all_features[5526]  | (~\all_features[5525]  & (new_n27605_ | ~new_n27610_ | ~\all_features[5524] )));
  assign new_n27622_ = new_n27615_ & new_n27623_ & new_n27603_ & new_n27611_;
  assign new_n27623_ = ~new_n27614_ & new_n27613_;
  assign new_n27624_ = new_n27603_ & new_n27615_ & (new_n27625_ | ~new_n27623_ | ~new_n27611_);
  assign new_n27625_ = new_n27613_ & \all_features[5525]  & ((~new_n27605_ & \all_features[5522] ) | \all_features[5524]  | \all_features[5523] );
  assign new_n27626_ = new_n27627_ & ~new_n27606_ & ~new_n27619_ & ~new_n27616_ & ~new_n27618_;
  assign new_n27627_ = ~new_n27608_ & (\all_features[5523]  | \all_features[5524]  | \all_features[5525]  | ~new_n27617_);
  assign new_n27628_ = ~new_n27620_ & ~new_n27621_;
  assign new_n27629_ = ~new_n27606_ & ~new_n27608_;
  assign new_n27630_ = new_n10681_ & ((~new_n27631_ & new_n27632_) | (~new_n16525_ & new_n6568_ & ~new_n27632_));
  assign new_n27631_ = new_n26891_ & ~new_n24259_ & ~new_n24955_;
  assign new_n27632_ = ~new_n12904_ & (~new_n12901_ | new_n16766_);
  assign new_n27633_ = ~new_n27634_ & new_n27637_ & (~new_n23150_ | ~new_n27638_ | new_n24905_ | new_n27636_);
  assign new_n27634_ = new_n27635_ & (new_n25747_ | new_n26997_) & (~new_n27565_ | ~new_n12143_ | ~new_n12147_ | ~new_n26997_);
  assign new_n27635_ = new_n18288_ & new_n18285_ & ~new_n25409_ & new_n27636_;
  assign new_n27636_ = ~new_n21834_ & (~new_n21836_ | ~new_n21809_);
  assign new_n27637_ = new_n27636_ | ((~new_n27639_ | new_n27638_) & (new_n23150_ | new_n25867_ | ~new_n27299_ | ~new_n27638_));
  assign new_n27638_ = ~new_n20342_ & new_n27573_;
  assign new_n27639_ = ~new_n26422_ & ~new_n15596_ & (~new_n26424_ | ~new_n26404_);
  assign new_n27640_ = new_n27641_ & (new_n21355_ ? ~new_n27645_ : (~new_n27646_ | (~new_n19764_ & new_n20846_)));
  assign new_n27641_ = ~new_n27642_ & (new_n21355_ | new_n6532_ | ~new_n27644_ | (new_n6529_ & new_n6498_));
  assign new_n27642_ = ~new_n23922_ & new_n27643_ & new_n21355_ & (new_n18000_ | ~new_n17975_);
  assign new_n27643_ = new_n21125_ & new_n21111_ & (new_n25619_ | (new_n21120_ & new_n21132_));
  assign new_n27644_ = new_n6568_ & new_n6597_;
  assign new_n27645_ = new_n8630_ & ~new_n24335_ & ~new_n27643_;
  assign new_n27646_ = ~new_n27644_ & new_n13556_ & new_n19766_ & (new_n13553_ | new_n13545_);
  assign new_n27647_ = new_n27648_ & (new_n10681_ ? new_n27652_ : (new_n27653_ | (new_n24009_ & new_n25936_)));
  assign new_n27648_ = ~new_n27649_ & ~new_n27650_ & (new_n23665_ | new_n12900_ | new_n14042_ | ~new_n10681_);
  assign new_n27649_ = new_n10681_ & new_n12900_ & ~new_n8854_ & ~new_n24395_ & ~new_n22949_;
  assign new_n27650_ = ~new_n10681_ & new_n27651_ & ((~new_n23583_ & new_n23823_) ? new_n13063_ : ~new_n8506_);
  assign new_n27651_ = new_n24009_ & new_n25936_;
  assign new_n27652_ = (new_n26390_ | ~new_n14042_ | new_n12900_) & (~new_n24395_ | ~new_n12900_ | (new_n10243_ & new_n6736_));
  assign new_n27653_ = (new_n19702_ & new_n21694_ & (new_n19679_ | ~new_n19720_)) | (~new_n24451_ & ~new_n21694_);
  assign new_n27654_ = new_n24395_ ? new_n27657_ : (new_n27655_ & (new_n26876_ | ~new_n24143_ | ~new_n27656_));
  assign new_n27655_ = (~new_n9725_ | ~new_n20570_ | ~new_n26876_) & (new_n27656_ | new_n11608_ | new_n26876_);
  assign new_n27656_ = ~new_n7251_ & (~new_n7229_ | ~new_n26902_);
  assign new_n27657_ = (new_n21012_ | new_n11169_ | ~new_n27658_) & (~new_n26777_ | ~new_n12980_ | new_n27658_);
  assign new_n27658_ = ~new_n10682_ & (~new_n13937_ | ~new_n24180_);
  assign new_n27659_ = ~new_n27660_ & new_n27673_;
  assign new_n27660_ = new_n27661_ & ((new_n25277_ & new_n27672_ & new_n27671_) | (new_n27665_ & new_n27664_));
  assign new_n27661_ = new_n27662_ & (~new_n27671_ | (new_n19846_ & ~new_n27672_) | (new_n25277_ & new_n27672_));
  assign new_n27662_ = (~new_n27667_ | ~new_n27666_) & (~new_n27669_ | ~new_n27668_) & (new_n27670_ | ~new_n27663_);
  assign new_n27663_ = ~new_n27665_ & new_n27664_;
  assign new_n27664_ = ~new_n21355_ & new_n25711_;
  assign new_n27665_ = ~new_n22872_ & (~new_n22874_ | new_n23162_);
  assign new_n27666_ = new_n21355_ & new_n25711_;
  assign new_n27667_ = (~new_n24516_ & ~new_n27188_) | (new_n9134_ & new_n24342_ & new_n27188_);
  assign new_n27668_ = new_n12908_ & ~new_n25711_ & new_n20845_;
  assign new_n27669_ = new_n23336_ & new_n17961_;
  assign new_n27670_ = ~new_n25386_ & new_n23200_;
  assign new_n27671_ = ~new_n12908_ & ~new_n25711_;
  assign new_n27672_ = ~new_n25668_ & new_n26163_;
  assign new_n27673_ = new_n27674_ & (new_n27669_ | ~new_n27668_) & (~new_n27666_ | new_n27667_);
  assign new_n27674_ = (new_n27672_ | ~new_n19846_ | ~new_n27671_) & (~new_n27670_ | ~new_n27663_);
  assign new_n27675_ = ~new_n27308_ & new_n27304_;
  assign new_n27676_ = ~new_n27677_ & new_n27684_;
  assign new_n27677_ = new_n27678_ & (~new_n18582_ | (~new_n27683_ & ~new_n18740_) | (new_n16233_ & new_n13134_ & new_n18740_));
  assign new_n27678_ = (~new_n27682_ | ~new_n27680_) & (~new_n27679_ | (new_n27681_ ? ~new_n10603_ : ~new_n9163_));
  assign new_n27679_ = ~new_n24178_ & ~new_n18582_;
  assign new_n27680_ = new_n18015_ & ~new_n18740_ & new_n18582_;
  assign new_n27681_ = ~new_n12865_ & new_n11940_;
  assign new_n27682_ = new_n16378_ & new_n16400_;
  assign new_n27683_ = new_n7558_ & ~new_n14391_ & ~new_n18015_;
  assign new_n27684_ = new_n27685_ & (new_n27686_ | new_n18582_) & (~new_n13134_ | ~new_n16233_ | ~new_n18740_ | ~new_n18582_);
  assign new_n27685_ = (~new_n27680_ | new_n27682_) & (new_n27681_ | new_n9163_ | ~new_n27679_);
  assign new_n27686_ = (~new_n24178_ & (new_n10603_ | ~new_n27681_)) | (new_n15874_ & new_n24401_ & new_n24178_);
  assign new_n27687_ = ~new_n27699_ & new_n27688_;
  assign new_n27688_ = new_n27689_ & (new_n27698_ | ~new_n27697_) & (~new_n27696_ | new_n10637_);
  assign new_n27689_ = ~new_n27690_ & (new_n27692_ | (new_n27695_ & new_n16776_) | (~new_n27694_ & ~new_n16776_));
  assign new_n27690_ = ~new_n17998_ & ~new_n20786_ & new_n27691_ & (~new_n18004_ | ~new_n27570_);
  assign new_n27691_ = ~new_n27693_ & new_n27692_;
  assign new_n27692_ = new_n12184_ & new_n16566_;
  assign new_n27693_ = ~new_n15786_ & (~new_n15763_ | ~new_n15788_);
  assign new_n27694_ = ~new_n25807_ & ~new_n21641_;
  assign new_n27695_ = new_n26730_ ? new_n16850_ : ~new_n16758_;
  assign new_n27696_ = new_n27691_ & new_n20786_;
  assign new_n27697_ = new_n27692_ & new_n27693_;
  assign new_n27698_ = (~new_n17770_ & ~new_n17800_ & ~new_n17802_) ? (new_n13735_ | new_n13765_) : new_n17588_;
  assign new_n27699_ = new_n27700_ & (~new_n10637_ | ~new_n27696_) & (~new_n27698_ | ~new_n27697_);
  assign new_n27700_ = new_n27692_ | (new_n16776_ ? (new_n26730_ ? ~new_n16850_ : new_n16758_) : new_n27694_);
  assign new_n27701_ = ~new_n27702_ & new_n27710_;
  assign new_n27702_ = new_n27703_ & (~new_n13349_ | (~new_n27708_ & (new_n27709_ | ~new_n12849_ | ~new_n7097_)));
  assign new_n27703_ = (~new_n27707_ | new_n27704_ | new_n13349_) & (new_n27706_ | new_n7097_ | new_n27705_ | ~new_n13349_);
  assign new_n27704_ = new_n12562_ ? new_n26768_ : new_n14070_;
  assign new_n27705_ = new_n25709_ & ~new_n26643_ & ~new_n20377_;
  assign new_n27706_ = new_n17631_ & (~new_n12855_ | ~new_n12851_);
  assign new_n27707_ = ~new_n21111_ & (~new_n25619_ | ~new_n25615_);
  assign new_n27708_ = ~new_n7097_ & new_n27705_ & (~new_n10333_ | (~new_n10311_ & ~new_n10339_));
  assign new_n27709_ = ~new_n21852_ & ~new_n6388_;
  assign new_n27710_ = new_n27711_ & (new_n13349_ | (~new_n27704_ & new_n27707_) | (new_n27713_ & ~new_n27707_));
  assign new_n27711_ = ~new_n13349_ | (~new_n27712_ & (~new_n7097_ | (new_n12849_ ? ~new_n27709_ : ~new_n22545_)));
  assign new_n27712_ = new_n27706_ & ~new_n27705_ & ~new_n7097_;
  assign new_n27713_ = (~new_n15214_ & ~new_n15264_) ? ~new_n27439_ : (~new_n10833_ | (~new_n10830_ & new_n24953_));
  assign new_n27714_ = new_n27202_ ? new_n27715_ : ((~new_n21201_ & new_n22036_ & ~new_n27201_) | (new_n27718_ & new_n27201_));
  assign new_n27715_ = (new_n27716_ | new_n17455_) & (new_n21706_ | new_n27717_ | new_n20693_ | ~new_n17455_);
  assign new_n27716_ = new_n25861_ & new_n26092_ & new_n25857_;
  assign new_n27717_ = new_n20689_ & new_n20662_ & new_n20684_;
  assign new_n27718_ = ~new_n19813_ & new_n12904_ & (new_n12901_ | new_n12871_);
  assign \o[64]  = new_n27720_ ^ new_n27721_;
  assign new_n27720_ = new_n27161_ & new_n27714_;
  assign new_n27721_ = new_n27722_ ? (new_n27723_ ^ new_n27775_) : (~new_n27723_ ^ new_n27775_);
  assign new_n27722_ = (new_n27687_ & new_n27701_) | (~new_n27162_ & (new_n27687_ | new_n27701_));
  assign new_n27723_ = new_n27724_ ? (~new_n27725_ ^ new_n27774_) : (new_n27725_ ^ new_n27774_);
  assign new_n27724_ = (~new_n27581_ & new_n27676_) | (~new_n27163_ & (~new_n27581_ | new_n27676_));
  assign new_n27725_ = new_n27726_ ? (new_n27727_ ^ new_n27761_) : (~new_n27727_ ^ new_n27761_);
  assign new_n27726_ = (~new_n27343_ & new_n27578_) | (~new_n27164_ & (~new_n27343_ | new_n27578_));
  assign new_n27727_ = new_n27728_ ? (new_n27741_ ^ new_n27742_) : (~new_n27741_ ^ new_n27742_);
  assign new_n27728_ = new_n27729_ ? (~new_n27730_ ^ new_n27740_) : (new_n27730_ ^ new_n27740_);
  assign new_n27729_ = (~new_n27196_ & new_n27302_) | (~new_n27166_ & (~new_n27196_ | new_n27302_));
  assign new_n27730_ = new_n27731_ ? (new_n27735_ ^ new_n27739_) : (~new_n27735_ ^ new_n27739_);
  assign new_n27731_ = new_n27732_ ? (new_n27733_ ^ new_n27734_) : (~new_n27733_ ^ new_n27734_);
  assign new_n27732_ = new_n27347_ & new_n27367_;
  assign new_n27733_ = new_n27372_ & new_n27377_;
  assign new_n27734_ = new_n27198_ & new_n27238_;
  assign new_n27735_ = new_n27736_ ? (new_n27737_ ^ new_n27738_) : (~new_n27737_ ^ new_n27738_);
  assign new_n27736_ = new_n27661_ & new_n27673_;
  assign new_n27737_ = ~new_n27566_ & new_n27558_;
  assign new_n27738_ = ~new_n27380_ & (new_n27384_ | ~new_n24077_ | new_n24023_) & (~new_n16026_ | new_n19147_ | ~new_n24023_);
  assign new_n27739_ = (new_n27242_ & new_n27254_) | (new_n27197_ & (new_n27242_ | new_n27254_));
  assign new_n27740_ = (new_n27386_ & new_n27427_) | (~new_n27345_ & (new_n27386_ | new_n27427_));
  assign new_n27741_ = (~new_n27428_ & new_n27303_) | (~new_n27344_ & (~new_n27428_ | new_n27303_));
  assign new_n27742_ = new_n27743_ ? (new_n27750_ ^ new_n27751_) : (~new_n27750_ ^ new_n27751_);
  assign new_n27743_ = new_n27744_ ? (~new_n27745_ ^ new_n27749_) : (new_n27745_ ^ new_n27749_);
  assign new_n27744_ = (~new_n27378_ & new_n27371_) | (new_n27346_ & (~new_n27378_ | new_n27371_));
  assign new_n27745_ = new_n27746_ ? (new_n27747_ ^ new_n27748_) : (~new_n27747_ ^ new_n27748_);
  assign new_n27746_ = new_n27546_ & new_n27555_;
  assign new_n27747_ = new_n27677_ & new_n27684_;
  assign new_n27748_ = new_n27568_ & new_n27576_;
  assign new_n27749_ = (new_n27557_ & new_n27567_) | (new_n27545_ & (new_n27557_ | new_n27567_));
  assign new_n27750_ = (~new_n27544_ & new_n27427_) | (~new_n27429_ & (~new_n27544_ | new_n27427_));
  assign new_n27751_ = new_n27752_ ? (new_n27753_ ^ new_n27757_) : (~new_n27753_ ^ new_n27757_);
  assign new_n27752_ = (new_n27453_ & new_n27533_) | (new_n27430_ & (new_n27453_ | new_n27533_));
  assign new_n27753_ = new_n27754_ ^ new_n27755_;
  assign new_n27754_ = new_n27431_ & new_n27451_;
  assign new_n27755_ = new_n27500_ & ~new_n27756_ & new_n27454_;
  assign new_n27756_ = ~new_n27494_ & new_n27495_;
  assign new_n27757_ = new_n27758_ ? (new_n27759_ ^ new_n27760_) : (~new_n27759_ ^ new_n27760_);
  assign new_n27758_ = new_n27688_ & new_n27699_;
  assign new_n27759_ = new_n27534_ & new_n27541_;
  assign new_n27760_ = new_n27702_ & new_n27710_;
  assign new_n27761_ = new_n27762_ ? (~new_n27772_ ^ new_n27773_) : (new_n27772_ ^ new_n27773_);
  assign new_n27762_ = new_n27763_ ? (~new_n27770_ ^ new_n27771_) : (new_n27770_ ^ new_n27771_);
  assign new_n27763_ = new_n27764_ ? (~new_n27768_ ^ new_n27769_) : (new_n27768_ ^ new_n27769_);
  assign new_n27764_ = new_n27765_ ? (new_n27766_ ^ new_n27767_) : (~new_n27766_ ^ new_n27767_);
  assign new_n27765_ = new_n27168_ & new_n27178_;
  assign new_n27766_ = new_n27312_ & new_n27341_;
  assign new_n27767_ = new_n27255_ & new_n27300_;
  assign new_n27768_ = (new_n27181_ & new_n27191_) | (new_n27167_ & (new_n27181_ | new_n27191_));
  assign new_n27769_ = (new_n27596_ & new_n27633_) | (new_n27585_ & (new_n27596_ | new_n27633_));
  assign new_n27770_ = (new_n27302_ & new_n27640_) | (~new_n27584_ & (new_n27302_ | new_n27640_));
  assign new_n27771_ = new_n27586_ & new_n27594_;
  assign new_n27772_ = (new_n27303_ & new_n27311_) | (~new_n27165_ & (new_n27303_ | new_n27311_));
  assign new_n27773_ = (new_n27647_ & new_n27654_) | (~new_n27583_ & (new_n27647_ | new_n27654_));
  assign new_n27774_ = (new_n27659_ & new_n27675_) | (~new_n27582_ & (new_n27659_ | new_n27675_));
  assign new_n27775_ = new_n27387_ & new_n27426_;
  assign \o[65]  = ~new_n27777_ ^ new_n27778_;
  assign new_n27777_ = new_n27720_ & new_n27721_;
  assign new_n27778_ = new_n27779_ ^ new_n27780_;
  assign new_n27779_ = (~new_n27723_ & new_n27775_) | (new_n27722_ & (~new_n27723_ | new_n27775_));
  assign new_n27780_ = ~new_n27781_ ^ new_n27782_;
  assign new_n27781_ = (~new_n27725_ & new_n27774_) | (new_n27724_ & (~new_n27725_ | new_n27774_));
  assign new_n27782_ = new_n27783_ ? (new_n27784_ ^ new_n27810_) : (~new_n27784_ ^ new_n27810_);
  assign new_n27783_ = (~new_n27727_ & ~new_n27761_) | (new_n27726_ & (~new_n27727_ | ~new_n27761_));
  assign new_n27784_ = new_n27785_ ? (new_n27793_ ^ new_n27794_) : (~new_n27793_ ^ new_n27794_);
  assign new_n27785_ = new_n27786_ ? (~new_n27791_ ^ new_n27792_) : (new_n27791_ ^ new_n27792_);
  assign new_n27786_ = ~new_n27787_ ^ new_n27790_;
  assign new_n27787_ = new_n27788_ ^ new_n27789_;
  assign new_n27788_ = (new_n27766_ & new_n27767_) | (new_n27765_ & (new_n27766_ | new_n27767_));
  assign new_n27789_ = (new_n27733_ & new_n27734_) | (new_n27732_ & (new_n27733_ | new_n27734_));
  assign new_n27790_ = (new_n27768_ & new_n27769_) | (~new_n27764_ & (new_n27768_ | new_n27769_));
  assign new_n27791_ = (~new_n27730_ & new_n27740_) | (new_n27729_ & (~new_n27730_ | new_n27740_));
  assign new_n27792_ = (new_n27770_ & new_n27771_) | (~new_n27763_ & (new_n27770_ | new_n27771_));
  assign new_n27793_ = (~new_n27742_ & new_n27741_) | (~new_n27728_ & (~new_n27742_ | new_n27741_));
  assign new_n27794_ = new_n27795_ ? (new_n27799_ ^ new_n27800_) : (~new_n27799_ ^ new_n27800_);
  assign new_n27795_ = new_n27796_ ? (new_n27797_ ^ new_n27798_) : (~new_n27797_ ^ new_n27798_);
  assign new_n27796_ = (~new_n27735_ & new_n27739_) | (~new_n27731_ & (~new_n27735_ | new_n27739_));
  assign new_n27797_ = (~new_n27745_ & new_n27749_) | (new_n27744_ & (~new_n27745_ | new_n27749_));
  assign new_n27798_ = (new_n27737_ & new_n27738_) | (new_n27736_ & (new_n27737_ | new_n27738_));
  assign new_n27799_ = (~new_n27751_ & new_n27750_) | (~new_n27743_ & (~new_n27751_ | new_n27750_));
  assign new_n27800_ = new_n27801_ ? (new_n27802_ ^ new_n27807_) : (~new_n27802_ ^ new_n27807_);
  assign new_n27801_ = (~new_n27753_ & ~new_n27757_) | (new_n27752_ & (~new_n27753_ | ~new_n27757_));
  assign new_n27802_ = ~new_n27803_ ^ new_n27804_;
  assign new_n27803_ = ~new_n27754_ & ~new_n27755_;
  assign new_n27804_ = ~new_n27805_ ^ new_n27806_;
  assign new_n27805_ = new_n27500_ & new_n27454_ & new_n27756_;
  assign new_n27806_ = new_n27451_ & new_n27432_ & new_n27448_;
  assign new_n27807_ = ~new_n27808_ ^ new_n27809_;
  assign new_n27808_ = (new_n27747_ & new_n27748_) | (new_n27746_ & (new_n27747_ | new_n27748_));
  assign new_n27809_ = (new_n27759_ & new_n27760_) | (new_n27758_ & (new_n27759_ | new_n27760_));
  assign new_n27810_ = (new_n27772_ & new_n27773_) | (~new_n27762_ & (new_n27772_ | new_n27773_));
  assign \o[66]  = ((new_n27812_ | new_n27813_) & (new_n27814_ ^ new_n27815_)) | (~new_n27812_ & ~new_n27813_ & (~new_n27814_ ^ new_n27815_));
  assign new_n27812_ = ~new_n27778_ & new_n27777_;
  assign new_n27813_ = ~new_n27780_ & new_n27779_;
  assign new_n27814_ = new_n27781_ & new_n27782_;
  assign new_n27815_ = ~new_n27816_ ^ new_n27817_;
  assign new_n27816_ = (~new_n27784_ & new_n27810_) | (new_n27783_ & (~new_n27784_ | new_n27810_));
  assign new_n27817_ = new_n27818_ ? (new_n27819_ ^ new_n27831_) : (~new_n27819_ ^ new_n27831_);
  assign new_n27818_ = (~new_n27794_ & new_n27793_) | (~new_n27785_ & (~new_n27794_ | new_n27793_));
  assign new_n27819_ = new_n27820_ ? (new_n27824_ ^ new_n27825_) : (~new_n27824_ ^ new_n27825_);
  assign new_n27820_ = new_n27821_ ? (new_n27822_ ^ new_n27823_) : (~new_n27822_ ^ new_n27823_);
  assign new_n27821_ = new_n27787_ & new_n27790_;
  assign new_n27822_ = new_n27788_ & new_n27789_;
  assign new_n27823_ = (new_n27797_ & new_n27798_) | (new_n27796_ & (new_n27797_ | new_n27798_));
  assign new_n27824_ = (~new_n27800_ & new_n27799_) | (~new_n27795_ & (~new_n27800_ | new_n27799_));
  assign new_n27825_ = new_n27826_ ? (~new_n27827_ ^ new_n27830_) : (new_n27827_ ^ new_n27830_);
  assign new_n27826_ = (~new_n27802_ & ~new_n27807_) | (new_n27801_ & (~new_n27802_ | ~new_n27807_));
  assign new_n27827_ = ~new_n27828_ ^ new_n27829_;
  assign new_n27828_ = ~new_n27803_ & ~new_n27804_;
  assign new_n27829_ = new_n27805_ & new_n27806_;
  assign new_n27830_ = new_n27808_ & new_n27809_;
  assign new_n27831_ = (new_n27791_ & new_n27792_) | (~new_n27786_ & (new_n27791_ | new_n27792_));
  assign \o[67]  = ~new_n27833_ ^ new_n27834_;
  assign new_n27833_ = (new_n27814_ | (~new_n27815_ & (new_n27813_ | new_n27812_))) & (new_n27813_ | new_n27812_ | ~new_n27815_);
  assign new_n27834_ = new_n27835_ ^ new_n27836_;
  assign new_n27835_ = new_n27816_ & new_n27817_;
  assign new_n27836_ = ~new_n27837_ ^ new_n27838_;
  assign new_n27837_ = (~new_n27819_ & new_n27831_) | (new_n27818_ & (~new_n27819_ | new_n27831_));
  assign new_n27838_ = new_n27839_ ? (new_n27840_ ^ new_n27841_) : (~new_n27840_ ^ new_n27841_);
  assign new_n27839_ = (~new_n27825_ & new_n27824_) | (~new_n27820_ & (~new_n27825_ | new_n27824_));
  assign new_n27840_ = (new_n27822_ & new_n27823_) | (new_n27821_ & (new_n27822_ | new_n27823_));
  assign new_n27841_ = ~new_n27842_ ^ new_n27843_;
  assign new_n27842_ = (~new_n27827_ & new_n27830_) | (new_n27826_ & (~new_n27827_ | new_n27830_));
  assign new_n27843_ = new_n27828_ & new_n27829_;
  assign \o[68]  = ((new_n27848_ ^ new_n27849_) & ((~new_n27845_ & ~new_n27846_ & ~new_n27847_) | (new_n27847_ & (new_n27845_ | new_n27846_)))) | (((~new_n27847_ & (new_n27845_ | new_n27846_)) | (~new_n27845_ & ~new_n27846_ & new_n27847_)) & (new_n27848_ ^ ~new_n27849_));
  assign new_n27845_ = ~new_n27834_ & new_n27833_;
  assign new_n27846_ = ~new_n27836_ & new_n27835_;
  assign new_n27847_ = new_n27837_ & new_n27838_;
  assign new_n27848_ = (~new_n27841_ & new_n27840_) | (new_n27839_ & (~new_n27841_ | new_n27840_));
  assign new_n27849_ = new_n27842_ & new_n27843_;
  assign \o[69]  = (~new_n27847_ | ~new_n27848_ | ~new_n27849_ | (~new_n27845_ & ~new_n27846_)) & (new_n27847_ | new_n27848_ | new_n27849_) & (new_n27845_ | new_n27846_ | ((new_n27848_ | new_n27849_) & (new_n27847_ | (new_n27848_ & new_n27849_))));
endmodule


