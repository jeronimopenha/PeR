// Benchmark "TreeLUT" written by ABC on Fri Sep  5 17:00:20 2025

module TreeLUT ( 
    \i[0] , \i[1] , \i[2] , \i[3] , \i[4] , \i[5] , \i[6] , \i[7] , \i[8] ,
    \i[9] , \i[10] , \i[11] , \i[12] , \i[13] , \i[14] , \i[15] , \i[16] ,
    \i[17] , \i[18] , \i[19] , \i[20] , \i[21] , \i[22] , \i[23] , \i[24] ,
    \i[25] , \i[26] , \i[27] , \i[28] , \i[29] , \i[30] , \i[31] , \i[32] ,
    \i[33] , \i[34] , \i[35] , \i[36] , \i[37] , \i[38] , \i[39] , \i[40] ,
    \i[41] , \i[42] , \i[43] , \i[44] , \i[45] , \i[46] , \i[47] , \i[48] ,
    \i[49] , \i[50] , \i[51] , \i[52] , \i[53] , \i[54] , \i[55] , \i[56] ,
    \i[57] , \i[58] , \i[59] , \i[60] , \i[61] , \i[62] , \i[63] , \i[64] ,
    \i[65] , \i[66] , \i[67] , \i[68] , \i[69] , \i[70] , \i[71] , \i[72] ,
    \i[73] , \i[74] , \i[75] , \i[76] , \i[77] , \i[78] , \i[79] , \i[80] ,
    \i[81] , \i[82] , \i[83] , \i[84] , \i[85] , \i[86] , \i[87] , \i[88] ,
    \i[89] , \i[90] , \i[91] , \i[92] , \i[93] , \i[94] , \i[95] , \i[96] ,
    \i[97] , \i[98] , \i[99] , \i[100] , \i[101] , \i[102] , \i[103] ,
    \i[104] , \i[105] , \i[106] , \i[107] , \i[108] , \i[109] , \i[110] ,
    \i[111] , \i[112] , \i[113] , \i[114] , \i[115] , \i[116] , \i[117] ,
    \i[118] , \i[119] , \i[120] , \i[121] , \i[122] , \i[123] , \i[124] ,
    \i[125] , \i[126] , \i[127] , \i[128] , \i[129] , \i[130] , \i[131] ,
    \i[132] , \i[133] , \i[134] , \i[135] , \i[136] , \i[137] , \i[138] ,
    \i[139] , \i[140] , \i[141] , \i[142] , \i[143] , \i[144] , \i[145] ,
    \i[146] , \i[147] , \i[148] , \i[149] , \i[150] , \i[151] , \i[152] ,
    \i[153] , \i[154] , \i[155] , \i[156] , \i[157] , \i[158] , \i[159] ,
    \i[160] , \i[161] , \i[162] , \i[163] , \i[164] , \i[165] , \i[166] ,
    \i[167] , \i[168] , \i[169] , \i[170] , \i[171] , \i[172] , \i[173] ,
    \i[174] , \i[175] , \i[176] , \i[177] , \i[178] , \i[179] , \i[180] ,
    \i[181] , \i[182] , \i[183] , \i[184] , \i[185] , \i[186] , \i[187] ,
    \i[188] , \i[189] , \i[190] , \i[191] , \i[192] , \i[193] , \i[194] ,
    \i[195] , \i[196] , \i[197] , \i[198] , \i[199] , \i[200] , \i[201] ,
    \i[202] , \i[203] , \i[204] , \i[205] , \i[206] , \i[207] , \i[208] ,
    \i[209] , \i[210] , \i[211] , \i[212] , \i[213] , \i[214] , \i[215] ,
    \i[216] , \i[217] , \i[218] , \i[219] , \i[220] , \i[221] , \i[222] ,
    \i[223] , \i[224] , \i[225] , \i[226] , \i[227] , \i[228] , \i[229] ,
    \i[230] , \i[231] , \i[232] , \i[233] , \i[234] , \i[235] , \i[236] ,
    \i[237] , \i[238] , \i[239] , \i[240] , \i[241] , \i[242] , \i[243] ,
    \i[244] , \i[245] , \i[246] , \i[247] , \i[248] , \i[249] , \i[250] ,
    \i[251] , \i[252] , \i[253] , \i[254] , \i[255] , \i[256] , \i[257] ,
    \i[258] , \i[259] , \i[260] , \i[261] , \i[262] , \i[263] , \i[264] ,
    \i[265] , \i[266] , \i[267] , \i[268] , \i[269] , \i[270] , \i[271] ,
    \i[272] , \i[273] , \i[274] , \i[275] , \i[276] , \i[277] , \i[278] ,
    \i[279] , \i[280] , \i[281] , \i[282] , \i[283] , \i[284] , \i[285] ,
    \i[286] , \i[287] , \i[288] , \i[289] , \i[290] , \i[291] , \i[292] ,
    \i[293] , \i[294] , \i[295] , \i[296] , \i[297] , \i[298] , \i[299] ,
    \i[300] , \i[301] , \i[302] , \i[303] , \i[304] , \i[305] , \i[306] ,
    \i[307] , \i[308] , \i[309] , \i[310] , \i[311] , \i[312] , \i[313] ,
    \i[314] , \i[315] , \i[316] , \i[317] , \i[318] , \i[319] , \i[320] ,
    \i[321] , \i[322] , \i[323] , \i[324] , \i[325] , \i[326] , \i[327] ,
    \i[328] , \i[329] , \i[330] , \i[331] , \i[332] , \i[333] , \i[334] ,
    \i[335] , \i[336] , \i[337] , \i[338] , \i[339] , \i[340] , \i[341] ,
    \i[342] , \i[343] , \i[344] , \i[345] , \i[346] , \i[347] , \i[348] ,
    \i[349] , \i[350] , \i[351] , \i[352] , \i[353] , \i[354] , \i[355] ,
    \i[356] , \i[357] , \i[358] , \i[359] , \i[360] , \i[361] , \i[362] ,
    \i[363] , \i[364] , \i[365] , \i[366] , \i[367] , \i[368] , \i[369] ,
    \i[370] , \i[371] , \i[372] , \i[373] , \i[374] , \i[375] , \i[376] ,
    \i[377] , \i[378] , \i[379] , \i[380] , \i[381] , \i[382] , \i[383] ,
    \i[384] , \i[385] , \i[386] , \i[387] , \i[388] , \i[389] , \i[390] ,
    \i[391] , \i[392] , \i[393] , \i[394] , \i[395] , \i[396] , \i[397] ,
    \i[398] , \i[399] , \i[400] , \i[401] , \i[402] , \i[403] , \i[404] ,
    \i[405] , \i[406] , \i[407] , \i[408] , \i[409] , \i[410] , \i[411] ,
    \i[412] , \i[413] , \i[414] , \i[415] , \i[416] , \i[417] , \i[418] ,
    \i[419] , \i[420] , \i[421] , \i[422] , \i[423] , \i[424] , \i[425] ,
    \i[426] , \i[427] , \i[428] , \i[429] , \i[430] , \i[431] , \i[432] ,
    \i[433] , \i[434] , \i[435] , \i[436] , \i[437] , \i[438] , \i[439] ,
    \i[440] , \i[441] , \i[442] , \i[443] , \i[444] , \i[445] , \i[446] ,
    \i[447] , \i[448] , \i[449] , \i[450] , \i[451] , \i[452] , \i[453] ,
    \i[454] , \i[455] , \i[456] , \i[457] , \i[458] , \i[459] , \i[460] ,
    \i[461] , \i[462] , \i[463] , \i[464] , \i[465] , \i[466] , \i[467] ,
    \i[468] , \i[469] , \i[470] , \i[471] , \i[472] , \i[473] , \i[474] ,
    \i[475] , \i[476] , \i[477] , \i[478] , \i[479] , \i[480] , \i[481] ,
    \i[482] , \i[483] , \i[484] , \i[485] , \i[486] , \i[487] , \i[488] ,
    \i[489] , \i[490] , \i[491] , \i[492] , \i[493] , \i[494] , \i[495] ,
    \i[496] , \i[497] , \i[498] , \i[499] , \i[500] , \i[501] , \i[502] ,
    \i[503] , \i[504] , \i[505] , \i[506] , \i[507] , \i[508] , \i[509] ,
    \i[510] , \i[511] , \i[512] , \i[513] , \i[514] , \i[515] , \i[516] ,
    \i[517] , \i[518] , \i[519] , \i[520] , \i[521] , \i[522] , \i[523] ,
    \i[524] , \i[525] , \i[526] , \i[527] , \i[528] , \i[529] , \i[530] ,
    \i[531] , \i[532] , \i[533] , \i[534] , \i[535] , \i[536] , \i[537] ,
    \i[538] , \i[539] , \i[540] , \i[541] , \i[542] , \i[543] , \i[544] ,
    \i[545] , \i[546] , \i[547] , \i[548] , \i[549] , \i[550] , \i[551] ,
    \i[552] , \i[553] , \i[554] , \i[555] , \i[556] , \i[557] , \i[558] ,
    \i[559] , \i[560] , \i[561] , \i[562] , \i[563] , \i[564] , \i[565] ,
    \i[566] , \i[567] , \i[568] , \i[569] , \i[570] , \i[571] , \i[572] ,
    \i[573] , \i[574] , \i[575] , \i[576] , \i[577] , \i[578] , \i[579] ,
    \i[580] , \i[581] , \i[582] , \i[583] , \i[584] , \i[585] , \i[586] ,
    \i[587] , \i[588] , \i[589] , \i[590] , \i[591] , \i[592] , \i[593] ,
    \i[594] , \i[595] , \i[596] , \i[597] , \i[598] , \i[599] , \i[600] ,
    \i[601] , \i[602] , \i[603] , \i[604] , \i[605] , \i[606] , \i[607] ,
    \i[608] , \i[609] , \i[610] , \i[611] , \i[612] , \i[613] , \i[614] ,
    \i[615] , \i[616] , \i[617] , \i[618] , \i[619] , \i[620] , \i[621] ,
    \i[622] , \i[623] , \i[624] , \i[625] , \i[626] , \i[627] , \i[628] ,
    \i[629] , \i[630] , \i[631] , \i[632] , \i[633] , \i[634] , \i[635] ,
    \i[636] , \i[637] , \i[638] , \i[639] , \i[640] , \i[641] , \i[642] ,
    \i[643] , \i[644] , \i[645] , \i[646] , \i[647] , \i[648] , \i[649] ,
    \i[650] , \i[651] , \i[652] , \i[653] , \i[654] , \i[655] , \i[656] ,
    \i[657] , \i[658] , \i[659] , \i[660] , \i[661] , \i[662] , \i[663] ,
    \i[664] , \i[665] , \i[666] , \i[667] , \i[668] , \i[669] , \i[670] ,
    \i[671] , \i[672] , \i[673] , \i[674] , \i[675] , \i[676] , \i[677] ,
    \i[678] , \i[679] , \i[680] , \i[681] , \i[682] , \i[683] , \i[684] ,
    \i[685] , \i[686] , \i[687] , \i[688] , \i[689] , \i[690] , \i[691] ,
    \i[692] , \i[693] , \i[694] , \i[695] , \i[696] , \i[697] , \i[698] ,
    \i[699] , \i[700] , \i[701] , \i[702] , \i[703] , \i[704] , \i[705] ,
    \i[706] , \i[707] , \i[708] , \i[709] , \i[710] , \i[711] , \i[712] ,
    \i[713] , \i[714] , \i[715] , \i[716] , \i[717] , \i[718] , \i[719] ,
    \i[720] , \i[721] , \i[722] , \i[723] , \i[724] , \i[725] , \i[726] ,
    \i[727] , \i[728] , \i[729] , \i[730] , \i[731] , \i[732] , \i[733] ,
    \i[734] , \i[735] , \i[736] , \i[737] , \i[738] , \i[739] , \i[740] ,
    \i[741] , \i[742] , \i[743] , \i[744] , \i[745] , \i[746] , \i[747] ,
    \i[748] , \i[749] , \i[750] , \i[751] , \i[752] , \i[753] , \i[754] ,
    \i[755] , \i[756] , \i[757] , \i[758] , \i[759] , \i[760] , \i[761] ,
    \i[762] , \i[763] , \i[764] , \i[765] , \i[766] , \i[767] , \i[768] ,
    \i[769] , \i[770] , \i[771] , \i[772] , \i[773] , \i[774] , \i[775] ,
    \i[776] , \i[777] , \i[778] , \i[779] , \i[780] , \i[781] , \i[782] ,
    \i[783] , \i[784] , \i[785] , \i[786] , \i[787] , \i[788] , \i[789] ,
    \i[790] , \i[791] , \i[792] , \i[793] , \i[794] , \i[795] , \i[796] ,
    \i[797] , \i[798] , \i[799] , \i[800] , \i[801] , \i[802] , \i[803] ,
    \i[804] , \i[805] , \i[806] , \i[807] , \i[808] , \i[809] , \i[810] ,
    \i[811] , \i[812] , \i[813] , \i[814] , \i[815] , \i[816] , \i[817] ,
    \i[818] , \i[819] , \i[820] , \i[821] , \i[822] , \i[823] , \i[824] ,
    \i[825] , \i[826] , \i[827] , \i[828] , \i[829] , \i[830] , \i[831] ,
    \i[832] , \i[833] , \i[834] , \i[835] , \i[836] , \i[837] , \i[838] ,
    \i[839] , \i[840] , \i[841] , \i[842] , \i[843] , \i[844] , \i[845] ,
    \i[846] , \i[847] , \i[848] , \i[849] , \i[850] , \i[851] , \i[852] ,
    \i[853] , \i[854] , \i[855] , \i[856] , \i[857] , \i[858] , \i[859] ,
    \i[860] , \i[861] , \i[862] , \i[863] , \i[864] , \i[865] , \i[866] ,
    \i[867] , \i[868] , \i[869] , \i[870] , \i[871] , \i[872] , \i[873] ,
    \i[874] , \i[875] , \i[876] , \i[877] , \i[878] , \i[879] , \i[880] ,
    \i[881] , \i[882] , \i[883] , \i[884] , \i[885] , \i[886] , \i[887] ,
    \i[888] , \i[889] , \i[890] , \i[891] , \i[892] , \i[893] , \i[894] ,
    \i[895] , \i[896] , \i[897] , \i[898] , \i[899] , \i[900] , \i[901] ,
    \i[902] , \i[903] , \i[904] , \i[905] , \i[906] , \i[907] , \i[908] ,
    \i[909] , \i[910] , \i[911] , \i[912] , \i[913] , \i[914] , \i[915] ,
    \i[916] , \i[917] , \i[918] , \i[919] , \i[920] , \i[921] , \i[922] ,
    \i[923] , \i[924] , \i[925] , \i[926] , \i[927] , \i[928] , \i[929] ,
    \i[930] , \i[931] , \i[932] , \i[933] , \i[934] , \i[935] , \i[936] ,
    \i[937] , \i[938] , \i[939] , \i[940] , \i[941] , \i[942] , \i[943] ,
    \i[944] , \i[945] , \i[946] , \i[947] , \i[948] , \i[949] , \i[950] ,
    \i[951] , \i[952] , \i[953] , \i[954] , \i[955] , \i[956] , \i[957] ,
    \i[958] , \i[959] , \i[960] , \i[961] , \i[962] , \i[963] , \i[964] ,
    \i[965] , \i[966] , \i[967] , \i[968] , \i[969] , \i[970] , \i[971] ,
    \i[972] , \i[973] , \i[974] , \i[975] , \i[976] , \i[977] , \i[978] ,
    \i[979] , \i[980] , \i[981] , \i[982] , \i[983] , \i[984] , \i[985] ,
    \i[986] , \i[987] , \i[988] , \i[989] , \i[990] , \i[991] , \i[992] ,
    \i[993] , \i[994] , \i[995] , \i[996] , \i[997] , \i[998] , \i[999] ,
    \i[1000] , \i[1001] , \i[1002] , \i[1003] , \i[1004] , \i[1005] ,
    \i[1006] , \i[1007] , \i[1008] , \i[1009] , \i[1010] , \i[1011] ,
    \i[1012] , \i[1013] , \i[1014] , \i[1015] , \i[1016] , \i[1017] ,
    \i[1018] , \i[1019] , \i[1020] , \i[1021] , \i[1022] , \i[1023] ,
    \i[1024] , \i[1025] , \i[1026] , \i[1027] , \i[1028] , \i[1029] ,
    \i[1030] , \i[1031] , \i[1032] , \i[1033] , \i[1034] , \i[1035] ,
    \i[1036] , \i[1037] , \i[1038] , \i[1039] , \i[1040] , \i[1041] ,
    \i[1042] , \i[1043] , \i[1044] , \i[1045] , \i[1046] , \i[1047] ,
    \i[1048] , \i[1049] , \i[1050] , \i[1051] , \i[1052] , \i[1053] ,
    \i[1054] , \i[1055] , \i[1056] , \i[1057] , \i[1058] , \i[1059] ,
    \i[1060] , \i[1061] , \i[1062] , \i[1063] , \i[1064] , \i[1065] ,
    \i[1066] , \i[1067] , \i[1068] , \i[1069] , \i[1070] , \i[1071] ,
    \i[1072] , \i[1073] , \i[1074] , \i[1075] , \i[1076] , \i[1077] ,
    \i[1078] , \i[1079] , \i[1080] , \i[1081] , \i[1082] , \i[1083] ,
    \i[1084] , \i[1085] , \i[1086] , \i[1087] , \i[1088] , \i[1089] ,
    \i[1090] , \i[1091] , \i[1092] , \i[1093] , \i[1094] , \i[1095] ,
    \i[1096] , \i[1097] , \i[1098] , \i[1099] , \i[1100] , \i[1101] ,
    \i[1102] , \i[1103] , \i[1104] , \i[1105] , \i[1106] , \i[1107] ,
    \i[1108] , \i[1109] , \i[1110] , \i[1111] , \i[1112] , \i[1113] ,
    \i[1114] , \i[1115] , \i[1116] , \i[1117] , \i[1118] , \i[1119] ,
    \i[1120] , \i[1121] , \i[1122] , \i[1123] , \i[1124] , \i[1125] ,
    \i[1126] , \i[1127] , \i[1128] , \i[1129] , \i[1130] , \i[1131] ,
    \i[1132] , \i[1133] , \i[1134] , \i[1135] , \i[1136] , \i[1137] ,
    \i[1138] , \i[1139] , \i[1140] , \i[1141] , \i[1142] , \i[1143] ,
    \i[1144] , \i[1145] , \i[1146] , \i[1147] , \i[1148] , \i[1149] ,
    \i[1150] , \i[1151] , \i[1152] , \i[1153] , \i[1154] , \i[1155] ,
    \i[1156] , \i[1157] , \i[1158] , \i[1159] , \i[1160] , \i[1161] ,
    \i[1162] , \i[1163] , \i[1164] , \i[1165] , \i[1166] , \i[1167] ,
    \i[1168] , \i[1169] , \i[1170] , \i[1171] , \i[1172] , \i[1173] ,
    \i[1174] , \i[1175] , \i[1176] , \i[1177] , \i[1178] , \i[1179] ,
    \i[1180] , \i[1181] , \i[1182] , \i[1183] , \i[1184] , \i[1185] ,
    \i[1186] , \i[1187] , \i[1188] , \i[1189] , \i[1190] , \i[1191] ,
    \i[1192] , \i[1193] , \i[1194] , \i[1195] , \i[1196] , \i[1197] ,
    \i[1198] , \i[1199] , \i[1200] , \i[1201] , \i[1202] , \i[1203] ,
    \i[1204] , \i[1205] , \i[1206] , \i[1207] , \i[1208] , \i[1209] ,
    \i[1210] , \i[1211] , \i[1212] , \i[1213] , \i[1214] , \i[1215] ,
    \i[1216] , \i[1217] , \i[1218] , \i[1219] , \i[1220] , \i[1221] ,
    \i[1222] , \i[1223] , \i[1224] , \i[1225] , \i[1226] , \i[1227] ,
    \i[1228] , \i[1229] , \i[1230] , \i[1231] , \i[1232] , \i[1233] ,
    \i[1234] , \i[1235] , \i[1236] , \i[1237] , \i[1238] , \i[1239] ,
    \i[1240] , \i[1241] , \i[1242] , \i[1243] , \i[1244] , \i[1245] ,
    \i[1246] , \i[1247] , \i[1248] , \i[1249] , \i[1250] , \i[1251] ,
    \i[1252] , \i[1253] , \i[1254] , \i[1255] , \i[1256] , \i[1257] ,
    \i[1258] , \i[1259] , \i[1260] , \i[1261] , \i[1262] , \i[1263] ,
    \i[1264] , \i[1265] , \i[1266] , \i[1267] , \i[1268] , \i[1269] ,
    \i[1270] , \i[1271] , \i[1272] , \i[1273] , \i[1274] , \i[1275] ,
    \i[1276] , \i[1277] , \i[1278] , \i[1279] , \i[1280] , \i[1281] ,
    \i[1282] , \i[1283] , \i[1284] , \i[1285] , \i[1286] , \i[1287] ,
    \i[1288] , \i[1289] , \i[1290] , \i[1291] , \i[1292] , \i[1293] ,
    \i[1294] , \i[1295] , \i[1296] , \i[1297] , \i[1298] , \i[1299] ,
    \i[1300] , \i[1301] , \i[1302] , \i[1303] , \i[1304] , \i[1305] ,
    \i[1306] , \i[1307] , \i[1308] , \i[1309] , \i[1310] , \i[1311] ,
    \i[1312] , \i[1313] , \i[1314] , \i[1315] , \i[1316] , \i[1317] ,
    \i[1318] , \i[1319] , \i[1320] , \i[1321] , \i[1322] , \i[1323] ,
    \i[1324] , \i[1325] , \i[1326] , \i[1327] , \i[1328] , \i[1329] ,
    \i[1330] , \i[1331] , \i[1332] , \i[1333] , \i[1334] , \i[1335] ,
    \i[1336] , \i[1337] , \i[1338] , \i[1339] , \i[1340] , \i[1341] ,
    \i[1342] , \i[1343] , \i[1344] , \i[1345] , \i[1346] , \i[1347] ,
    \i[1348] , \i[1349] , \i[1350] , \i[1351] , \i[1352] , \i[1353] ,
    \i[1354] , \i[1355] , \i[1356] , \i[1357] , \i[1358] , \i[1359] ,
    \i[1360] , \i[1361] , \i[1362] , \i[1363] , \i[1364] , \i[1365] ,
    \i[1366] , \i[1367] , \i[1368] , \i[1369] , \i[1370] , \i[1371] ,
    \i[1372] , \i[1373] , \i[1374] , \i[1375] , \i[1376] , \i[1377] ,
    \i[1378] , \i[1379] , \i[1380] , \i[1381] , \i[1382] , \i[1383] ,
    \i[1384] , \i[1385] , \i[1386] , \i[1387] , \i[1388] , \i[1389] ,
    \i[1390] , \i[1391] , \i[1392] , \i[1393] , \i[1394] , \i[1395] ,
    \i[1396] , \i[1397] , \i[1398] , \i[1399] , \i[1400] , \i[1401] ,
    \i[1402] , \i[1403] , \i[1404] , \i[1405] , \i[1406] , \i[1407] ,
    \i[1408] , \i[1409] , \i[1410] , \i[1411] , \i[1412] , \i[1413] ,
    \i[1414] , \i[1415] , \i[1416] , \i[1417] , \i[1418] , \i[1419] ,
    \i[1420] , \i[1421] , \i[1422] , \i[1423] , \i[1424] , \i[1425] ,
    \i[1426] , \i[1427] , \i[1428] , \i[1429] , \i[1430] , \i[1431] ,
    \i[1432] , \i[1433] , \i[1434] , \i[1435] , \i[1436] , \i[1437] ,
    \i[1438] , \i[1439] , \i[1440] , \i[1441] , \i[1442] , \i[1443] ,
    \i[1444] , \i[1445] , \i[1446] , \i[1447] , \i[1448] , \i[1449] ,
    \i[1450] , \i[1451] , \i[1452] , \i[1453] , \i[1454] , \i[1455] ,
    \i[1456] , \i[1457] , \i[1458] , \i[1459] , \i[1460] , \i[1461] ,
    \i[1462] , \i[1463] , \i[1464] , \i[1465] , \i[1466] , \i[1467] ,
    \i[1468] , \i[1469] , \i[1470] , \i[1471] , \i[1472] , \i[1473] ,
    \i[1474] , \i[1475] , \i[1476] , \i[1477] , \i[1478] , \i[1479] ,
    \i[1480] , \i[1481] , \i[1482] , \i[1483] , \i[1484] , \i[1485] ,
    \i[1486] , \i[1487] , \i[1488] , \i[1489] , \i[1490] , \i[1491] ,
    \i[1492] , \i[1493] , \i[1494] , \i[1495] , \i[1496] , \i[1497] ,
    \i[1498] , \i[1499] , \i[1500] , \i[1501] , \i[1502] , \i[1503] ,
    \i[1504] , \i[1505] , \i[1506] , \i[1507] , \i[1508] , \i[1509] ,
    \i[1510] , \i[1511] , \i[1512] , \i[1513] , \i[1514] , \i[1515] ,
    \i[1516] , \i[1517] , \i[1518] , \i[1519] , \i[1520] , \i[1521] ,
    \i[1522] , \i[1523] , \i[1524] , \i[1525] , \i[1526] , \i[1527] ,
    \i[1528] , \i[1529] , \i[1530] , \i[1531] , \i[1532] , \i[1533] ,
    \i[1534] , \i[1535] , \i[1536] , \i[1537] , \i[1538] , \i[1539] ,
    \i[1540] , \i[1541] , \i[1542] , \i[1543] , \i[1544] , \i[1545] ,
    \i[1546] , \i[1547] , \i[1548] , \i[1549] , \i[1550] , \i[1551] ,
    \i[1552] , \i[1553] , \i[1554] , \i[1555] , \i[1556] , \i[1557] ,
    \i[1558] , \i[1559] , \i[1560] , \i[1561] , \i[1562] , \i[1563] ,
    \i[1564] , \i[1565] , \i[1566] , \i[1567] , \i[1568] , \i[1569] ,
    \i[1570] , \i[1571] , \i[1572] , \i[1573] , \i[1574] , \i[1575] ,
    \i[1576] , \i[1577] , \i[1578] , \i[1579] , \i[1580] , \i[1581] ,
    \i[1582] , \i[1583] , \i[1584] , \i[1585] , \i[1586] , \i[1587] ,
    \i[1588] , \i[1589] , \i[1590] , \i[1591] , \i[1592] , \i[1593] ,
    \i[1594] , \i[1595] , \i[1596] , \i[1597] , \i[1598] , \i[1599] ,
    \i[1600] , \i[1601] , \i[1602] , \i[1603] , \i[1604] , \i[1605] ,
    \i[1606] , \i[1607] , \i[1608] , \i[1609] , \i[1610] , \i[1611] ,
    \i[1612] , \i[1613] , \i[1614] , \i[1615] , \i[1616] , \i[1617] ,
    \i[1618] , \i[1619] , \i[1620] , \i[1621] , \i[1622] , \i[1623] ,
    \i[1624] , \i[1625] , \i[1626] , \i[1627] , \i[1628] , \i[1629] ,
    \i[1630] , \i[1631] , \i[1632] , \i[1633] , \i[1634] , \i[1635] ,
    \i[1636] , \i[1637] , \i[1638] , \i[1639] , \i[1640] , \i[1641] ,
    \i[1642] , \i[1643] , \i[1644] , \i[1645] , \i[1646] , \i[1647] ,
    \i[1648] , \i[1649] , \i[1650] , \i[1651] , \i[1652] , \i[1653] ,
    \i[1654] , \i[1655] , \i[1656] , \i[1657] , \i[1658] , \i[1659] ,
    \i[1660] , \i[1661] , \i[1662] , \i[1663] , \i[1664] , \i[1665] ,
    \i[1666] , \i[1667] , \i[1668] , \i[1669] , \i[1670] , \i[1671] ,
    \i[1672] , \i[1673] , \i[1674] , \i[1675] , \i[1676] , \i[1677] ,
    \i[1678] , \i[1679] , \i[1680] , \i[1681] , \i[1682] , \i[1683] ,
    \i[1684] , \i[1685] , \i[1686] , \i[1687] , \i[1688] , \i[1689] ,
    \i[1690] , \i[1691] , \i[1692] , \i[1693] , \i[1694] , \i[1695] ,
    \i[1696] , \i[1697] , \i[1698] , \i[1699] , \i[1700] , \i[1701] ,
    \i[1702] , \i[1703] , \i[1704] , \i[1705] , \i[1706] , \i[1707] ,
    \i[1708] , \i[1709] , \i[1710] , \i[1711] , \i[1712] , \i[1713] ,
    \i[1714] , \i[1715] , \i[1716] , \i[1717] , \i[1718] , \i[1719] ,
    \i[1720] , \i[1721] , \i[1722] , \i[1723] , \i[1724] , \i[1725] ,
    \i[1726] , \i[1727] , \i[1728] , \i[1729] , \i[1730] , \i[1731] ,
    \i[1732] , \i[1733] , \i[1734] , \i[1735] , \i[1736] , \i[1737] ,
    \i[1738] , \i[1739] , \i[1740] , \i[1741] , \i[1742] , \i[1743] ,
    \i[1744] , \i[1745] , \i[1746] , \i[1747] , \i[1748] , \i[1749] ,
    \i[1750] , \i[1751] , \i[1752] , \i[1753] , \i[1754] , \i[1755] ,
    \i[1756] , \i[1757] , \i[1758] , \i[1759] , \i[1760] , \i[1761] ,
    \i[1762] , \i[1763] , \i[1764] , \i[1765] , \i[1766] , \i[1767] ,
    \i[1768] , \i[1769] , \i[1770] , \i[1771] , \i[1772] , \i[1773] ,
    \i[1774] , \i[1775] , \i[1776] , \i[1777] , \i[1778] , \i[1779] ,
    \i[1780] , \i[1781] , \i[1782] , \i[1783] , \i[1784] , \i[1785] ,
    \i[1786] , \i[1787] , \i[1788] , \i[1789] , \i[1790] , \i[1791] ,
    \i[1792] , \i[1793] , \i[1794] , \i[1795] , \i[1796] , \i[1797] ,
    \i[1798] , \i[1799] , \i[1800] , \i[1801] , \i[1802] , \i[1803] ,
    \i[1804] , \i[1805] , \i[1806] , \i[1807] , \i[1808] , \i[1809] ,
    \i[1810] , \i[1811] , \i[1812] , \i[1813] , \i[1814] , \i[1815] ,
    \i[1816] , \i[1817] , \i[1818] , \i[1819] , \i[1820] , \i[1821] ,
    \i[1822] , \i[1823] , \i[1824] , \i[1825] , \i[1826] , \i[1827] ,
    \i[1828] , \i[1829] , \i[1830] , \i[1831] , \i[1832] , \i[1833] ,
    \i[1834] , \i[1835] , \i[1836] , \i[1837] , \i[1838] , \i[1839] ,
    \i[1840] , \i[1841] , \i[1842] , \i[1843] , \i[1844] , \i[1845] ,
    \i[1846] , \i[1847] , \i[1848] , \i[1849] , \i[1850] , \i[1851] ,
    \i[1852] , \i[1853] , \i[1854] , \i[1855] , \i[1856] , \i[1857] ,
    \i[1858] , \i[1859] , \i[1860] , \i[1861] , \i[1862] , \i[1863] ,
    \i[1864] , \i[1865] , \i[1866] , \i[1867] , \i[1868] , \i[1869] ,
    \i[1870] , \i[1871] , \i[1872] , \i[1873] , \i[1874] , \i[1875] ,
    \i[1876] , \i[1877] , \i[1878] , \i[1879] , \i[1880] , \i[1881] ,
    \i[1882] , \i[1883] , \i[1884] , \i[1885] , \i[1886] , \i[1887] ,
    \i[1888] , \i[1889] , \i[1890] , \i[1891] , \i[1892] , \i[1893] ,
    \i[1894] , \i[1895] , \i[1896] , \i[1897] , \i[1898] , \i[1899] ,
    \i[1900] , \i[1901] , \i[1902] , \i[1903] , \i[1904] , \i[1905] ,
    \i[1906] , \i[1907] , \i[1908] , \i[1909] , \i[1910] , \i[1911] ,
    \i[1912] , \i[1913] , \i[1914] , \i[1915] , \i[1916] , \i[1917] ,
    \i[1918] , \i[1919] , \i[1920] , \i[1921] , \i[1922] , \i[1923] ,
    \i[1924] , \i[1925] , \i[1926] , \i[1927] , \i[1928] , \i[1929] ,
    \i[1930] , \i[1931] , \i[1932] , \i[1933] , \i[1934] , \i[1935] ,
    \i[1936] , \i[1937] , \i[1938] , \i[1939] , \i[1940] , \i[1941] ,
    \i[1942] , \i[1943] , \i[1944] , \i[1945] , \i[1946] , \i[1947] ,
    \i[1948] , \i[1949] , \i[1950] , \i[1951] , \i[1952] , \i[1953] ,
    \i[1954] , \i[1955] , \i[1956] , \i[1957] , \i[1958] , \i[1959] ,
    \i[1960] , \i[1961] , \i[1962] , \i[1963] , \i[1964] , \i[1965] ,
    \i[1966] , \i[1967] , \i[1968] , \i[1969] , \i[1970] , \i[1971] ,
    \i[1972] , \i[1973] , \i[1974] , \i[1975] , \i[1976] , \i[1977] ,
    \i[1978] , \i[1979] , \i[1980] , \i[1981] , \i[1982] , \i[1983] ,
    \i[1984] , \i[1985] , \i[1986] , \i[1987] , \i[1988] , \i[1989] ,
    \i[1990] , \i[1991] , \i[1992] , \i[1993] , \i[1994] , \i[1995] ,
    \i[1996] , \i[1997] , \i[1998] , \i[1999] , \i[2000] , \i[2001] ,
    \i[2002] , \i[2003] , \i[2004] , \i[2005] , \i[2006] , \i[2007] ,
    \i[2008] , \i[2009] , \i[2010] , \i[2011] , \i[2012] , \i[2013] ,
    \i[2014] , \i[2015] , \i[2016] , \i[2017] , \i[2018] , \i[2019] ,
    \i[2020] , \i[2021] , \i[2022] , \i[2023] , \i[2024] , \i[2025] ,
    \i[2026] , \i[2027] , \i[2028] , \i[2029] , \i[2030] , \i[2031] ,
    \i[2032] , \i[2033] , \i[2034] , \i[2035] , \i[2036] , \i[2037] ,
    \i[2038] , \i[2039] , \i[2040] , \i[2041] , \i[2042] , \i[2043] ,
    \i[2044] , \i[2045] , \i[2046] , \i[2047] , \i[2048] , \i[2049] ,
    \i[2050] , \i[2051] , \i[2052] , \i[2053] , \i[2054] , \i[2055] ,
    \i[2056] , \i[2057] , \i[2058] , \i[2059] , \i[2060] , \i[2061] ,
    \i[2062] , \i[2063] , \i[2064] , \i[2065] , \i[2066] , \i[2067] ,
    \i[2068] , \i[2069] , \i[2070] , \i[2071] , \i[2072] , \i[2073] ,
    \i[2074] , \i[2075] , \i[2076] , \i[2077] , \i[2078] , \i[2079] ,
    \i[2080] , \i[2081] , \i[2082] , \i[2083] , \i[2084] , \i[2085] ,
    \i[2086] , \i[2087] , \i[2088] , \i[2089] , \i[2090] , \i[2091] ,
    \i[2092] , \i[2093] , \i[2094] , \i[2095] , \i[2096] , \i[2097] ,
    \i[2098] , \i[2099] , \i[2100] , \i[2101] , \i[2102] , \i[2103] ,
    \i[2104] , \i[2105] , \i[2106] , \i[2107] , \i[2108] , \i[2109] ,
    \i[2110] , \i[2111] , \i[2112] , \i[2113] , \i[2114] , \i[2115] ,
    \i[2116] , \i[2117] , \i[2118] , \i[2119] , \i[2120] , \i[2121] ,
    \i[2122] , \i[2123] , \i[2124] , \i[2125] , \i[2126] , \i[2127] ,
    \i[2128] , \i[2129] , \i[2130] , \i[2131] , \i[2132] , \i[2133] ,
    \i[2134] , \i[2135] , \i[2136] , \i[2137] , \i[2138] , \i[2139] ,
    \i[2140] , \i[2141] , \i[2142] , \i[2143] , \i[2144] , \i[2145] ,
    \i[2146] , \i[2147] , \i[2148] , \i[2149] , \i[2150] , \i[2151] ,
    \i[2152] , \i[2153] , \i[2154] , \i[2155] , \i[2156] , \i[2157] ,
    \i[2158] , \i[2159] , \i[2160] , \i[2161] , \i[2162] , \i[2163] ,
    \i[2164] , \i[2165] , \i[2166] , \i[2167] , \i[2168] , \i[2169] ,
    \i[2170] , \i[2171] , \i[2172] , \i[2173] , \i[2174] , \i[2175] ,
    \i[2176] , \i[2177] , \i[2178] , \i[2179] , \i[2180] , \i[2181] ,
    \i[2182] , \i[2183] , \i[2184] , \i[2185] , \i[2186] , \i[2187] ,
    \i[2188] , \i[2189] , \i[2190] , \i[2191] , \i[2192] , \i[2193] ,
    \i[2194] , \i[2195] , \i[2196] , \i[2197] , \i[2198] , \i[2199] ,
    \i[2200] , \i[2201] , \i[2202] , \i[2203] , \i[2204] , \i[2205] ,
    \i[2206] , \i[2207] , \i[2208] , \i[2209] , \i[2210] , \i[2211] ,
    \i[2212] , \i[2213] , \i[2214] , \i[2215] , \i[2216] , \i[2217] ,
    \i[2218] , \i[2219] , \i[2220] , \i[2221] , \i[2222] , \i[2223] ,
    \i[2224] , \i[2225] , \i[2226] , \i[2227] , \i[2228] , \i[2229] ,
    \i[2230] , \i[2231] , \i[2232] , \i[2233] , \i[2234] , \i[2235] ,
    \i[2236] , \i[2237] , \i[2238] , \i[2239] , \i[2240] , \i[2241] ,
    \i[2242] , \i[2243] , \i[2244] , \i[2245] , \i[2246] , \i[2247] ,
    \i[2248] , \i[2249] , \i[2250] , \i[2251] , \i[2252] , \i[2253] ,
    \i[2254] , \i[2255] , \i[2256] , \i[2257] , \i[2258] , \i[2259] ,
    \i[2260] , \i[2261] , \i[2262] , \i[2263] , \i[2264] , \i[2265] ,
    \i[2266] , \i[2267] , \i[2268] , \i[2269] , \i[2270] , \i[2271] ,
    \i[2272] , \i[2273] , \i[2274] , \i[2275] , \i[2276] , \i[2277] ,
    \i[2278] , \i[2279] , \i[2280] , \i[2281] , \i[2282] , \i[2283] ,
    \i[2284] , \i[2285] , \i[2286] , \i[2287] , \i[2288] , \i[2289] ,
    \i[2290] , \i[2291] , \i[2292] , \i[2293] , \i[2294] , \i[2295] ,
    \i[2296] , \i[2297] , \i[2298] , \i[2299] , \i[2300] , \i[2301] ,
    \i[2302] , \i[2303] , \i[2304] , \i[2305] , \i[2306] , \i[2307] ,
    \i[2308] , \i[2309] , \i[2310] , \i[2311] , \i[2312] , \i[2313] ,
    \i[2314] , \i[2315] , \i[2316] , \i[2317] , \i[2318] , \i[2319] ,
    \i[2320] , \i[2321] , \i[2322] , \i[2323] , \i[2324] , \i[2325] ,
    \i[2326] , \i[2327] , \i[2328] , \i[2329] , \i[2330] , \i[2331] ,
    \i[2332] , \i[2333] , \i[2334] , \i[2335] , \i[2336] , \i[2337] ,
    \i[2338] , \i[2339] , \i[2340] , \i[2341] , \i[2342] , \i[2343] ,
    \i[2344] , \i[2345] , \i[2346] , \i[2347] , \i[2348] , \i[2349] ,
    \i[2350] , \i[2351] , \i[2352] , \i[2353] , \i[2354] , \i[2355] ,
    \i[2356] , \i[2357] , \i[2358] , \i[2359] , \i[2360] , \i[2361] ,
    \i[2362] , \i[2363] , \i[2364] , \i[2365] , \i[2366] , \i[2367] ,
    \i[2368] , \i[2369] , \i[2370] , \i[2371] , \i[2372] , \i[2373] ,
    \i[2374] , \i[2375] , \i[2376] , \i[2377] , \i[2378] , \i[2379] ,
    \i[2380] , \i[2381] , \i[2382] , \i[2383] , \i[2384] , \i[2385] ,
    \i[2386] , \i[2387] , \i[2388] , \i[2389] , \i[2390] , \i[2391] ,
    \i[2392] , \i[2393] , \i[2394] , \i[2395] , \i[2396] , \i[2397] ,
    \i[2398] , \i[2399] , \i[2400] , \i[2401] , \i[2402] , \i[2403] ,
    \i[2404] , \i[2405] , \i[2406] , \i[2407] , \i[2408] , \i[2409] ,
    \i[2410] , \i[2411] , \i[2412] , \i[2413] , \i[2414] , \i[2415] ,
    \i[2416] , \i[2417] , \i[2418] , \i[2419] , \i[2420] , \i[2421] ,
    \i[2422] , \i[2423] , \i[2424] , \i[2425] , \i[2426] , \i[2427] ,
    \i[2428] , \i[2429] , \i[2430] , \i[2431] , \i[2432] , \i[2433] ,
    \i[2434] , \i[2435] , \i[2436] , \i[2437] , \i[2438] , \i[2439] ,
    \i[2440] , \i[2441] , \i[2442] , \i[2443] , \i[2444] , \i[2445] ,
    \i[2446] , \i[2447] , \i[2448] , \i[2449] , \i[2450] , \i[2451] ,
    \i[2452] , \i[2453] , \i[2454] , \i[2455] , \i[2456] , \i[2457] ,
    \i[2458] , \i[2459] , \i[2460] , \i[2461] , \i[2462] , \i[2463] ,
    \i[2464] , \i[2465] , \i[2466] , \i[2467] , \i[2468] , \i[2469] ,
    \i[2470] , \i[2471] , \i[2472] , \i[2473] , \i[2474] , \i[2475] ,
    \i[2476] , \i[2477] , \i[2478] , \i[2479] , \i[2480] , \i[2481] ,
    \i[2482] , \i[2483] , \i[2484] , \i[2485] , \i[2486] , \i[2487] ,
    \i[2488] , \i[2489] , \i[2490] , \i[2491] , \i[2492] , \i[2493] ,
    \i[2494] , \i[2495] , \i[2496] , \i[2497] , \i[2498] , \i[2499] ,
    \i[2500] , \i[2501] , \i[2502] , \i[2503] , \i[2504] , \i[2505] ,
    \i[2506] , \i[2507] , \i[2508] , \i[2509] , \i[2510] , \i[2511] ,
    \i[2512] , \i[2513] , \i[2514] , \i[2515] , \i[2516] , \i[2517] ,
    \i[2518] , \i[2519] , \i[2520] , \i[2521] , \i[2522] , \i[2523] ,
    \i[2524] , \i[2525] , \i[2526] , \i[2527] , \i[2528] , \i[2529] ,
    \i[2530] , \i[2531] , \i[2532] , \i[2533] , \i[2534] , \i[2535] ,
    \i[2536] , \i[2537] , \i[2538] , \i[2539] , \i[2540] , \i[2541] ,
    \i[2542] , \i[2543] , \i[2544] , \i[2545] , \i[2546] , \i[2547] ,
    \i[2548] , \i[2549] , \i[2550] , \i[2551] , \i[2552] , \i[2553] ,
    \i[2554] , \i[2555] , \i[2556] , \i[2557] , \i[2558] , \i[2559] ,
    \i[2560] , \i[2561] , \i[2562] , \i[2563] , \i[2564] , \i[2565] ,
    \i[2566] , \i[2567] , \i[2568] , \i[2569] , \i[2570] , \i[2571] ,
    \i[2572] , \i[2573] , \i[2574] , \i[2575] , \i[2576] , \i[2577] ,
    \i[2578] , \i[2579] , \i[2580] , \i[2581] , \i[2582] , \i[2583] ,
    \i[2584] , \i[2585] , \i[2586] , \i[2587] , \i[2588] , \i[2589] ,
    \i[2590] , \i[2591] , \i[2592] , \i[2593] , \i[2594] , \i[2595] ,
    \i[2596] , \i[2597] , \i[2598] , \i[2599] , \i[2600] , \i[2601] ,
    \i[2602] , \i[2603] , \i[2604] , \i[2605] , \i[2606] , \i[2607] ,
    \i[2608] , \i[2609] , \i[2610] , \i[2611] , \i[2612] , \i[2613] ,
    \i[2614] , \i[2615] , \i[2616] , \i[2617] , \i[2618] , \i[2619] ,
    \i[2620] , \i[2621] , \i[2622] , \i[2623] , \i[2624] , \i[2625] ,
    \i[2626] , \i[2627] , \i[2628] , \i[2629] , \i[2630] , \i[2631] ,
    \i[2632] , \i[2633] , \i[2634] , \i[2635] , \i[2636] , \i[2637] ,
    \i[2638] , \i[2639] , \i[2640] , \i[2641] , \i[2642] , \i[2643] ,
    \i[2644] , \i[2645] , \i[2646] , \i[2647] , \i[2648] , \i[2649] ,
    \i[2650] , \i[2651] , \i[2652] , \i[2653] , \i[2654] , \i[2655] ,
    \i[2656] , \i[2657] , \i[2658] , \i[2659] , \i[2660] , \i[2661] ,
    \i[2662] , \i[2663] , \i[2664] , \i[2665] , \i[2666] , \i[2667] ,
    \i[2668] , \i[2669] , \i[2670] , \i[2671] , \i[2672] , \i[2673] ,
    \i[2674] , \i[2675] , \i[2676] , \i[2677] , \i[2678] , \i[2679] ,
    \i[2680] , \i[2681] , \i[2682] , \i[2683] , \i[2684] , \i[2685] ,
    \i[2686] , \i[2687] , \i[2688] , \i[2689] , \i[2690] , \i[2691] ,
    \i[2692] , \i[2693] , \i[2694] , \i[2695] , \i[2696] , \i[2697] ,
    \i[2698] , \i[2699] , \i[2700] , \i[2701] , \i[2702] , \i[2703] ,
    \i[2704] , \i[2705] , \i[2706] , \i[2707] , \i[2708] , \i[2709] ,
    \i[2710] , \i[2711] , \i[2712] , \i[2713] , \i[2714] , \i[2715] ,
    \i[2716] , \i[2717] , \i[2718] , \i[2719] , \i[2720] , \i[2721] ,
    \i[2722] , \i[2723] , \i[2724] , \i[2725] , \i[2726] , \i[2727] ,
    \i[2728] , \i[2729] , \i[2730] , \i[2731] , \i[2732] , \i[2733] ,
    \i[2734] , \i[2735] , \i[2736] , \i[2737] , \i[2738] , \i[2739] ,
    \i[2740] , \i[2741] , \i[2742] , \i[2743] , \i[2744] , \i[2745] ,
    \i[2746] , \i[2747] , \i[2748] , \i[2749] , \i[2750] , \i[2751] ,
    \i[2752] , \i[2753] , \i[2754] , \i[2755] , \i[2756] , \i[2757] ,
    \i[2758] , \i[2759] , \i[2760] , \i[2761] , \i[2762] , \i[2763] ,
    \i[2764] , \i[2765] , \i[2766] , \i[2767] , \i[2768] , \i[2769] ,
    \i[2770] , \i[2771] , \i[2772] , \i[2773] , \i[2774] , \i[2775] ,
    \i[2776] , \i[2777] , \i[2778] , \i[2779] , \i[2780] , \i[2781] ,
    \i[2782] , \i[2783] , \i[2784] , \i[2785] , \i[2786] , \i[2787] ,
    \i[2788] , \i[2789] , \i[2790] , \i[2791] , \i[2792] , \i[2793] ,
    \i[2794] , \i[2795] , \i[2796] , \i[2797] , \i[2798] , \i[2799] ,
    \i[2800] , \i[2801] , \i[2802] , \i[2803] , \i[2804] , \i[2805] ,
    \i[2806] , \i[2807] , \i[2808] , \i[2809] , \i[2810] , \i[2811] ,
    \i[2812] , \i[2813] , \i[2814] , \i[2815] , \i[2816] , \i[2817] ,
    \i[2818] , \i[2819] , \i[2820] , \i[2821] , \i[2822] , \i[2823] ,
    \i[2824] , \i[2825] , \i[2826] , \i[2827] , \i[2828] , \i[2829] ,
    \i[2830] , \i[2831] , \i[2832] , \i[2833] , \i[2834] , \i[2835] ,
    \i[2836] , \i[2837] , \i[2838] , \i[2839] , \i[2840] , \i[2841] ,
    \i[2842] , \i[2843] , \i[2844] , \i[2845] , \i[2846] , \i[2847] ,
    \i[2848] , \i[2849] , \i[2850] , \i[2851] , \i[2852] , \i[2853] ,
    \i[2854] , \i[2855] , \i[2856] , \i[2857] , \i[2858] , \i[2859] ,
    \i[2860] , \i[2861] , \i[2862] , \i[2863] , \i[2864] , \i[2865] ,
    \i[2866] , \i[2867] , \i[2868] , \i[2869] , \i[2870] , \i[2871] ,
    \i[2872] , \i[2873] , \i[2874] , \i[2875] , \i[2876] , \i[2877] ,
    \i[2878] , \i[2879] , \i[2880] , \i[2881] , \i[2882] , \i[2883] ,
    \i[2884] , \i[2885] , \i[2886] , \i[2887] , \i[2888] , \i[2889] ,
    \i[2890] , \i[2891] , \i[2892] , \i[2893] , \i[2894] , \i[2895] ,
    \i[2896] , \i[2897] , \i[2898] , \i[2899] , \i[2900] , \i[2901] ,
    \i[2902] , \i[2903] , \i[2904] , \i[2905] , \i[2906] , \i[2907] ,
    \i[2908] , \i[2909] , \i[2910] , \i[2911] , \i[2912] , \i[2913] ,
    \i[2914] , \i[2915] , \i[2916] , \i[2917] , \i[2918] , \i[2919] ,
    \i[2920] , \i[2921] , \i[2922] , \i[2923] , \i[2924] , \i[2925] ,
    \i[2926] , \i[2927] , \i[2928] , \i[2929] , \i[2930] , \i[2931] ,
    \i[2932] , \i[2933] , \i[2934] , \i[2935] , \i[2936] , \i[2937] ,
    \i[2938] , \i[2939] , \i[2940] , \i[2941] , \i[2942] , \i[2943] ,
    \i[2944] , \i[2945] , \i[2946] , \i[2947] , \i[2948] , \i[2949] ,
    \i[2950] , \i[2951] , \i[2952] , \i[2953] , \i[2954] , \i[2955] ,
    \i[2956] , \i[2957] , \i[2958] , \i[2959] , \i[2960] , \i[2961] ,
    \i[2962] , \i[2963] , \i[2964] , \i[2965] , \i[2966] , \i[2967] ,
    \i[2968] , \i[2969] , \i[2970] , \i[2971] , \i[2972] , \i[2973] ,
    \i[2974] , \i[2975] , \i[2976] , \i[2977] , \i[2978] , \i[2979] ,
    \i[2980] , \i[2981] , \i[2982] , \i[2983] , \i[2984] , \i[2985] ,
    \i[2986] , \i[2987] , \i[2988] , \i[2989] , \i[2990] , \i[2991] ,
    \i[2992] , \i[2993] , \i[2994] , \i[2995] , \i[2996] , \i[2997] ,
    \i[2998] , \i[2999] , \i[3000] , \i[3001] , \i[3002] , \i[3003] ,
    \i[3004] , \i[3005] , \i[3006] , \i[3007] , \i[3008] , \i[3009] ,
    \i[3010] , \i[3011] , \i[3012] , \i[3013] , \i[3014] , \i[3015] ,
    \i[3016] , \i[3017] , \i[3018] , \i[3019] , \i[3020] , \i[3021] ,
    \i[3022] , \i[3023] , \i[3024] , \i[3025] , \i[3026] , \i[3027] ,
    \i[3028] , \i[3029] , \i[3030] , \i[3031] , \i[3032] , \i[3033] ,
    \i[3034] , \i[3035] , \i[3036] , \i[3037] , \i[3038] , \i[3039] ,
    \i[3040] , \i[3041] , \i[3042] , \i[3043] , \i[3044] , \i[3045] ,
    \i[3046] , \i[3047] , \i[3048] , \i[3049] , \i[3050] , \i[3051] ,
    \i[3052] , \i[3053] , \i[3054] , \i[3055] , \i[3056] , \i[3057] ,
    \i[3058] , \i[3059] , \i[3060] , \i[3061] , \i[3062] , \i[3063] ,
    \i[3064] , \i[3065] , \i[3066] , \i[3067] , \i[3068] , \i[3069] ,
    \i[3070] , \i[3071] , \i[3072] , \i[3073] , \i[3074] , \i[3075] ,
    \i[3076] , \i[3077] , \i[3078] , \i[3079] , \i[3080] , \i[3081] ,
    \i[3082] , \i[3083] , \i[3084] , \i[3085] , \i[3086] , \i[3087] ,
    \i[3088] , \i[3089] , \i[3090] , \i[3091] , \i[3092] , \i[3093] ,
    \i[3094] , \i[3095] , \i[3096] , \i[3097] , \i[3098] , \i[3099] ,
    \i[3100] , \i[3101] , \i[3102] , \i[3103] , \i[3104] , \i[3105] ,
    \i[3106] , \i[3107] , \i[3108] , \i[3109] , \i[3110] , \i[3111] ,
    \i[3112] , \i[3113] , \i[3114] , \i[3115] , \i[3116] , \i[3117] ,
    \i[3118] , \i[3119] , \i[3120] , \i[3121] , \i[3122] , \i[3123] ,
    \i[3124] , \i[3125] , \i[3126] , \i[3127] , \i[3128] , \i[3129] ,
    \i[3130] , \i[3131] , \i[3132] , \i[3133] , \i[3134] , \i[3135] ,
    \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] , \o[8] ,
    \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] , \o[16] ,
    \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] , \o[24] ,
    \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] , \o[32] ,
    \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] , \o[40] ,
    \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] , \o[48] ,
    \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] , \o[56] ,
    \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] , \o[64] ,
    \o[65] , \o[66] , \o[67] , \o[68] , \o[69]   );
  input  \i[0] , \i[1] , \i[2] , \i[3] , \i[4] , \i[5] , \i[6] , \i[7] ,
    \i[8] , \i[9] , \i[10] , \i[11] , \i[12] , \i[13] , \i[14] , \i[15] ,
    \i[16] , \i[17] , \i[18] , \i[19] , \i[20] , \i[21] , \i[22] , \i[23] ,
    \i[24] , \i[25] , \i[26] , \i[27] , \i[28] , \i[29] , \i[30] , \i[31] ,
    \i[32] , \i[33] , \i[34] , \i[35] , \i[36] , \i[37] , \i[38] , \i[39] ,
    \i[40] , \i[41] , \i[42] , \i[43] , \i[44] , \i[45] , \i[46] , \i[47] ,
    \i[48] , \i[49] , \i[50] , \i[51] , \i[52] , \i[53] , \i[54] , \i[55] ,
    \i[56] , \i[57] , \i[58] , \i[59] , \i[60] , \i[61] , \i[62] , \i[63] ,
    \i[64] , \i[65] , \i[66] , \i[67] , \i[68] , \i[69] , \i[70] , \i[71] ,
    \i[72] , \i[73] , \i[74] , \i[75] , \i[76] , \i[77] , \i[78] , \i[79] ,
    \i[80] , \i[81] , \i[82] , \i[83] , \i[84] , \i[85] , \i[86] , \i[87] ,
    \i[88] , \i[89] , \i[90] , \i[91] , \i[92] , \i[93] , \i[94] , \i[95] ,
    \i[96] , \i[97] , \i[98] , \i[99] , \i[100] , \i[101] , \i[102] ,
    \i[103] , \i[104] , \i[105] , \i[106] , \i[107] , \i[108] , \i[109] ,
    \i[110] , \i[111] , \i[112] , \i[113] , \i[114] , \i[115] , \i[116] ,
    \i[117] , \i[118] , \i[119] , \i[120] , \i[121] , \i[122] , \i[123] ,
    \i[124] , \i[125] , \i[126] , \i[127] , \i[128] , \i[129] , \i[130] ,
    \i[131] , \i[132] , \i[133] , \i[134] , \i[135] , \i[136] , \i[137] ,
    \i[138] , \i[139] , \i[140] , \i[141] , \i[142] , \i[143] , \i[144] ,
    \i[145] , \i[146] , \i[147] , \i[148] , \i[149] , \i[150] , \i[151] ,
    \i[152] , \i[153] , \i[154] , \i[155] , \i[156] , \i[157] , \i[158] ,
    \i[159] , \i[160] , \i[161] , \i[162] , \i[163] , \i[164] , \i[165] ,
    \i[166] , \i[167] , \i[168] , \i[169] , \i[170] , \i[171] , \i[172] ,
    \i[173] , \i[174] , \i[175] , \i[176] , \i[177] , \i[178] , \i[179] ,
    \i[180] , \i[181] , \i[182] , \i[183] , \i[184] , \i[185] , \i[186] ,
    \i[187] , \i[188] , \i[189] , \i[190] , \i[191] , \i[192] , \i[193] ,
    \i[194] , \i[195] , \i[196] , \i[197] , \i[198] , \i[199] , \i[200] ,
    \i[201] , \i[202] , \i[203] , \i[204] , \i[205] , \i[206] , \i[207] ,
    \i[208] , \i[209] , \i[210] , \i[211] , \i[212] , \i[213] , \i[214] ,
    \i[215] , \i[216] , \i[217] , \i[218] , \i[219] , \i[220] , \i[221] ,
    \i[222] , \i[223] , \i[224] , \i[225] , \i[226] , \i[227] , \i[228] ,
    \i[229] , \i[230] , \i[231] , \i[232] , \i[233] , \i[234] , \i[235] ,
    \i[236] , \i[237] , \i[238] , \i[239] , \i[240] , \i[241] , \i[242] ,
    \i[243] , \i[244] , \i[245] , \i[246] , \i[247] , \i[248] , \i[249] ,
    \i[250] , \i[251] , \i[252] , \i[253] , \i[254] , \i[255] , \i[256] ,
    \i[257] , \i[258] , \i[259] , \i[260] , \i[261] , \i[262] , \i[263] ,
    \i[264] , \i[265] , \i[266] , \i[267] , \i[268] , \i[269] , \i[270] ,
    \i[271] , \i[272] , \i[273] , \i[274] , \i[275] , \i[276] , \i[277] ,
    \i[278] , \i[279] , \i[280] , \i[281] , \i[282] , \i[283] , \i[284] ,
    \i[285] , \i[286] , \i[287] , \i[288] , \i[289] , \i[290] , \i[291] ,
    \i[292] , \i[293] , \i[294] , \i[295] , \i[296] , \i[297] , \i[298] ,
    \i[299] , \i[300] , \i[301] , \i[302] , \i[303] , \i[304] , \i[305] ,
    \i[306] , \i[307] , \i[308] , \i[309] , \i[310] , \i[311] , \i[312] ,
    \i[313] , \i[314] , \i[315] , \i[316] , \i[317] , \i[318] , \i[319] ,
    \i[320] , \i[321] , \i[322] , \i[323] , \i[324] , \i[325] , \i[326] ,
    \i[327] , \i[328] , \i[329] , \i[330] , \i[331] , \i[332] , \i[333] ,
    \i[334] , \i[335] , \i[336] , \i[337] , \i[338] , \i[339] , \i[340] ,
    \i[341] , \i[342] , \i[343] , \i[344] , \i[345] , \i[346] , \i[347] ,
    \i[348] , \i[349] , \i[350] , \i[351] , \i[352] , \i[353] , \i[354] ,
    \i[355] , \i[356] , \i[357] , \i[358] , \i[359] , \i[360] , \i[361] ,
    \i[362] , \i[363] , \i[364] , \i[365] , \i[366] , \i[367] , \i[368] ,
    \i[369] , \i[370] , \i[371] , \i[372] , \i[373] , \i[374] , \i[375] ,
    \i[376] , \i[377] , \i[378] , \i[379] , \i[380] , \i[381] , \i[382] ,
    \i[383] , \i[384] , \i[385] , \i[386] , \i[387] , \i[388] , \i[389] ,
    \i[390] , \i[391] , \i[392] , \i[393] , \i[394] , \i[395] , \i[396] ,
    \i[397] , \i[398] , \i[399] , \i[400] , \i[401] , \i[402] , \i[403] ,
    \i[404] , \i[405] , \i[406] , \i[407] , \i[408] , \i[409] , \i[410] ,
    \i[411] , \i[412] , \i[413] , \i[414] , \i[415] , \i[416] , \i[417] ,
    \i[418] , \i[419] , \i[420] , \i[421] , \i[422] , \i[423] , \i[424] ,
    \i[425] , \i[426] , \i[427] , \i[428] , \i[429] , \i[430] , \i[431] ,
    \i[432] , \i[433] , \i[434] , \i[435] , \i[436] , \i[437] , \i[438] ,
    \i[439] , \i[440] , \i[441] , \i[442] , \i[443] , \i[444] , \i[445] ,
    \i[446] , \i[447] , \i[448] , \i[449] , \i[450] , \i[451] , \i[452] ,
    \i[453] , \i[454] , \i[455] , \i[456] , \i[457] , \i[458] , \i[459] ,
    \i[460] , \i[461] , \i[462] , \i[463] , \i[464] , \i[465] , \i[466] ,
    \i[467] , \i[468] , \i[469] , \i[470] , \i[471] , \i[472] , \i[473] ,
    \i[474] , \i[475] , \i[476] , \i[477] , \i[478] , \i[479] , \i[480] ,
    \i[481] , \i[482] , \i[483] , \i[484] , \i[485] , \i[486] , \i[487] ,
    \i[488] , \i[489] , \i[490] , \i[491] , \i[492] , \i[493] , \i[494] ,
    \i[495] , \i[496] , \i[497] , \i[498] , \i[499] , \i[500] , \i[501] ,
    \i[502] , \i[503] , \i[504] , \i[505] , \i[506] , \i[507] , \i[508] ,
    \i[509] , \i[510] , \i[511] , \i[512] , \i[513] , \i[514] , \i[515] ,
    \i[516] , \i[517] , \i[518] , \i[519] , \i[520] , \i[521] , \i[522] ,
    \i[523] , \i[524] , \i[525] , \i[526] , \i[527] , \i[528] , \i[529] ,
    \i[530] , \i[531] , \i[532] , \i[533] , \i[534] , \i[535] , \i[536] ,
    \i[537] , \i[538] , \i[539] , \i[540] , \i[541] , \i[542] , \i[543] ,
    \i[544] , \i[545] , \i[546] , \i[547] , \i[548] , \i[549] , \i[550] ,
    \i[551] , \i[552] , \i[553] , \i[554] , \i[555] , \i[556] , \i[557] ,
    \i[558] , \i[559] , \i[560] , \i[561] , \i[562] , \i[563] , \i[564] ,
    \i[565] , \i[566] , \i[567] , \i[568] , \i[569] , \i[570] , \i[571] ,
    \i[572] , \i[573] , \i[574] , \i[575] , \i[576] , \i[577] , \i[578] ,
    \i[579] , \i[580] , \i[581] , \i[582] , \i[583] , \i[584] , \i[585] ,
    \i[586] , \i[587] , \i[588] , \i[589] , \i[590] , \i[591] , \i[592] ,
    \i[593] , \i[594] , \i[595] , \i[596] , \i[597] , \i[598] , \i[599] ,
    \i[600] , \i[601] , \i[602] , \i[603] , \i[604] , \i[605] , \i[606] ,
    \i[607] , \i[608] , \i[609] , \i[610] , \i[611] , \i[612] , \i[613] ,
    \i[614] , \i[615] , \i[616] , \i[617] , \i[618] , \i[619] , \i[620] ,
    \i[621] , \i[622] , \i[623] , \i[624] , \i[625] , \i[626] , \i[627] ,
    \i[628] , \i[629] , \i[630] , \i[631] , \i[632] , \i[633] , \i[634] ,
    \i[635] , \i[636] , \i[637] , \i[638] , \i[639] , \i[640] , \i[641] ,
    \i[642] , \i[643] , \i[644] , \i[645] , \i[646] , \i[647] , \i[648] ,
    \i[649] , \i[650] , \i[651] , \i[652] , \i[653] , \i[654] , \i[655] ,
    \i[656] , \i[657] , \i[658] , \i[659] , \i[660] , \i[661] , \i[662] ,
    \i[663] , \i[664] , \i[665] , \i[666] , \i[667] , \i[668] , \i[669] ,
    \i[670] , \i[671] , \i[672] , \i[673] , \i[674] , \i[675] , \i[676] ,
    \i[677] , \i[678] , \i[679] , \i[680] , \i[681] , \i[682] , \i[683] ,
    \i[684] , \i[685] , \i[686] , \i[687] , \i[688] , \i[689] , \i[690] ,
    \i[691] , \i[692] , \i[693] , \i[694] , \i[695] , \i[696] , \i[697] ,
    \i[698] , \i[699] , \i[700] , \i[701] , \i[702] , \i[703] , \i[704] ,
    \i[705] , \i[706] , \i[707] , \i[708] , \i[709] , \i[710] , \i[711] ,
    \i[712] , \i[713] , \i[714] , \i[715] , \i[716] , \i[717] , \i[718] ,
    \i[719] , \i[720] , \i[721] , \i[722] , \i[723] , \i[724] , \i[725] ,
    \i[726] , \i[727] , \i[728] , \i[729] , \i[730] , \i[731] , \i[732] ,
    \i[733] , \i[734] , \i[735] , \i[736] , \i[737] , \i[738] , \i[739] ,
    \i[740] , \i[741] , \i[742] , \i[743] , \i[744] , \i[745] , \i[746] ,
    \i[747] , \i[748] , \i[749] , \i[750] , \i[751] , \i[752] , \i[753] ,
    \i[754] , \i[755] , \i[756] , \i[757] , \i[758] , \i[759] , \i[760] ,
    \i[761] , \i[762] , \i[763] , \i[764] , \i[765] , \i[766] , \i[767] ,
    \i[768] , \i[769] , \i[770] , \i[771] , \i[772] , \i[773] , \i[774] ,
    \i[775] , \i[776] , \i[777] , \i[778] , \i[779] , \i[780] , \i[781] ,
    \i[782] , \i[783] , \i[784] , \i[785] , \i[786] , \i[787] , \i[788] ,
    \i[789] , \i[790] , \i[791] , \i[792] , \i[793] , \i[794] , \i[795] ,
    \i[796] , \i[797] , \i[798] , \i[799] , \i[800] , \i[801] , \i[802] ,
    \i[803] , \i[804] , \i[805] , \i[806] , \i[807] , \i[808] , \i[809] ,
    \i[810] , \i[811] , \i[812] , \i[813] , \i[814] , \i[815] , \i[816] ,
    \i[817] , \i[818] , \i[819] , \i[820] , \i[821] , \i[822] , \i[823] ,
    \i[824] , \i[825] , \i[826] , \i[827] , \i[828] , \i[829] , \i[830] ,
    \i[831] , \i[832] , \i[833] , \i[834] , \i[835] , \i[836] , \i[837] ,
    \i[838] , \i[839] , \i[840] , \i[841] , \i[842] , \i[843] , \i[844] ,
    \i[845] , \i[846] , \i[847] , \i[848] , \i[849] , \i[850] , \i[851] ,
    \i[852] , \i[853] , \i[854] , \i[855] , \i[856] , \i[857] , \i[858] ,
    \i[859] , \i[860] , \i[861] , \i[862] , \i[863] , \i[864] , \i[865] ,
    \i[866] , \i[867] , \i[868] , \i[869] , \i[870] , \i[871] , \i[872] ,
    \i[873] , \i[874] , \i[875] , \i[876] , \i[877] , \i[878] , \i[879] ,
    \i[880] , \i[881] , \i[882] , \i[883] , \i[884] , \i[885] , \i[886] ,
    \i[887] , \i[888] , \i[889] , \i[890] , \i[891] , \i[892] , \i[893] ,
    \i[894] , \i[895] , \i[896] , \i[897] , \i[898] , \i[899] , \i[900] ,
    \i[901] , \i[902] , \i[903] , \i[904] , \i[905] , \i[906] , \i[907] ,
    \i[908] , \i[909] , \i[910] , \i[911] , \i[912] , \i[913] , \i[914] ,
    \i[915] , \i[916] , \i[917] , \i[918] , \i[919] , \i[920] , \i[921] ,
    \i[922] , \i[923] , \i[924] , \i[925] , \i[926] , \i[927] , \i[928] ,
    \i[929] , \i[930] , \i[931] , \i[932] , \i[933] , \i[934] , \i[935] ,
    \i[936] , \i[937] , \i[938] , \i[939] , \i[940] , \i[941] , \i[942] ,
    \i[943] , \i[944] , \i[945] , \i[946] , \i[947] , \i[948] , \i[949] ,
    \i[950] , \i[951] , \i[952] , \i[953] , \i[954] , \i[955] , \i[956] ,
    \i[957] , \i[958] , \i[959] , \i[960] , \i[961] , \i[962] , \i[963] ,
    \i[964] , \i[965] , \i[966] , \i[967] , \i[968] , \i[969] , \i[970] ,
    \i[971] , \i[972] , \i[973] , \i[974] , \i[975] , \i[976] , \i[977] ,
    \i[978] , \i[979] , \i[980] , \i[981] , \i[982] , \i[983] , \i[984] ,
    \i[985] , \i[986] , \i[987] , \i[988] , \i[989] , \i[990] , \i[991] ,
    \i[992] , \i[993] , \i[994] , \i[995] , \i[996] , \i[997] , \i[998] ,
    \i[999] , \i[1000] , \i[1001] , \i[1002] , \i[1003] , \i[1004] ,
    \i[1005] , \i[1006] , \i[1007] , \i[1008] , \i[1009] , \i[1010] ,
    \i[1011] , \i[1012] , \i[1013] , \i[1014] , \i[1015] , \i[1016] ,
    \i[1017] , \i[1018] , \i[1019] , \i[1020] , \i[1021] , \i[1022] ,
    \i[1023] , \i[1024] , \i[1025] , \i[1026] , \i[1027] , \i[1028] ,
    \i[1029] , \i[1030] , \i[1031] , \i[1032] , \i[1033] , \i[1034] ,
    \i[1035] , \i[1036] , \i[1037] , \i[1038] , \i[1039] , \i[1040] ,
    \i[1041] , \i[1042] , \i[1043] , \i[1044] , \i[1045] , \i[1046] ,
    \i[1047] , \i[1048] , \i[1049] , \i[1050] , \i[1051] , \i[1052] ,
    \i[1053] , \i[1054] , \i[1055] , \i[1056] , \i[1057] , \i[1058] ,
    \i[1059] , \i[1060] , \i[1061] , \i[1062] , \i[1063] , \i[1064] ,
    \i[1065] , \i[1066] , \i[1067] , \i[1068] , \i[1069] , \i[1070] ,
    \i[1071] , \i[1072] , \i[1073] , \i[1074] , \i[1075] , \i[1076] ,
    \i[1077] , \i[1078] , \i[1079] , \i[1080] , \i[1081] , \i[1082] ,
    \i[1083] , \i[1084] , \i[1085] , \i[1086] , \i[1087] , \i[1088] ,
    \i[1089] , \i[1090] , \i[1091] , \i[1092] , \i[1093] , \i[1094] ,
    \i[1095] , \i[1096] , \i[1097] , \i[1098] , \i[1099] , \i[1100] ,
    \i[1101] , \i[1102] , \i[1103] , \i[1104] , \i[1105] , \i[1106] ,
    \i[1107] , \i[1108] , \i[1109] , \i[1110] , \i[1111] , \i[1112] ,
    \i[1113] , \i[1114] , \i[1115] , \i[1116] , \i[1117] , \i[1118] ,
    \i[1119] , \i[1120] , \i[1121] , \i[1122] , \i[1123] , \i[1124] ,
    \i[1125] , \i[1126] , \i[1127] , \i[1128] , \i[1129] , \i[1130] ,
    \i[1131] , \i[1132] , \i[1133] , \i[1134] , \i[1135] , \i[1136] ,
    \i[1137] , \i[1138] , \i[1139] , \i[1140] , \i[1141] , \i[1142] ,
    \i[1143] , \i[1144] , \i[1145] , \i[1146] , \i[1147] , \i[1148] ,
    \i[1149] , \i[1150] , \i[1151] , \i[1152] , \i[1153] , \i[1154] ,
    \i[1155] , \i[1156] , \i[1157] , \i[1158] , \i[1159] , \i[1160] ,
    \i[1161] , \i[1162] , \i[1163] , \i[1164] , \i[1165] , \i[1166] ,
    \i[1167] , \i[1168] , \i[1169] , \i[1170] , \i[1171] , \i[1172] ,
    \i[1173] , \i[1174] , \i[1175] , \i[1176] , \i[1177] , \i[1178] ,
    \i[1179] , \i[1180] , \i[1181] , \i[1182] , \i[1183] , \i[1184] ,
    \i[1185] , \i[1186] , \i[1187] , \i[1188] , \i[1189] , \i[1190] ,
    \i[1191] , \i[1192] , \i[1193] , \i[1194] , \i[1195] , \i[1196] ,
    \i[1197] , \i[1198] , \i[1199] , \i[1200] , \i[1201] , \i[1202] ,
    \i[1203] , \i[1204] , \i[1205] , \i[1206] , \i[1207] , \i[1208] ,
    \i[1209] , \i[1210] , \i[1211] , \i[1212] , \i[1213] , \i[1214] ,
    \i[1215] , \i[1216] , \i[1217] , \i[1218] , \i[1219] , \i[1220] ,
    \i[1221] , \i[1222] , \i[1223] , \i[1224] , \i[1225] , \i[1226] ,
    \i[1227] , \i[1228] , \i[1229] , \i[1230] , \i[1231] , \i[1232] ,
    \i[1233] , \i[1234] , \i[1235] , \i[1236] , \i[1237] , \i[1238] ,
    \i[1239] , \i[1240] , \i[1241] , \i[1242] , \i[1243] , \i[1244] ,
    \i[1245] , \i[1246] , \i[1247] , \i[1248] , \i[1249] , \i[1250] ,
    \i[1251] , \i[1252] , \i[1253] , \i[1254] , \i[1255] , \i[1256] ,
    \i[1257] , \i[1258] , \i[1259] , \i[1260] , \i[1261] , \i[1262] ,
    \i[1263] , \i[1264] , \i[1265] , \i[1266] , \i[1267] , \i[1268] ,
    \i[1269] , \i[1270] , \i[1271] , \i[1272] , \i[1273] , \i[1274] ,
    \i[1275] , \i[1276] , \i[1277] , \i[1278] , \i[1279] , \i[1280] ,
    \i[1281] , \i[1282] , \i[1283] , \i[1284] , \i[1285] , \i[1286] ,
    \i[1287] , \i[1288] , \i[1289] , \i[1290] , \i[1291] , \i[1292] ,
    \i[1293] , \i[1294] , \i[1295] , \i[1296] , \i[1297] , \i[1298] ,
    \i[1299] , \i[1300] , \i[1301] , \i[1302] , \i[1303] , \i[1304] ,
    \i[1305] , \i[1306] , \i[1307] , \i[1308] , \i[1309] , \i[1310] ,
    \i[1311] , \i[1312] , \i[1313] , \i[1314] , \i[1315] , \i[1316] ,
    \i[1317] , \i[1318] , \i[1319] , \i[1320] , \i[1321] , \i[1322] ,
    \i[1323] , \i[1324] , \i[1325] , \i[1326] , \i[1327] , \i[1328] ,
    \i[1329] , \i[1330] , \i[1331] , \i[1332] , \i[1333] , \i[1334] ,
    \i[1335] , \i[1336] , \i[1337] , \i[1338] , \i[1339] , \i[1340] ,
    \i[1341] , \i[1342] , \i[1343] , \i[1344] , \i[1345] , \i[1346] ,
    \i[1347] , \i[1348] , \i[1349] , \i[1350] , \i[1351] , \i[1352] ,
    \i[1353] , \i[1354] , \i[1355] , \i[1356] , \i[1357] , \i[1358] ,
    \i[1359] , \i[1360] , \i[1361] , \i[1362] , \i[1363] , \i[1364] ,
    \i[1365] , \i[1366] , \i[1367] , \i[1368] , \i[1369] , \i[1370] ,
    \i[1371] , \i[1372] , \i[1373] , \i[1374] , \i[1375] , \i[1376] ,
    \i[1377] , \i[1378] , \i[1379] , \i[1380] , \i[1381] , \i[1382] ,
    \i[1383] , \i[1384] , \i[1385] , \i[1386] , \i[1387] , \i[1388] ,
    \i[1389] , \i[1390] , \i[1391] , \i[1392] , \i[1393] , \i[1394] ,
    \i[1395] , \i[1396] , \i[1397] , \i[1398] , \i[1399] , \i[1400] ,
    \i[1401] , \i[1402] , \i[1403] , \i[1404] , \i[1405] , \i[1406] ,
    \i[1407] , \i[1408] , \i[1409] , \i[1410] , \i[1411] , \i[1412] ,
    \i[1413] , \i[1414] , \i[1415] , \i[1416] , \i[1417] , \i[1418] ,
    \i[1419] , \i[1420] , \i[1421] , \i[1422] , \i[1423] , \i[1424] ,
    \i[1425] , \i[1426] , \i[1427] , \i[1428] , \i[1429] , \i[1430] ,
    \i[1431] , \i[1432] , \i[1433] , \i[1434] , \i[1435] , \i[1436] ,
    \i[1437] , \i[1438] , \i[1439] , \i[1440] , \i[1441] , \i[1442] ,
    \i[1443] , \i[1444] , \i[1445] , \i[1446] , \i[1447] , \i[1448] ,
    \i[1449] , \i[1450] , \i[1451] , \i[1452] , \i[1453] , \i[1454] ,
    \i[1455] , \i[1456] , \i[1457] , \i[1458] , \i[1459] , \i[1460] ,
    \i[1461] , \i[1462] , \i[1463] , \i[1464] , \i[1465] , \i[1466] ,
    \i[1467] , \i[1468] , \i[1469] , \i[1470] , \i[1471] , \i[1472] ,
    \i[1473] , \i[1474] , \i[1475] , \i[1476] , \i[1477] , \i[1478] ,
    \i[1479] , \i[1480] , \i[1481] , \i[1482] , \i[1483] , \i[1484] ,
    \i[1485] , \i[1486] , \i[1487] , \i[1488] , \i[1489] , \i[1490] ,
    \i[1491] , \i[1492] , \i[1493] , \i[1494] , \i[1495] , \i[1496] ,
    \i[1497] , \i[1498] , \i[1499] , \i[1500] , \i[1501] , \i[1502] ,
    \i[1503] , \i[1504] , \i[1505] , \i[1506] , \i[1507] , \i[1508] ,
    \i[1509] , \i[1510] , \i[1511] , \i[1512] , \i[1513] , \i[1514] ,
    \i[1515] , \i[1516] , \i[1517] , \i[1518] , \i[1519] , \i[1520] ,
    \i[1521] , \i[1522] , \i[1523] , \i[1524] , \i[1525] , \i[1526] ,
    \i[1527] , \i[1528] , \i[1529] , \i[1530] , \i[1531] , \i[1532] ,
    \i[1533] , \i[1534] , \i[1535] , \i[1536] , \i[1537] , \i[1538] ,
    \i[1539] , \i[1540] , \i[1541] , \i[1542] , \i[1543] , \i[1544] ,
    \i[1545] , \i[1546] , \i[1547] , \i[1548] , \i[1549] , \i[1550] ,
    \i[1551] , \i[1552] , \i[1553] , \i[1554] , \i[1555] , \i[1556] ,
    \i[1557] , \i[1558] , \i[1559] , \i[1560] , \i[1561] , \i[1562] ,
    \i[1563] , \i[1564] , \i[1565] , \i[1566] , \i[1567] , \i[1568] ,
    \i[1569] , \i[1570] , \i[1571] , \i[1572] , \i[1573] , \i[1574] ,
    \i[1575] , \i[1576] , \i[1577] , \i[1578] , \i[1579] , \i[1580] ,
    \i[1581] , \i[1582] , \i[1583] , \i[1584] , \i[1585] , \i[1586] ,
    \i[1587] , \i[1588] , \i[1589] , \i[1590] , \i[1591] , \i[1592] ,
    \i[1593] , \i[1594] , \i[1595] , \i[1596] , \i[1597] , \i[1598] ,
    \i[1599] , \i[1600] , \i[1601] , \i[1602] , \i[1603] , \i[1604] ,
    \i[1605] , \i[1606] , \i[1607] , \i[1608] , \i[1609] , \i[1610] ,
    \i[1611] , \i[1612] , \i[1613] , \i[1614] , \i[1615] , \i[1616] ,
    \i[1617] , \i[1618] , \i[1619] , \i[1620] , \i[1621] , \i[1622] ,
    \i[1623] , \i[1624] , \i[1625] , \i[1626] , \i[1627] , \i[1628] ,
    \i[1629] , \i[1630] , \i[1631] , \i[1632] , \i[1633] , \i[1634] ,
    \i[1635] , \i[1636] , \i[1637] , \i[1638] , \i[1639] , \i[1640] ,
    \i[1641] , \i[1642] , \i[1643] , \i[1644] , \i[1645] , \i[1646] ,
    \i[1647] , \i[1648] , \i[1649] , \i[1650] , \i[1651] , \i[1652] ,
    \i[1653] , \i[1654] , \i[1655] , \i[1656] , \i[1657] , \i[1658] ,
    \i[1659] , \i[1660] , \i[1661] , \i[1662] , \i[1663] , \i[1664] ,
    \i[1665] , \i[1666] , \i[1667] , \i[1668] , \i[1669] , \i[1670] ,
    \i[1671] , \i[1672] , \i[1673] , \i[1674] , \i[1675] , \i[1676] ,
    \i[1677] , \i[1678] , \i[1679] , \i[1680] , \i[1681] , \i[1682] ,
    \i[1683] , \i[1684] , \i[1685] , \i[1686] , \i[1687] , \i[1688] ,
    \i[1689] , \i[1690] , \i[1691] , \i[1692] , \i[1693] , \i[1694] ,
    \i[1695] , \i[1696] , \i[1697] , \i[1698] , \i[1699] , \i[1700] ,
    \i[1701] , \i[1702] , \i[1703] , \i[1704] , \i[1705] , \i[1706] ,
    \i[1707] , \i[1708] , \i[1709] , \i[1710] , \i[1711] , \i[1712] ,
    \i[1713] , \i[1714] , \i[1715] , \i[1716] , \i[1717] , \i[1718] ,
    \i[1719] , \i[1720] , \i[1721] , \i[1722] , \i[1723] , \i[1724] ,
    \i[1725] , \i[1726] , \i[1727] , \i[1728] , \i[1729] , \i[1730] ,
    \i[1731] , \i[1732] , \i[1733] , \i[1734] , \i[1735] , \i[1736] ,
    \i[1737] , \i[1738] , \i[1739] , \i[1740] , \i[1741] , \i[1742] ,
    \i[1743] , \i[1744] , \i[1745] , \i[1746] , \i[1747] , \i[1748] ,
    \i[1749] , \i[1750] , \i[1751] , \i[1752] , \i[1753] , \i[1754] ,
    \i[1755] , \i[1756] , \i[1757] , \i[1758] , \i[1759] , \i[1760] ,
    \i[1761] , \i[1762] , \i[1763] , \i[1764] , \i[1765] , \i[1766] ,
    \i[1767] , \i[1768] , \i[1769] , \i[1770] , \i[1771] , \i[1772] ,
    \i[1773] , \i[1774] , \i[1775] , \i[1776] , \i[1777] , \i[1778] ,
    \i[1779] , \i[1780] , \i[1781] , \i[1782] , \i[1783] , \i[1784] ,
    \i[1785] , \i[1786] , \i[1787] , \i[1788] , \i[1789] , \i[1790] ,
    \i[1791] , \i[1792] , \i[1793] , \i[1794] , \i[1795] , \i[1796] ,
    \i[1797] , \i[1798] , \i[1799] , \i[1800] , \i[1801] , \i[1802] ,
    \i[1803] , \i[1804] , \i[1805] , \i[1806] , \i[1807] , \i[1808] ,
    \i[1809] , \i[1810] , \i[1811] , \i[1812] , \i[1813] , \i[1814] ,
    \i[1815] , \i[1816] , \i[1817] , \i[1818] , \i[1819] , \i[1820] ,
    \i[1821] , \i[1822] , \i[1823] , \i[1824] , \i[1825] , \i[1826] ,
    \i[1827] , \i[1828] , \i[1829] , \i[1830] , \i[1831] , \i[1832] ,
    \i[1833] , \i[1834] , \i[1835] , \i[1836] , \i[1837] , \i[1838] ,
    \i[1839] , \i[1840] , \i[1841] , \i[1842] , \i[1843] , \i[1844] ,
    \i[1845] , \i[1846] , \i[1847] , \i[1848] , \i[1849] , \i[1850] ,
    \i[1851] , \i[1852] , \i[1853] , \i[1854] , \i[1855] , \i[1856] ,
    \i[1857] , \i[1858] , \i[1859] , \i[1860] , \i[1861] , \i[1862] ,
    \i[1863] , \i[1864] , \i[1865] , \i[1866] , \i[1867] , \i[1868] ,
    \i[1869] , \i[1870] , \i[1871] , \i[1872] , \i[1873] , \i[1874] ,
    \i[1875] , \i[1876] , \i[1877] , \i[1878] , \i[1879] , \i[1880] ,
    \i[1881] , \i[1882] , \i[1883] , \i[1884] , \i[1885] , \i[1886] ,
    \i[1887] , \i[1888] , \i[1889] , \i[1890] , \i[1891] , \i[1892] ,
    \i[1893] , \i[1894] , \i[1895] , \i[1896] , \i[1897] , \i[1898] ,
    \i[1899] , \i[1900] , \i[1901] , \i[1902] , \i[1903] , \i[1904] ,
    \i[1905] , \i[1906] , \i[1907] , \i[1908] , \i[1909] , \i[1910] ,
    \i[1911] , \i[1912] , \i[1913] , \i[1914] , \i[1915] , \i[1916] ,
    \i[1917] , \i[1918] , \i[1919] , \i[1920] , \i[1921] , \i[1922] ,
    \i[1923] , \i[1924] , \i[1925] , \i[1926] , \i[1927] , \i[1928] ,
    \i[1929] , \i[1930] , \i[1931] , \i[1932] , \i[1933] , \i[1934] ,
    \i[1935] , \i[1936] , \i[1937] , \i[1938] , \i[1939] , \i[1940] ,
    \i[1941] , \i[1942] , \i[1943] , \i[1944] , \i[1945] , \i[1946] ,
    \i[1947] , \i[1948] , \i[1949] , \i[1950] , \i[1951] , \i[1952] ,
    \i[1953] , \i[1954] , \i[1955] , \i[1956] , \i[1957] , \i[1958] ,
    \i[1959] , \i[1960] , \i[1961] , \i[1962] , \i[1963] , \i[1964] ,
    \i[1965] , \i[1966] , \i[1967] , \i[1968] , \i[1969] , \i[1970] ,
    \i[1971] , \i[1972] , \i[1973] , \i[1974] , \i[1975] , \i[1976] ,
    \i[1977] , \i[1978] , \i[1979] , \i[1980] , \i[1981] , \i[1982] ,
    \i[1983] , \i[1984] , \i[1985] , \i[1986] , \i[1987] , \i[1988] ,
    \i[1989] , \i[1990] , \i[1991] , \i[1992] , \i[1993] , \i[1994] ,
    \i[1995] , \i[1996] , \i[1997] , \i[1998] , \i[1999] , \i[2000] ,
    \i[2001] , \i[2002] , \i[2003] , \i[2004] , \i[2005] , \i[2006] ,
    \i[2007] , \i[2008] , \i[2009] , \i[2010] , \i[2011] , \i[2012] ,
    \i[2013] , \i[2014] , \i[2015] , \i[2016] , \i[2017] , \i[2018] ,
    \i[2019] , \i[2020] , \i[2021] , \i[2022] , \i[2023] , \i[2024] ,
    \i[2025] , \i[2026] , \i[2027] , \i[2028] , \i[2029] , \i[2030] ,
    \i[2031] , \i[2032] , \i[2033] , \i[2034] , \i[2035] , \i[2036] ,
    \i[2037] , \i[2038] , \i[2039] , \i[2040] , \i[2041] , \i[2042] ,
    \i[2043] , \i[2044] , \i[2045] , \i[2046] , \i[2047] , \i[2048] ,
    \i[2049] , \i[2050] , \i[2051] , \i[2052] , \i[2053] , \i[2054] ,
    \i[2055] , \i[2056] , \i[2057] , \i[2058] , \i[2059] , \i[2060] ,
    \i[2061] , \i[2062] , \i[2063] , \i[2064] , \i[2065] , \i[2066] ,
    \i[2067] , \i[2068] , \i[2069] , \i[2070] , \i[2071] , \i[2072] ,
    \i[2073] , \i[2074] , \i[2075] , \i[2076] , \i[2077] , \i[2078] ,
    \i[2079] , \i[2080] , \i[2081] , \i[2082] , \i[2083] , \i[2084] ,
    \i[2085] , \i[2086] , \i[2087] , \i[2088] , \i[2089] , \i[2090] ,
    \i[2091] , \i[2092] , \i[2093] , \i[2094] , \i[2095] , \i[2096] ,
    \i[2097] , \i[2098] , \i[2099] , \i[2100] , \i[2101] , \i[2102] ,
    \i[2103] , \i[2104] , \i[2105] , \i[2106] , \i[2107] , \i[2108] ,
    \i[2109] , \i[2110] , \i[2111] , \i[2112] , \i[2113] , \i[2114] ,
    \i[2115] , \i[2116] , \i[2117] , \i[2118] , \i[2119] , \i[2120] ,
    \i[2121] , \i[2122] , \i[2123] , \i[2124] , \i[2125] , \i[2126] ,
    \i[2127] , \i[2128] , \i[2129] , \i[2130] , \i[2131] , \i[2132] ,
    \i[2133] , \i[2134] , \i[2135] , \i[2136] , \i[2137] , \i[2138] ,
    \i[2139] , \i[2140] , \i[2141] , \i[2142] , \i[2143] , \i[2144] ,
    \i[2145] , \i[2146] , \i[2147] , \i[2148] , \i[2149] , \i[2150] ,
    \i[2151] , \i[2152] , \i[2153] , \i[2154] , \i[2155] , \i[2156] ,
    \i[2157] , \i[2158] , \i[2159] , \i[2160] , \i[2161] , \i[2162] ,
    \i[2163] , \i[2164] , \i[2165] , \i[2166] , \i[2167] , \i[2168] ,
    \i[2169] , \i[2170] , \i[2171] , \i[2172] , \i[2173] , \i[2174] ,
    \i[2175] , \i[2176] , \i[2177] , \i[2178] , \i[2179] , \i[2180] ,
    \i[2181] , \i[2182] , \i[2183] , \i[2184] , \i[2185] , \i[2186] ,
    \i[2187] , \i[2188] , \i[2189] , \i[2190] , \i[2191] , \i[2192] ,
    \i[2193] , \i[2194] , \i[2195] , \i[2196] , \i[2197] , \i[2198] ,
    \i[2199] , \i[2200] , \i[2201] , \i[2202] , \i[2203] , \i[2204] ,
    \i[2205] , \i[2206] , \i[2207] , \i[2208] , \i[2209] , \i[2210] ,
    \i[2211] , \i[2212] , \i[2213] , \i[2214] , \i[2215] , \i[2216] ,
    \i[2217] , \i[2218] , \i[2219] , \i[2220] , \i[2221] , \i[2222] ,
    \i[2223] , \i[2224] , \i[2225] , \i[2226] , \i[2227] , \i[2228] ,
    \i[2229] , \i[2230] , \i[2231] , \i[2232] , \i[2233] , \i[2234] ,
    \i[2235] , \i[2236] , \i[2237] , \i[2238] , \i[2239] , \i[2240] ,
    \i[2241] , \i[2242] , \i[2243] , \i[2244] , \i[2245] , \i[2246] ,
    \i[2247] , \i[2248] , \i[2249] , \i[2250] , \i[2251] , \i[2252] ,
    \i[2253] , \i[2254] , \i[2255] , \i[2256] , \i[2257] , \i[2258] ,
    \i[2259] , \i[2260] , \i[2261] , \i[2262] , \i[2263] , \i[2264] ,
    \i[2265] , \i[2266] , \i[2267] , \i[2268] , \i[2269] , \i[2270] ,
    \i[2271] , \i[2272] , \i[2273] , \i[2274] , \i[2275] , \i[2276] ,
    \i[2277] , \i[2278] , \i[2279] , \i[2280] , \i[2281] , \i[2282] ,
    \i[2283] , \i[2284] , \i[2285] , \i[2286] , \i[2287] , \i[2288] ,
    \i[2289] , \i[2290] , \i[2291] , \i[2292] , \i[2293] , \i[2294] ,
    \i[2295] , \i[2296] , \i[2297] , \i[2298] , \i[2299] , \i[2300] ,
    \i[2301] , \i[2302] , \i[2303] , \i[2304] , \i[2305] , \i[2306] ,
    \i[2307] , \i[2308] , \i[2309] , \i[2310] , \i[2311] , \i[2312] ,
    \i[2313] , \i[2314] , \i[2315] , \i[2316] , \i[2317] , \i[2318] ,
    \i[2319] , \i[2320] , \i[2321] , \i[2322] , \i[2323] , \i[2324] ,
    \i[2325] , \i[2326] , \i[2327] , \i[2328] , \i[2329] , \i[2330] ,
    \i[2331] , \i[2332] , \i[2333] , \i[2334] , \i[2335] , \i[2336] ,
    \i[2337] , \i[2338] , \i[2339] , \i[2340] , \i[2341] , \i[2342] ,
    \i[2343] , \i[2344] , \i[2345] , \i[2346] , \i[2347] , \i[2348] ,
    \i[2349] , \i[2350] , \i[2351] , \i[2352] , \i[2353] , \i[2354] ,
    \i[2355] , \i[2356] , \i[2357] , \i[2358] , \i[2359] , \i[2360] ,
    \i[2361] , \i[2362] , \i[2363] , \i[2364] , \i[2365] , \i[2366] ,
    \i[2367] , \i[2368] , \i[2369] , \i[2370] , \i[2371] , \i[2372] ,
    \i[2373] , \i[2374] , \i[2375] , \i[2376] , \i[2377] , \i[2378] ,
    \i[2379] , \i[2380] , \i[2381] , \i[2382] , \i[2383] , \i[2384] ,
    \i[2385] , \i[2386] , \i[2387] , \i[2388] , \i[2389] , \i[2390] ,
    \i[2391] , \i[2392] , \i[2393] , \i[2394] , \i[2395] , \i[2396] ,
    \i[2397] , \i[2398] , \i[2399] , \i[2400] , \i[2401] , \i[2402] ,
    \i[2403] , \i[2404] , \i[2405] , \i[2406] , \i[2407] , \i[2408] ,
    \i[2409] , \i[2410] , \i[2411] , \i[2412] , \i[2413] , \i[2414] ,
    \i[2415] , \i[2416] , \i[2417] , \i[2418] , \i[2419] , \i[2420] ,
    \i[2421] , \i[2422] , \i[2423] , \i[2424] , \i[2425] , \i[2426] ,
    \i[2427] , \i[2428] , \i[2429] , \i[2430] , \i[2431] , \i[2432] ,
    \i[2433] , \i[2434] , \i[2435] , \i[2436] , \i[2437] , \i[2438] ,
    \i[2439] , \i[2440] , \i[2441] , \i[2442] , \i[2443] , \i[2444] ,
    \i[2445] , \i[2446] , \i[2447] , \i[2448] , \i[2449] , \i[2450] ,
    \i[2451] , \i[2452] , \i[2453] , \i[2454] , \i[2455] , \i[2456] ,
    \i[2457] , \i[2458] , \i[2459] , \i[2460] , \i[2461] , \i[2462] ,
    \i[2463] , \i[2464] , \i[2465] , \i[2466] , \i[2467] , \i[2468] ,
    \i[2469] , \i[2470] , \i[2471] , \i[2472] , \i[2473] , \i[2474] ,
    \i[2475] , \i[2476] , \i[2477] , \i[2478] , \i[2479] , \i[2480] ,
    \i[2481] , \i[2482] , \i[2483] , \i[2484] , \i[2485] , \i[2486] ,
    \i[2487] , \i[2488] , \i[2489] , \i[2490] , \i[2491] , \i[2492] ,
    \i[2493] , \i[2494] , \i[2495] , \i[2496] , \i[2497] , \i[2498] ,
    \i[2499] , \i[2500] , \i[2501] , \i[2502] , \i[2503] , \i[2504] ,
    \i[2505] , \i[2506] , \i[2507] , \i[2508] , \i[2509] , \i[2510] ,
    \i[2511] , \i[2512] , \i[2513] , \i[2514] , \i[2515] , \i[2516] ,
    \i[2517] , \i[2518] , \i[2519] , \i[2520] , \i[2521] , \i[2522] ,
    \i[2523] , \i[2524] , \i[2525] , \i[2526] , \i[2527] , \i[2528] ,
    \i[2529] , \i[2530] , \i[2531] , \i[2532] , \i[2533] , \i[2534] ,
    \i[2535] , \i[2536] , \i[2537] , \i[2538] , \i[2539] , \i[2540] ,
    \i[2541] , \i[2542] , \i[2543] , \i[2544] , \i[2545] , \i[2546] ,
    \i[2547] , \i[2548] , \i[2549] , \i[2550] , \i[2551] , \i[2552] ,
    \i[2553] , \i[2554] , \i[2555] , \i[2556] , \i[2557] , \i[2558] ,
    \i[2559] , \i[2560] , \i[2561] , \i[2562] , \i[2563] , \i[2564] ,
    \i[2565] , \i[2566] , \i[2567] , \i[2568] , \i[2569] , \i[2570] ,
    \i[2571] , \i[2572] , \i[2573] , \i[2574] , \i[2575] , \i[2576] ,
    \i[2577] , \i[2578] , \i[2579] , \i[2580] , \i[2581] , \i[2582] ,
    \i[2583] , \i[2584] , \i[2585] , \i[2586] , \i[2587] , \i[2588] ,
    \i[2589] , \i[2590] , \i[2591] , \i[2592] , \i[2593] , \i[2594] ,
    \i[2595] , \i[2596] , \i[2597] , \i[2598] , \i[2599] , \i[2600] ,
    \i[2601] , \i[2602] , \i[2603] , \i[2604] , \i[2605] , \i[2606] ,
    \i[2607] , \i[2608] , \i[2609] , \i[2610] , \i[2611] , \i[2612] ,
    \i[2613] , \i[2614] , \i[2615] , \i[2616] , \i[2617] , \i[2618] ,
    \i[2619] , \i[2620] , \i[2621] , \i[2622] , \i[2623] , \i[2624] ,
    \i[2625] , \i[2626] , \i[2627] , \i[2628] , \i[2629] , \i[2630] ,
    \i[2631] , \i[2632] , \i[2633] , \i[2634] , \i[2635] , \i[2636] ,
    \i[2637] , \i[2638] , \i[2639] , \i[2640] , \i[2641] , \i[2642] ,
    \i[2643] , \i[2644] , \i[2645] , \i[2646] , \i[2647] , \i[2648] ,
    \i[2649] , \i[2650] , \i[2651] , \i[2652] , \i[2653] , \i[2654] ,
    \i[2655] , \i[2656] , \i[2657] , \i[2658] , \i[2659] , \i[2660] ,
    \i[2661] , \i[2662] , \i[2663] , \i[2664] , \i[2665] , \i[2666] ,
    \i[2667] , \i[2668] , \i[2669] , \i[2670] , \i[2671] , \i[2672] ,
    \i[2673] , \i[2674] , \i[2675] , \i[2676] , \i[2677] , \i[2678] ,
    \i[2679] , \i[2680] , \i[2681] , \i[2682] , \i[2683] , \i[2684] ,
    \i[2685] , \i[2686] , \i[2687] , \i[2688] , \i[2689] , \i[2690] ,
    \i[2691] , \i[2692] , \i[2693] , \i[2694] , \i[2695] , \i[2696] ,
    \i[2697] , \i[2698] , \i[2699] , \i[2700] , \i[2701] , \i[2702] ,
    \i[2703] , \i[2704] , \i[2705] , \i[2706] , \i[2707] , \i[2708] ,
    \i[2709] , \i[2710] , \i[2711] , \i[2712] , \i[2713] , \i[2714] ,
    \i[2715] , \i[2716] , \i[2717] , \i[2718] , \i[2719] , \i[2720] ,
    \i[2721] , \i[2722] , \i[2723] , \i[2724] , \i[2725] , \i[2726] ,
    \i[2727] , \i[2728] , \i[2729] , \i[2730] , \i[2731] , \i[2732] ,
    \i[2733] , \i[2734] , \i[2735] , \i[2736] , \i[2737] , \i[2738] ,
    \i[2739] , \i[2740] , \i[2741] , \i[2742] , \i[2743] , \i[2744] ,
    \i[2745] , \i[2746] , \i[2747] , \i[2748] , \i[2749] , \i[2750] ,
    \i[2751] , \i[2752] , \i[2753] , \i[2754] , \i[2755] , \i[2756] ,
    \i[2757] , \i[2758] , \i[2759] , \i[2760] , \i[2761] , \i[2762] ,
    \i[2763] , \i[2764] , \i[2765] , \i[2766] , \i[2767] , \i[2768] ,
    \i[2769] , \i[2770] , \i[2771] , \i[2772] , \i[2773] , \i[2774] ,
    \i[2775] , \i[2776] , \i[2777] , \i[2778] , \i[2779] , \i[2780] ,
    \i[2781] , \i[2782] , \i[2783] , \i[2784] , \i[2785] , \i[2786] ,
    \i[2787] , \i[2788] , \i[2789] , \i[2790] , \i[2791] , \i[2792] ,
    \i[2793] , \i[2794] , \i[2795] , \i[2796] , \i[2797] , \i[2798] ,
    \i[2799] , \i[2800] , \i[2801] , \i[2802] , \i[2803] , \i[2804] ,
    \i[2805] , \i[2806] , \i[2807] , \i[2808] , \i[2809] , \i[2810] ,
    \i[2811] , \i[2812] , \i[2813] , \i[2814] , \i[2815] , \i[2816] ,
    \i[2817] , \i[2818] , \i[2819] , \i[2820] , \i[2821] , \i[2822] ,
    \i[2823] , \i[2824] , \i[2825] , \i[2826] , \i[2827] , \i[2828] ,
    \i[2829] , \i[2830] , \i[2831] , \i[2832] , \i[2833] , \i[2834] ,
    \i[2835] , \i[2836] , \i[2837] , \i[2838] , \i[2839] , \i[2840] ,
    \i[2841] , \i[2842] , \i[2843] , \i[2844] , \i[2845] , \i[2846] ,
    \i[2847] , \i[2848] , \i[2849] , \i[2850] , \i[2851] , \i[2852] ,
    \i[2853] , \i[2854] , \i[2855] , \i[2856] , \i[2857] , \i[2858] ,
    \i[2859] , \i[2860] , \i[2861] , \i[2862] , \i[2863] , \i[2864] ,
    \i[2865] , \i[2866] , \i[2867] , \i[2868] , \i[2869] , \i[2870] ,
    \i[2871] , \i[2872] , \i[2873] , \i[2874] , \i[2875] , \i[2876] ,
    \i[2877] , \i[2878] , \i[2879] , \i[2880] , \i[2881] , \i[2882] ,
    \i[2883] , \i[2884] , \i[2885] , \i[2886] , \i[2887] , \i[2888] ,
    \i[2889] , \i[2890] , \i[2891] , \i[2892] , \i[2893] , \i[2894] ,
    \i[2895] , \i[2896] , \i[2897] , \i[2898] , \i[2899] , \i[2900] ,
    \i[2901] , \i[2902] , \i[2903] , \i[2904] , \i[2905] , \i[2906] ,
    \i[2907] , \i[2908] , \i[2909] , \i[2910] , \i[2911] , \i[2912] ,
    \i[2913] , \i[2914] , \i[2915] , \i[2916] , \i[2917] , \i[2918] ,
    \i[2919] , \i[2920] , \i[2921] , \i[2922] , \i[2923] , \i[2924] ,
    \i[2925] , \i[2926] , \i[2927] , \i[2928] , \i[2929] , \i[2930] ,
    \i[2931] , \i[2932] , \i[2933] , \i[2934] , \i[2935] , \i[2936] ,
    \i[2937] , \i[2938] , \i[2939] , \i[2940] , \i[2941] , \i[2942] ,
    \i[2943] , \i[2944] , \i[2945] , \i[2946] , \i[2947] , \i[2948] ,
    \i[2949] , \i[2950] , \i[2951] , \i[2952] , \i[2953] , \i[2954] ,
    \i[2955] , \i[2956] , \i[2957] , \i[2958] , \i[2959] , \i[2960] ,
    \i[2961] , \i[2962] , \i[2963] , \i[2964] , \i[2965] , \i[2966] ,
    \i[2967] , \i[2968] , \i[2969] , \i[2970] , \i[2971] , \i[2972] ,
    \i[2973] , \i[2974] , \i[2975] , \i[2976] , \i[2977] , \i[2978] ,
    \i[2979] , \i[2980] , \i[2981] , \i[2982] , \i[2983] , \i[2984] ,
    \i[2985] , \i[2986] , \i[2987] , \i[2988] , \i[2989] , \i[2990] ,
    \i[2991] , \i[2992] , \i[2993] , \i[2994] , \i[2995] , \i[2996] ,
    \i[2997] , \i[2998] , \i[2999] , \i[3000] , \i[3001] , \i[3002] ,
    \i[3003] , \i[3004] , \i[3005] , \i[3006] , \i[3007] , \i[3008] ,
    \i[3009] , \i[3010] , \i[3011] , \i[3012] , \i[3013] , \i[3014] ,
    \i[3015] , \i[3016] , \i[3017] , \i[3018] , \i[3019] , \i[3020] ,
    \i[3021] , \i[3022] , \i[3023] , \i[3024] , \i[3025] , \i[3026] ,
    \i[3027] , \i[3028] , \i[3029] , \i[3030] , \i[3031] , \i[3032] ,
    \i[3033] , \i[3034] , \i[3035] , \i[3036] , \i[3037] , \i[3038] ,
    \i[3039] , \i[3040] , \i[3041] , \i[3042] , \i[3043] , \i[3044] ,
    \i[3045] , \i[3046] , \i[3047] , \i[3048] , \i[3049] , \i[3050] ,
    \i[3051] , \i[3052] , \i[3053] , \i[3054] , \i[3055] , \i[3056] ,
    \i[3057] , \i[3058] , \i[3059] , \i[3060] , \i[3061] , \i[3062] ,
    \i[3063] , \i[3064] , \i[3065] , \i[3066] , \i[3067] , \i[3068] ,
    \i[3069] , \i[3070] , \i[3071] , \i[3072] , \i[3073] , \i[3074] ,
    \i[3075] , \i[3076] , \i[3077] , \i[3078] , \i[3079] , \i[3080] ,
    \i[3081] , \i[3082] , \i[3083] , \i[3084] , \i[3085] , \i[3086] ,
    \i[3087] , \i[3088] , \i[3089] , \i[3090] , \i[3091] , \i[3092] ,
    \i[3093] , \i[3094] , \i[3095] , \i[3096] , \i[3097] , \i[3098] ,
    \i[3099] , \i[3100] , \i[3101] , \i[3102] , \i[3103] , \i[3104] ,
    \i[3105] , \i[3106] , \i[3107] , \i[3108] , \i[3109] , \i[3110] ,
    \i[3111] , \i[3112] , \i[3113] , \i[3114] , \i[3115] , \i[3116] ,
    \i[3117] , \i[3118] , \i[3119] , \i[3120] , \i[3121] , \i[3122] ,
    \i[3123] , \i[3124] , \i[3125] , \i[3126] , \i[3127] , \i[3128] ,
    \i[3129] , \i[3130] , \i[3131] , \i[3132] , \i[3133] , \i[3134] ,
    \i[3135] ;
  output \o[0] , \o[1] , \o[2] , \o[3] , \o[4] , \o[5] , \o[6] , \o[7] ,
    \o[8] , \o[9] , \o[10] , \o[11] , \o[12] , \o[13] , \o[14] , \o[15] ,
    \o[16] , \o[17] , \o[18] , \o[19] , \o[20] , \o[21] , \o[22] , \o[23] ,
    \o[24] , \o[25] , \o[26] , \o[27] , \o[28] , \o[29] , \o[30] , \o[31] ,
    \o[32] , \o[33] , \o[34] , \o[35] , \o[36] , \o[37] , \o[38] , \o[39] ,
    \o[40] , \o[41] , \o[42] , \o[43] , \o[44] , \o[45] , \o[46] , \o[47] ,
    \o[48] , \o[49] , \o[50] , \o[51] , \o[52] , \o[53] , \o[54] , \o[55] ,
    \o[56] , \o[57] , \o[58] , \o[59] , \o[60] , \o[61] , \o[62] , \o[63] ,
    \o[64] , \o[65] , \o[66] , \o[67] , \o[68] , \o[69] ;
  wire new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_,
    new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_,
    new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_,
    new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_,
    new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_,
    new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_,
    new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_,
    new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_,
    new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_,
    new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_,
    new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_,
    new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_,
    new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_,
    new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_,
    new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_,
    new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_,
    new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_,
    new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_,
    new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_,
    new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_,
    new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_,
    new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_,
    new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_,
    new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_,
    new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_,
    new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_,
    new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_,
    new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_,
    new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_,
    new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_,
    new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_,
    new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_,
    new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_,
    new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_,
    new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_,
    new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_,
    new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_,
    new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_,
    new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_,
    new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_,
    new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_,
    new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_,
    new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_,
    new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_,
    new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_,
    new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_,
    new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_,
    new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_,
    new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_,
    new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_,
    new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_,
    new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_,
    new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4469_, new_n4470_, new_n4471_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4570_, new_n4571_, new_n4572_,
    new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_, new_n4578_,
    new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_, new_n4584_,
    new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_, new_n4590_,
    new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_, new_n4596_,
    new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_, new_n4602_,
    new_n4603_, new_n4604_, new_n4605_, new_n4607_, new_n4608_, new_n4609_,
    new_n4610_, new_n4611_, new_n4612_, new_n4613_, new_n4614_, new_n4615_,
    new_n4616_, new_n4617_, new_n4618_, new_n4619_, new_n4620_, new_n4621_,
    new_n4622_, new_n4623_, new_n4624_, new_n4626_, new_n4627_, new_n4628_,
    new_n4629_, new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_, new_n5214_,
    new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_,
    new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_,
    new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_,
    new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_,
    new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_,
    new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_,
    new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_,
    new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_,
    new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_,
    new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_,
    new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_,
    new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_,
    new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_,
    new_n5293_, new_n5294_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_,
    new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_,
    new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_,
    new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_,
    new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_,
    new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_,
    new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_,
    new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_,
    new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_,
    new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_,
    new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_,
    new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_,
    new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_,
    new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_,
    new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_,
    new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_,
    new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5544_,
    new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_, new_n5550_,
    new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_, new_n5556_,
    new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_, new_n5562_,
    new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_, new_n5568_,
    new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_, new_n5574_,
    new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_, new_n5580_,
    new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_, new_n5586_,
    new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_, new_n5592_,
    new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_, new_n5598_,
    new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_, new_n5604_,
    new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_, new_n5610_,
    new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_, new_n5616_,
    new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_, new_n5622_,
    new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_, new_n5628_,
    new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_, new_n5634_,
    new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_, new_n5640_,
    new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_, new_n5646_,
    new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_, new_n5652_,
    new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_, new_n5658_,
    new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_, new_n5664_,
    new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_, new_n5670_,
    new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6033_, new_n6034_,
    new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_,
    new_n6041_, new_n6042_, new_n6043_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_,
    new_n6068_, new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_,
    new_n6074_, new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_,
    new_n6080_, new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_,
    new_n6086_, new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_,
    new_n6092_, new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_,
    new_n6098_, new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_,
    new_n6104_, new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_,
    new_n6110_, new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_,
    new_n6116_, new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_,
    new_n6122_, new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_,
    new_n6128_, new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_,
    new_n6134_, new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_,
    new_n6140_, new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_,
    new_n6146_, new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_,
    new_n6152_, new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_,
    new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_,
    new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_,
    new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_,
    new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_,
    new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_,
    new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_,
    new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_,
    new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_,
    new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_,
    new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_,
    new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_,
    new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_,
    new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_,
    new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_,
    new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_,
    new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_,
    new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_,
    new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_,
    new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_,
    new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_,
    new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_,
    new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_,
    new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_,
    new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_,
    new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_,
    new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_,
    new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_,
    new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_,
    new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_,
    new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_,
    new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_,
    new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_,
    new_n6350_, new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_,
    new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_,
    new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_,
    new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_,
    new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_,
    new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_,
    new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_,
    new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_,
    new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_,
    new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_,
    new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_,
    new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_,
    new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_,
    new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_,
    new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_,
    new_n6573_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6638_, new_n6639_, new_n6640_, new_n6641_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_,
    new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_,
    new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_,
    new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_,
    new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_,
    new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_,
    new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_,
    new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6741_, new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_,
    new_n6747_, new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_,
    new_n6753_, new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_,
    new_n6759_, new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_,
    new_n6765_, new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_,
    new_n6771_, new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_,
    new_n6777_, new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_,
    new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_,
    new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_,
    new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_,
    new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_,
    new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_,
    new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_,
    new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_,
    new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_,
    new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_,
    new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_,
    new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_,
    new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_,
    new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_,
    new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_,
    new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_,
    new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_,
    new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_,
    new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_,
    new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_,
    new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_,
    new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_,
    new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_,
    new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_,
    new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_,
    new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_,
    new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_,
    new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_,
    new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_,
    new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_,
    new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_,
    new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_,
    new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_,
    new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_,
    new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_,
    new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_,
    new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_,
    new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_,
    new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_,
    new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_,
    new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_,
    new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_,
    new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_,
    new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_,
    new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_,
    new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_,
    new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_,
    new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7131_, new_n7132_,
    new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_,
    new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_,
    new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_,
    new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_,
    new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_,
    new_n7163_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7181_, new_n7182_,
    new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_,
    new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_,
    new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7662_,
    new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_,
    new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_,
    new_n7675_, new_n7676_, new_n7677_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_,
    new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_,
    new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_,
    new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_,
    new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_,
    new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_,
    new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_,
    new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_,
    new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_,
    new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_,
    new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_,
    new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_,
    new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_,
    new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_,
    new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_,
    new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_,
    new_n8009_, new_n8010_, new_n8011_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_, new_n8677_,
    new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8683_, new_n8684_,
    new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_,
    new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_,
    new_n8697_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8708_, new_n8709_, new_n8710_,
    new_n8711_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_, new_n8766_,
    new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_,
    new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_,
    new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_,
    new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_,
    new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_,
    new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_,
    new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_,
    new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_,
    new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_,
    new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_,
    new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_,
    new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_,
    new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_,
    new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_,
    new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_,
    new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_,
    new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_,
    new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_,
    new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9183_, new_n9184_,
    new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_,
    new_n9191_, new_n9193_, new_n9194_, new_n9195_, new_n9196_;
  assign \o[0]  = new_n3209_ ? (new_n3764_ ^ new_n3783_) : (~new_n3764_ ^ new_n3783_);
  assign new_n3209_ = new_n3210_ ? (~new_n3723_ ^ new_n3746_) : (new_n3723_ ^ new_n3746_);
  assign new_n3210_ = new_n3211_ ? (~new_n3653_ ^ new_n3699_) : (new_n3653_ ^ new_n3699_);
  assign new_n3211_ = new_n3212_ ? (new_n3481_ ^ new_n3642_) : (~new_n3481_ ^ new_n3642_);
  assign new_n3212_ = new_n3213_ ? (new_n3329_ ^ new_n3464_) : (~new_n3329_ ^ new_n3464_);
  assign new_n3213_ = new_n3214_ ? (~new_n3296_ ^ new_n3315_) : (new_n3296_ ^ new_n3315_);
  assign new_n3214_ = new_n3215_ ? (~new_n3245_ ^ new_n3270_) : (new_n3245_ ^ new_n3270_);
  assign new_n3215_ = new_n3243_ ? new_n3216_ : new_n3231_;
  assign new_n3216_ = new_n3229_ ? (~new_n3226_ & (new_n3230_ | ~new_n3227_ | ~\i[763] )) : new_n3217_;
  assign new_n3217_ = (~\i[1043]  & (new_n3225_ | ~\i[1042] )) ? new_n3222_ : new_n3218_;
  assign new_n3218_ = (~new_n3221_ | ~new_n3219_) & (~\i[1880]  | ~\i[1881]  | ~\i[1882]  | ~\i[1883]  | new_n3219_);
  assign new_n3219_ = new_n3220_ & (~\i[1757]  | ~\i[1756] );
  assign new_n3220_ = ~\i[1758]  & ~\i[1759] ;
  assign new_n3221_ = ~\i[1503]  & ~\i[1502]  & ~\i[1500]  & ~\i[1501] ;
  assign new_n3222_ = new_n3223_ ? new_n3224_ : (\i[607]  | (\i[605]  & \i[606] ));
  assign new_n3223_ = ~\i[2279]  & ~\i[2278]  & ~\i[2276]  & ~\i[2277] ;
  assign new_n3224_ = ~\i[2383]  & (~\i[2381]  | ~\i[2382]  | ~\i[2380] );
  assign new_n3225_ = ~\i[1040]  & ~\i[1041] ;
  assign new_n3226_ = \i[935]  & \i[934]  & \i[933]  & \i[932]  & ~new_n3227_ & new_n3228_;
  assign new_n3227_ = ~\i[1527]  & (~\i[1525]  | ~\i[1526]  | ~\i[1524] );
  assign new_n3228_ = ~\i[1723]  & (~\i[1721]  | ~\i[1722]  | ~\i[1720] );
  assign new_n3229_ = ~\i[975]  & ~\i[974]  & ~\i[972]  & ~\i[973] ;
  assign new_n3230_ = ~\i[1822]  & ~\i[1823]  & (~\i[1821]  | ~\i[1820] );
  assign new_n3231_ = (\i[2515]  & (\i[2514]  | (\i[2512]  & \i[2513] ))) ? new_n3237_ : new_n3232_;
  assign new_n3232_ = (~new_n3233_ | ~new_n3236_ | (\i[1546]  & \i[1547] )) & (~new_n3235_ | ~\i[1546]  | ~\i[1547] );
  assign new_n3233_ = new_n3234_ & ~\i[1504]  & ~\i[1505] ;
  assign new_n3234_ = ~\i[1506]  & ~\i[1507] ;
  assign new_n3235_ = ~\i[1515]  & (~\i[1514]  | (~\i[1513]  & ~\i[1512] ));
  assign new_n3236_ = \i[1167]  & \i[1166]  & \i[1164]  & \i[1165] ;
  assign new_n3237_ = new_n3238_ ? ~new_n3242_ : (new_n3240_ ? ~new_n3239_ : ~new_n3241_);
  assign new_n3238_ = ~\i[1519]  & ~\i[1518]  & ~\i[1516]  & ~\i[1517] ;
  assign new_n3239_ = \i[1303]  & \i[1301]  & \i[1302] ;
  assign new_n3240_ = \i[2063]  & \i[2062]  & \i[2060]  & \i[2061] ;
  assign new_n3241_ = \i[1711]  & (\i[1710]  | \i[1709] );
  assign new_n3242_ = ~\i[935]  & ~\i[934]  & ~\i[932]  & ~\i[933] ;
  assign new_n3243_ = new_n3244_ & (~\i[1521]  | ~\i[1520] );
  assign new_n3244_ = ~\i[1522]  & ~\i[1523] ;
  assign new_n3245_ = ~new_n3246_ & (~new_n3253_ | ((new_n3262_ | new_n3267_ | ~new_n3269_) & (new_n3255_ | new_n3269_)));
  assign new_n3246_ = ~new_n3247_ & ~new_n3253_ & (new_n3249_ | \i[955]  | ~new_n3254_ | ~new_n3251_);
  assign new_n3247_ = new_n3248_ & ((~\i[1709]  & ~\i[1710]  & ~\i[1711]  & \i[1503] ) | (new_n3250_ & ~\i[1503] ));
  assign new_n3248_ = ~\i[1759]  & (new_n3249_ | \i[955] ) & (~\i[1758]  | (~\i[1756]  & ~\i[1757] ));
  assign new_n3249_ = \i[953]  & \i[954] ;
  assign new_n3250_ = ~\i[491]  & (~\i[490]  | (~\i[489]  & ~\i[488] ));
  assign new_n3251_ = ~new_n3252_ & ~\i[1923]  & (~\i[1922]  | ~\i[1921] );
  assign new_n3252_ = ~\i[1587]  & ~\i[1586]  & ~\i[1584]  & ~\i[1585] ;
  assign new_n3253_ = ~\i[1659]  & ~\i[1658]  & ~\i[1656]  & ~\i[1657] ;
  assign new_n3254_ = ~\i[2287]  & ~\i[2286]  & ~\i[2284]  & ~\i[2285] ;
  assign new_n3255_ = new_n3259_ ? new_n3256_ : ((~new_n3261_ | ~new_n3260_) & (~\i[1086]  | ~\i[1087]  | new_n3260_));
  assign new_n3256_ = new_n3257_ ? (~\i[1427]  & (~\i[1424]  | ~\i[1425]  | ~\i[1426] )) : ~new_n3258_;
  assign new_n3257_ = ~\i[1643]  & ~\i[1642]  & ~\i[1640]  & ~\i[1641] ;
  assign new_n3258_ = ~\i[1515]  & ~\i[1514]  & ~\i[1512]  & ~\i[1513] ;
  assign new_n3259_ = ~\i[1535]  & ~\i[1534]  & ~\i[1532]  & ~\i[1533] ;
  assign new_n3260_ = ~\i[1635]  & (~\i[1633]  | ~\i[1634]  | ~\i[1632] );
  assign new_n3261_ = ~\i[2859]  & ~\i[2858]  & ~\i[2856]  & ~\i[2857] ;
  assign new_n3262_ = ~new_n3266_ & ((new_n3265_ & (~\i[1268]  | ~\i[1269] )) ? ~\i[1615]  : ~new_n3263_);
  assign new_n3263_ = new_n3264_ & (~\i[2389]  | ~\i[2388] );
  assign new_n3264_ = ~\i[2390]  & ~\i[2391] ;
  assign new_n3265_ = ~\i[1270]  & ~\i[1271] ;
  assign new_n3266_ = \i[1167]  & \i[1165]  & \i[1166] ;
  assign new_n3267_ = new_n3266_ & new_n3268_ & ((~\i[1616]  & ~\i[1617] ) | ~\i[1619]  | ~\i[1618] );
  assign new_n3268_ = ~\i[2719]  & ~\i[2718]  & ~\i[2716]  & ~\i[2717] ;
  assign new_n3269_ = ~\i[1610]  & ~\i[1611] ;
  assign new_n3270_ = ~new_n3279_ & (new_n3271_ | new_n3291_ | new_n3290_);
  assign new_n3271_ = new_n3276_ & (new_n3277_ ? (\i[1291]  | new_n3278_) : new_n3272_);
  assign new_n3272_ = new_n3274_ ? ~new_n3273_ : ~new_n3275_;
  assign new_n3273_ = \i[1615]  & \i[1614]  & \i[1612]  & \i[1613] ;
  assign new_n3274_ = ~\i[1659]  & ~\i[1657]  & ~\i[1658] ;
  assign new_n3275_ = ~\i[1847]  & ~\i[1846]  & ~\i[1844]  & ~\i[1845] ;
  assign new_n3276_ = \i[1175]  & (\i[1173]  | \i[1174]  | \i[1172] );
  assign new_n3277_ = \i[1971]  & \i[1969]  & \i[1970] ;
  assign new_n3278_ = \i[1507]  & \i[1506]  & \i[1504]  & \i[1505] ;
  assign new_n3279_ = new_n3290_ & ((\i[1607]  & (~new_n3288_ | new_n3286_)) | (~new_n3280_ & ~new_n3283_ & ~\i[1607] ));
  assign new_n3280_ = new_n3282_ & new_n3281_ & (\i[1667]  | (\i[1664]  & \i[1665]  & \i[1666] ));
  assign new_n3281_ = ~\i[1859]  & ~\i[1858]  & ~\i[1856]  & ~\i[1857] ;
  assign new_n3282_ = ~\i[491]  & ~\i[490]  & ~\i[488]  & ~\i[489] ;
  assign new_n3283_ = ~new_n3284_ & ~\i[1667]  & new_n3285_ & (~\i[1666]  | ~\i[1665]  | ~\i[1664] );
  assign new_n3284_ = ~\i[2539]  & ~\i[2538]  & ~\i[2536]  & ~\i[2537] ;
  assign new_n3285_ = ~\i[2630]  & ~\i[2631]  & (~\i[2629]  | ~\i[2628] );
  assign new_n3286_ = ~\i[1155]  & ~\i[1154]  & ~new_n3287_ & ~\i[1153] ;
  assign new_n3287_ = \i[2058]  & \i[2059] ;
  assign new_n3288_ = new_n3289_ & ~\i[1936]  & ~\i[1937] ;
  assign new_n3289_ = ~\i[1938]  & ~\i[1939] ;
  assign new_n3290_ = ~\i[1634]  & ~\i[1635] ;
  assign new_n3291_ = ~new_n3276_ & ~new_n3295_ & (new_n3292_ ? ~new_n3294_ : ~new_n3293_);
  assign new_n3292_ = \i[499]  & (\i[498]  | (\i[497]  & \i[496] ));
  assign new_n3293_ = \i[2047]  & \i[2046]  & \i[2044]  & \i[2045] ;
  assign new_n3294_ = \i[2635]  & \i[2634]  & \i[2632]  & \i[2633] ;
  assign new_n3295_ = \i[883]  & (\i[881]  | \i[882]  | \i[880] );
  assign new_n3296_ = (new_n3297_ | \i[1622]  | \i[1623] ) & (new_n3313_ | new_n3314_ | ~new_n3312_ | (~\i[1622]  & ~\i[1623] ));
  assign new_n3297_ = (new_n3298_ | ~new_n3310_) & (new_n3311_ | ~new_n3307_ | new_n3310_);
  assign new_n3298_ = (new_n3303_ | (new_n3305_ ? ~new_n3304_ : new_n3306_)) & (~new_n3301_ | new_n3299_ | ~new_n3303_);
  assign new_n3299_ = ~\i[623]  & new_n3300_;
  assign new_n3300_ = ~\i[622]  & ~\i[620]  & ~\i[621] ;
  assign new_n3301_ = new_n3302_ & ~\i[2072]  & ~\i[2073] ;
  assign new_n3302_ = ~\i[2074]  & ~\i[2075] ;
  assign new_n3303_ = ~\i[1179]  & ~\i[1178]  & ~\i[1176]  & ~\i[1177] ;
  assign new_n3304_ = \i[1099]  & (\i[1097]  | \i[1098]  | \i[1096] );
  assign new_n3305_ = ~\i[1727]  & ~\i[1725]  & ~\i[1726] ;
  assign new_n3306_ = ~\i[2091]  & (~\i[2090]  | ~\i[2089] );
  assign new_n3307_ = ~new_n3308_ & ~\i[2526]  & ~\i[2527]  & (~\i[2525]  | ~\i[2524] );
  assign new_n3308_ = new_n3309_ & (~\i[1073]  | ~\i[1072] );
  assign new_n3309_ = ~\i[1074]  & ~\i[1075] ;
  assign new_n3310_ = ~\i[1967]  & (~\i[1966]  | ~\i[1965] );
  assign new_n3311_ = ~\i[1823]  & ~\i[1821]  & ~\i[1822] ;
  assign new_n3312_ = \i[1287]  & (\i[1286]  | \i[1285] );
  assign new_n3313_ = ~\i[867]  & ~\i[866]  & ~\i[864]  & ~\i[865] ;
  assign new_n3314_ = \i[2307]  & \i[2306]  & \i[2304]  & \i[2305] ;
  assign new_n3315_ = (new_n3316_ | new_n3326_) & (new_n3328_ | \i[2423]  | ~new_n3327_ | ~new_n3238_ | ~new_n3326_);
  assign new_n3316_ = (new_n3317_ | ~new_n3323_) & (new_n3324_ | ~new_n3325_ | ~\i[979]  | new_n3323_);
  assign new_n3317_ = new_n3319_ ? new_n3318_ : (new_n3321_ ? new_n3322_ : new_n3320_);
  assign new_n3318_ = ~\i[1435]  & ~\i[1434]  & ~\i[1432]  & ~\i[1433] ;
  assign new_n3319_ = \i[514]  & \i[515]  & (\i[513]  | \i[512] );
  assign new_n3320_ = \i[1979]  & (\i[1978]  | (\i[1977]  & \i[1976] ));
  assign new_n3321_ = \i[1607]  & (\i[1605]  | \i[1606]  | \i[1604] );
  assign new_n3322_ = ~\i[1827]  & ~\i[1826]  & ~\i[1824]  & ~\i[1825] ;
  assign new_n3323_ = ~\i[1515]  & (~\i[1514]  | ~\i[1513] );
  assign new_n3324_ = ~\i[2055]  & (~\i[2054]  | (~\i[2053]  & ~\i[2052] ));
  assign new_n3325_ = ~\i[1523]  & ~\i[1521]  & ~\i[1522] ;
  assign new_n3326_ = \i[1863]  & \i[1862]  & \i[1860]  & \i[1861] ;
  assign new_n3327_ = \i[1395]  & (\i[1394]  | (\i[1393]  & \i[1392] ));
  assign new_n3328_ = \i[2422]  & \i[2420]  & \i[2421] ;
  assign new_n3329_ = new_n3330_ ? (new_n3410_ ^ new_n3456_) : (~new_n3410_ ^ new_n3456_);
  assign new_n3330_ = new_n3331_ ? (~new_n3357_ ^ new_n3380_) : (new_n3357_ ^ new_n3380_);
  assign new_n3331_ = new_n3356_ ? new_n3332_ : (new_n3345_ | (~new_n3353_ & ~new_n3352_ & new_n3355_));
  assign new_n3332_ = (~new_n3341_ & ~new_n3337_ & (\i[2518]  | \i[2519] )) | (~\i[2518]  & ~\i[2519]  & ~new_n3333_ & ~new_n3343_);
  assign new_n3333_ = new_n3334_ & (~new_n3335_ | (\i[1494]  & \i[1495]  & (\i[1493]  | \i[1492] )));
  assign new_n3334_ = new_n3336_ & (new_n3335_ | (\i[1847]  & (\i[1846]  | \i[1845] )));
  assign new_n3335_ = \i[2199]  & (\i[2197]  | \i[2198]  | \i[2196] );
  assign new_n3336_ = \i[2383]  & (\i[2382]  | \i[2381] );
  assign new_n3337_ = ~new_n3338_ & ((new_n3340_ & (~\i[1828]  | ~\i[1829] )) ? ~\i[1275]  : ~new_n3323_);
  assign new_n3338_ = new_n3339_ & (~\i[2053]  | ~\i[2052] );
  assign new_n3339_ = ~\i[2054]  & ~\i[2055] ;
  assign new_n3340_ = ~\i[1830]  & ~\i[1831] ;
  assign new_n3341_ = new_n3338_ & (new_n3342_ | ~\i[2042]  | ~\i[2043]  | (~\i[2041]  & ~\i[2040] ));
  assign new_n3342_ = ~\i[1203]  & ~\i[1201]  & ~\i[1202] ;
  assign new_n3343_ = ~new_n3336_ & ~new_n3344_ & (\i[1499]  | \i[1498] );
  assign new_n3344_ = \i[1891]  & \i[1890]  & \i[1888]  & \i[1889] ;
  assign new_n3345_ = new_n3352_ & (new_n3348_ ? new_n3346_ : (new_n3350_ ? ~new_n3349_ : new_n3351_));
  assign new_n3346_ = (~new_n3347_ & (~\i[1773]  | ~\i[1774]  | ~\i[1775] )) | (~\i[607]  & \i[1773]  & \i[1774]  & \i[1775] );
  assign new_n3347_ = ~\i[1607]  & ~\i[1605]  & ~\i[1606] ;
  assign new_n3348_ = \i[1594]  & \i[1595] ;
  assign new_n3349_ = \i[835]  & \i[834]  & \i[832]  & \i[833] ;
  assign new_n3350_ = ~\i[1871]  & ~\i[1869]  & ~\i[1870] ;
  assign new_n3351_ = ~\i[1755]  & ~\i[1754]  & ~\i[1752]  & ~\i[1753] ;
  assign new_n3352_ = ~\i[1326]  & ~\i[1327]  & (~\i[1325]  | ~\i[1324] );
  assign new_n3353_ = \i[1531]  ? \i[1211]  : new_n3354_;
  assign new_n3354_ = \i[2751]  & (\i[2750]  | (\i[2749]  & \i[2748] ));
  assign new_n3355_ = ~\i[383]  & ~\i[382]  & ~\i[380]  & ~\i[381] ;
  assign new_n3356_ = ~\i[1551]  & (~\i[1550]  | ~\i[1549] );
  assign new_n3357_ = new_n3379_ ? new_n3358_ : new_n3370_;
  assign new_n3358_ = ~new_n3359_ & (new_n3368_ | new_n3369_ | ~new_n3366_ | ~new_n3367_);
  assign new_n3359_ = ~new_n3366_ & (new_n3364_ ? (new_n3365_ | new_n3311_) : new_n3360_);
  assign new_n3360_ = new_n3362_ ? new_n3363_ : ~new_n3361_;
  assign new_n3361_ = \i[1059]  & \i[1057]  & \i[1058] ;
  assign new_n3362_ = ~\i[2219]  & (~\i[2218]  | ~\i[2217] );
  assign new_n3363_ = \i[1723]  & \i[1722]  & \i[1720]  & \i[1721] ;
  assign new_n3364_ = ~\i[2767]  & ~\i[2766]  & ~\i[2764]  & ~\i[2765] ;
  assign new_n3365_ = \i[2083]  & \i[2082]  & \i[2080]  & \i[2081] ;
  assign new_n3366_ = ~\i[963]  & (~\i[962]  | ~\i[961] );
  assign new_n3367_ = ~\i[2071]  & (~\i[2070]  | (~\i[2069]  & ~\i[2068] ));
  assign new_n3368_ = ~\i[1291]  & ~\i[1290]  & ~\i[1288]  & ~\i[1289] ;
  assign new_n3369_ = ~\i[983]  & ~\i[982]  & ~\i[980]  & ~\i[981] ;
  assign new_n3370_ = (new_n3374_ | new_n3371_ | ~\i[2051] ) & (new_n3376_ | ~new_n3377_ | ~new_n3378_ | \i[2051] );
  assign new_n3371_ = ~new_n3372_ & (~new_n3373_ | (~\i[1318]  & ~\i[1319]  & (~\i[1317]  | ~\i[1316] )));
  assign new_n3372_ = \i[2511]  & (\i[2510]  | \i[2509] );
  assign new_n3373_ = \i[1079]  & \i[1078]  & \i[1076]  & \i[1077] ;
  assign new_n3374_ = new_n3372_ & ~\i[839]  & ~new_n3375_ & ~\i[838] ;
  assign new_n3375_ = ~\i[1087]  & (~\i[1086]  | ~\i[1085] );
  assign new_n3376_ = new_n3290_ & ~\i[1632]  & ~\i[1633] ;
  assign new_n3377_ = ~\i[611]  & ~\i[610]  & ~\i[608]  & ~\i[609] ;
  assign new_n3378_ = \i[507]  & \i[506]  & \i[504]  & \i[505] ;
  assign new_n3379_ = ~\i[1631]  & (~\i[1629]  | ~\i[1630]  | ~\i[1628] );
  assign new_n3380_ = new_n3408_ ? new_n3390_ : ((new_n3403_ | new_n3407_ | ~new_n3409_) & (new_n3381_ | new_n3409_));
  assign new_n3381_ = (new_n3382_ & (~\i[2389]  | ~\i[2390]  | ~\i[2391] )) | (new_n3386_ & \i[2389]  & \i[2390]  & \i[2391] );
  assign new_n3382_ = (~new_n3385_ & (~\i[1384]  | ~\i[1385]  | ~\i[1386]  | ~\i[1387] )) | (~new_n3383_ & \i[1384]  & \i[1385]  & \i[1386]  & \i[1387] );
  assign new_n3383_ = new_n3384_ & (~\i[1525]  | ~\i[1524] );
  assign new_n3384_ = ~\i[1526]  & ~\i[1527] ;
  assign new_n3385_ = \i[991]  & \i[990]  & \i[988]  & \i[989] ;
  assign new_n3386_ = new_n3388_ ? ~new_n3389_ : ~new_n3387_;
  assign new_n3387_ = \i[1083]  & (\i[1082]  | (\i[1081]  & \i[1080] ));
  assign new_n3388_ = \i[1939]  & \i[1938]  & \i[1936]  & \i[1937] ;
  assign new_n3389_ = \i[1635]  & \i[1634]  & \i[1632]  & \i[1633] ;
  assign new_n3390_ = new_n3394_ ? (~new_n3391_ & (new_n3396_ | ~new_n3392_ | ~new_n3402_)) : ~new_n3398_;
  assign new_n3391_ = ~new_n3392_ & \i[1863]  & (\i[2267]  | (\i[2266]  & (\i[2265]  | \i[2264] )));
  assign new_n3392_ = new_n3393_ & ~\i[1704]  & ~\i[1705] ;
  assign new_n3393_ = ~\i[1706]  & ~\i[1707] ;
  assign new_n3394_ = new_n3395_ & ~\i[1716]  & ~\i[1717] ;
  assign new_n3395_ = ~\i[1718]  & ~\i[1719] ;
  assign new_n3396_ = ~\i[1711]  & ~new_n3397_ & ~\i[1710] ;
  assign new_n3397_ = \i[1708]  & \i[1709] ;
  assign new_n3398_ = ~new_n3399_ & ((\i[1519]  & ~new_n3400_ & (\i[1518]  | \i[1517] )) | (new_n3401_ & new_n3400_));
  assign new_n3399_ = ~\i[2283]  & ~\i[2282]  & ~\i[2280]  & ~\i[2281] ;
  assign new_n3400_ = ~\i[1083]  & ~\i[1082]  & ~\i[1080]  & ~\i[1081] ;
  assign new_n3401_ = ~\i[979]  & ~\i[978]  & ~\i[976]  & ~\i[977] ;
  assign new_n3402_ = ~\i[1727]  & (~\i[1725]  | ~\i[1726]  | ~\i[1724] );
  assign new_n3403_ = new_n3406_ & (~new_n3404_ | (~\i[1735]  & (~\i[1734]  | ~\i[1733] )));
  assign new_n3404_ = new_n3405_ & (\i[1713]  | \i[1712] );
  assign new_n3405_ = \i[1714]  & \i[1715] ;
  assign new_n3406_ = \i[2395]  & \i[2394]  & \i[2392]  & \i[2393] ;
  assign new_n3407_ = ~new_n3406_ & ((~\i[2253]  & ~\i[2252] ) | ~\i[2255]  | ~\i[2254] );
  assign new_n3408_ = ~\i[1739]  & ~\i[1737]  & ~\i[1738] ;
  assign new_n3409_ = ~\i[1546]  & ~\i[1547] ;
  assign new_n3410_ = new_n3411_ ^ new_n3433_;
  assign new_n3411_ = (~new_n3432_ | (new_n3325_ ? new_n3412_ : new_n3419_)) & (new_n3424_ | new_n3429_ | new_n3432_);
  assign new_n3412_ = (~new_n3313_ | ~new_n3415_ | new_n3413_) & (new_n3418_ | ~new_n3417_ | ~new_n3413_);
  assign new_n3413_ = new_n3414_ & ~\i[1604]  & ~\i[1605] ;
  assign new_n3414_ = ~\i[1606]  & ~\i[1607] ;
  assign new_n3415_ = new_n3416_ & ~\i[968]  & ~\i[969] ;
  assign new_n3416_ = ~\i[970]  & ~\i[971] ;
  assign new_n3417_ = ~\i[1599]  & (~\i[1598]  | (~\i[1597]  & ~\i[1596] ));
  assign new_n3418_ = ~\i[1615]  & (~\i[1613]  | ~\i[1614]  | ~\i[1612] );
  assign new_n3419_ = (~new_n3423_ | ~\i[737]  | ~\i[738]  | ~\i[739]  | new_n3422_) & (new_n3420_ | ~new_n3422_);
  assign new_n3420_ = (~new_n3421_ | \i[2059] ) & (\i[2626]  | \i[2627]  | ~\i[2059] );
  assign new_n3421_ = \i[1935]  & (\i[1933]  | \i[1934]  | \i[1932] );
  assign new_n3422_ = \i[1063]  & (\i[1061]  | \i[1062]  | \i[1060] );
  assign new_n3423_ = ~\i[1518]  & ~\i[1519]  & (~\i[1517]  | ~\i[1516] );
  assign new_n3424_ = ~new_n3409_ & (new_n3425_ | (~new_n3427_ & (new_n3428_ | ~new_n3295_)));
  assign new_n3425_ = new_n3427_ & (~new_n3426_ | (\i[1278]  & (\i[1277]  | \i[1276] )));
  assign new_n3426_ = ~\i[1279]  & ((~\i[1741]  & ~\i[1740] ) | ~\i[1743]  | ~\i[1742] );
  assign new_n3427_ = \i[863]  & \i[861]  & \i[862] ;
  assign new_n3428_ = \i[959]  & \i[958]  & \i[956]  & \i[957] ;
  assign new_n3429_ = new_n3409_ & (new_n3430_ | ~new_n3431_ | ~\i[1538]  | ~\i[1539] );
  assign new_n3430_ = \i[1443]  & \i[1442]  & \i[1440]  & \i[1441] ;
  assign new_n3431_ = \i[2166]  & \i[2167] ;
  assign new_n3432_ = ~\i[1739]  & ~\i[1738]  & ~\i[1736]  & ~\i[1737] ;
  assign new_n3433_ = (~new_n3454_ | (new_n3455_ ? new_n3434_ : new_n3440_)) & (new_n3444_ | new_n3449_ | new_n3454_);
  assign new_n3434_ = (~new_n3439_ | ~new_n3438_ | (~\i[2171]  & (~\i[2169]  | ~\i[2170] ))) & (new_n3435_ | new_n3438_);
  assign new_n3435_ = (~new_n3436_ & new_n3437_) | (~\i[2611]  & ~new_n3437_ & (~\i[2610]  | ~\i[2609] ));
  assign new_n3436_ = ~\i[1315]  & ~\i[1313]  & ~\i[1314] ;
  assign new_n3437_ = ~\i[1959]  & ~\i[1958]  & ~\i[1956]  & ~\i[1957] ;
  assign new_n3438_ = ~\i[2050]  & ~\i[2051] ;
  assign new_n3439_ = ~\i[1443]  & ~\i[1442]  & ~\i[1440]  & ~\i[1441] ;
  assign new_n3440_ = (\i[2051]  & (\i[2050]  | (\i[2048]  & \i[2049] ))) ? new_n3441_ : ~new_n3443_;
  assign new_n3441_ = (~\i[2458]  & ~\i[2459]  & ~new_n3442_) | (new_n3442_ & (~\i[1423]  | ~\i[1422] ));
  assign new_n3442_ = \i[1179]  & \i[1177]  & \i[1178] ;
  assign new_n3443_ = \i[1442]  & \i[1443]  & (\i[1441]  | \i[1440] );
  assign new_n3444_ = new_n3445_ & ((~new_n3446_ & new_n3447_) | (~new_n3448_ & ~\i[1663]  & ~new_n3447_));
  assign new_n3445_ = ~\i[1743]  & ~\i[1742]  & ~\i[1740]  & ~\i[1741] ;
  assign new_n3446_ = ~\i[743]  & ~\i[742]  & ~\i[740]  & ~\i[741] ;
  assign new_n3447_ = ~\i[2159]  & ~\i[2158]  & ~\i[2156]  & ~\i[2157] ;
  assign new_n3448_ = ~\i[1846]  & ~\i[1847]  & (~\i[1845]  | ~\i[1844] );
  assign new_n3449_ = ~new_n3445_ & (new_n3451_ ? new_n3453_ : (~new_n3452_ | ~new_n3450_));
  assign new_n3450_ = ~\i[1635]  & (~\i[1634]  | (~\i[1633]  & ~\i[1632] ));
  assign new_n3451_ = \i[1291]  & \i[1289]  & \i[1290] ;
  assign new_n3452_ = \i[1287]  & (\i[1286]  | (\i[1285]  & \i[1284] ));
  assign new_n3453_ = ~\i[2155]  & (~\i[2154]  | (~\i[2153]  & ~\i[2152] ));
  assign new_n3454_ = ~\i[1434]  & ~\i[1435]  & (~\i[1433]  | ~\i[1432] );
  assign new_n3455_ = ~\i[1631]  & ~\i[1630]  & ~\i[1628]  & ~\i[1629] ;
  assign new_n3456_ = ~\i[1743]  & ((new_n3284_ & (new_n3460_ | new_n3457_)) | (~new_n3462_ & new_n3463_ & ~new_n3284_));
  assign new_n3457_ = ~new_n3459_ & ~new_n3458_ & ~\i[2323]  & (~\i[2322]  | (~\i[2320]  & ~\i[2321] ));
  assign new_n3458_ = \i[1299]  & (\i[1297]  | \i[1298]  | \i[1296] );
  assign new_n3459_ = ~\i[2167]  & ~\i[2165]  & ~\i[2166] ;
  assign new_n3460_ = ~new_n3461_ & new_n3458_ & (~\i[2407]  | (~\i[2406]  & (~\i[2405]  | ~\i[2404] )));
  assign new_n3461_ = ~\i[1715]  & (~\i[1714]  | ~\i[1713] );
  assign new_n3462_ = ~\i[2635]  & ~\i[2634]  & ~\i[2632]  & ~\i[2633] ;
  assign new_n3463_ = \i[938]  & \i[939]  & (\i[2287]  | \i[2286] );
  assign new_n3464_ = new_n3480_ ? (new_n3479_ ? ~new_n3472_ : ~new_n3465_) : new_n3475_;
  assign new_n3465_ = new_n3418_ ? ((new_n3471_ | new_n3470_) & (~\i[390]  | ~\i[391]  | ~new_n3470_)) : new_n3466_;
  assign new_n3466_ = (~\i[855]  & (~\i[854]  | (~\i[852]  & ~\i[853] ))) ? ~new_n3469_ : new_n3467_;
  assign new_n3467_ = new_n3468_ & ~\i[2056]  & ~\i[2057] ;
  assign new_n3468_ = ~\i[2058]  & ~\i[2059] ;
  assign new_n3469_ = \i[2290]  & \i[2291]  & (\i[2289]  | \i[2288] );
  assign new_n3470_ = ~\i[1711]  & (~\i[1710]  | ~new_n3397_);
  assign new_n3471_ = \i[2086]  & \i[2087]  & (\i[2085]  | \i[2084] );
  assign new_n3472_ = (~new_n3474_ | new_n3473_) & (\i[1966]  | \i[1967]  | ~new_n3473_);
  assign new_n3473_ = ~\i[1747]  & ~\i[1746]  & ~\i[1744]  & ~\i[1745] ;
  assign new_n3474_ = \i[2394]  & \i[2395]  & ((\i[1088]  & \i[1089] ) | \i[1091]  | \i[1090] );
  assign new_n3475_ = (new_n3478_ | new_n3476_) & (new_n3477_ | \i[2497]  | \i[2498]  | \i[2499]  | ~new_n3476_);
  assign new_n3476_ = ~\i[955]  & (~\i[954]  | (~\i[953]  & ~\i[952] ));
  assign new_n3477_ = \i[2162]  & \i[2163] ;
  assign new_n3478_ = ~\i[1639]  & (~\i[1638]  | (~\i[1637]  & ~\i[1636] ));
  assign new_n3479_ = \i[1607]  & (\i[1606]  | \i[1605] );
  assign new_n3480_ = ~\i[1591]  & ~\i[1589]  & ~\i[1590] ;
  assign new_n3481_ = new_n3482_ ? (~new_n3598_ ^ new_n3620_) : (new_n3598_ ^ new_n3620_);
  assign new_n3482_ = new_n3483_ ? (~new_n3551_ ^ new_n3589_) : (new_n3551_ ^ new_n3589_);
  assign new_n3483_ = new_n3484_ ? (~new_n3507_ ^ new_n3529_) : (new_n3507_ ^ new_n3529_);
  assign new_n3484_ = new_n3506_ ? new_n3485_ : new_n3500_;
  assign new_n3485_ = (new_n3499_ & (\i[1188]  | \i[1189] )) ? new_n3486_ : new_n3493_;
  assign new_n3486_ = (\i[2383]  & (\i[2380]  | \i[2381]  | \i[2382] )) ? new_n3487_ : new_n3489_;
  assign new_n3487_ = (new_n3488_ & (~\i[1637]  | ~\i[1638]  | ~\i[1639] )) | (\i[2207]  & \i[1637]  & \i[1638]  & \i[1639] );
  assign new_n3488_ = new_n3393_ & (~\i[1705]  | ~\i[1704] );
  assign new_n3489_ = (new_n3491_ & ~\i[2641] ) ? new_n3490_ : (~new_n3492_ | (~\i[940]  & ~\i[941] ));
  assign new_n3490_ = \i[1383]  & \i[1381]  & \i[1382] ;
  assign new_n3491_ = ~\i[2642]  & ~\i[2643] ;
  assign new_n3492_ = \i[942]  & \i[943] ;
  assign new_n3493_ = (new_n3494_ | (new_n3495_ ? new_n3369_ : ~new_n3496_)) & (~new_n3497_ | ~new_n3498_ | ~new_n3494_);
  assign new_n3494_ = ~\i[627]  & ~\i[626]  & ~\i[624]  & ~\i[625] ;
  assign new_n3495_ = ~\i[1087]  & ~\i[1085]  & ~\i[1086] ;
  assign new_n3496_ = ~\i[1190]  & ~\i[1191]  & (~\i[1189]  | ~\i[1188] );
  assign new_n3497_ = ~\i[831]  & (~\i[829]  | ~\i[830]  | ~\i[828] );
  assign new_n3498_ = \i[2386]  & \i[2387]  & (\i[2385]  | \i[2384] );
  assign new_n3499_ = \i[1190]  & \i[1191] ;
  assign new_n3500_ = (~\i[1925]  & ~\i[1926]  & ~\i[1927] ) ? (new_n3503_ | new_n3505_) : new_n3501_;
  assign new_n3501_ = ~new_n3502_ & ~\i[755]  & (~\i[754]  | ~\i[753] );
  assign new_n3502_ = ~\i[1423]  & ~\i[1421]  & ~\i[1422] ;
  assign new_n3503_ = new_n3504_ & (~\i[861]  | ~\i[860] );
  assign new_n3504_ = ~\i[862]  & ~\i[863] ;
  assign new_n3505_ = ~\i[1934]  & ~\i[1935]  & (~\i[1933]  | ~\i[1932] );
  assign new_n3506_ = ~\i[1214]  & ~\i[1215]  & (~\i[1213]  | ~\i[1212] );
  assign new_n3507_ = new_n3528_ ? new_n3522_ : ((new_n3519_ | new_n3514_ | ~new_n3527_) & (new_n3508_ | new_n3527_));
  assign new_n3508_ = (new_n3513_ | new_n3509_) & (new_n3511_ | ~new_n3512_ | ~new_n3509_);
  assign new_n3509_ = new_n3510_ & ~\i[2528]  & ~\i[2529] ;
  assign new_n3510_ = ~\i[2530]  & ~\i[2531] ;
  assign new_n3511_ = ~\i[1175]  & ~\i[1174]  & ~\i[1172]  & ~\i[1173] ;
  assign new_n3512_ = ~\i[2731]  & ~\i[2730]  & ~\i[2728]  & ~\i[2729] ;
  assign new_n3513_ = ~\i[1883]  & ~\i[1881]  & ~\i[1882] ;
  assign new_n3514_ = new_n3515_ & (new_n3516_ ? ~new_n3517_ : ~new_n3518_);
  assign new_n3515_ = \i[1299]  & (\i[1298]  | \i[1297] );
  assign new_n3516_ = ~\i[1947]  & (~\i[1945]  | ~\i[1946]  | ~\i[1944] );
  assign new_n3517_ = \i[946]  & \i[947]  & (\i[945]  | \i[944] );
  assign new_n3518_ = \i[1607]  & (\i[1606]  | (\i[1605]  & \i[1604] ));
  assign new_n3519_ = new_n3521_ & ~new_n3515_ & ~new_n3520_;
  assign new_n3520_ = ~\i[2067]  & (~\i[2066]  | ~\i[2065] );
  assign new_n3521_ = ~\i[939]  & ~\i[937]  & ~\i[938] ;
  assign new_n3522_ = (new_n3523_ | ~new_n3524_) & (new_n3525_ | ~new_n3405_ | ~new_n3526_ | new_n3524_);
  assign new_n3523_ = ~\i[2627]  & ~\i[2626]  & ~\i[2624]  & ~\i[2625] ;
  assign new_n3524_ = \i[2067]  & (\i[2066]  | (\i[2065]  & \i[2064] ));
  assign new_n3525_ = \i[1615]  & (\i[1613]  | \i[1614]  | \i[1612] );
  assign new_n3526_ = \i[1712]  & \i[1713] ;
  assign new_n3527_ = ~\i[1967]  & (~\i[1965]  | ~\i[1966]  | ~\i[1964] );
  assign new_n3528_ = \i[1523]  & (\i[1522]  | \i[1521] );
  assign new_n3529_ = (new_n3530_ | new_n3537_ | ~new_n3243_) & (new_n3243_ | (~new_n3547_ & (new_n3541_ | new_n3550_)));
  assign new_n3530_ = ~new_n3534_ & ((new_n3531_ & new_n3535_) | (~new_n3536_ & new_n3369_ & ~new_n3535_));
  assign new_n3531_ = new_n3532_ ? ~new_n3533_ : (\i[399]  | (\i[397]  & \i[398] ));
  assign new_n3532_ = ~\i[2399]  & ~\i[2397]  & ~\i[2398] ;
  assign new_n3533_ = ~\i[2079]  & (~\i[2078]  | ~\i[2077] );
  assign new_n3534_ = \i[2194]  & \i[2195] ;
  assign new_n3535_ = ~\i[1175]  & (~\i[1174]  | (~\i[1173]  & ~\i[1172] ));
  assign new_n3536_ = \i[1411]  & (\i[1409]  | \i[1410]  | \i[1408] );
  assign new_n3537_ = new_n3534_ & (\i[2411]  | ~\i[1551]  | new_n3538_) & (new_n3540_ | new_n3257_ | ~new_n3538_);
  assign new_n3538_ = \i[1393]  & new_n3539_ & \i[1392] ;
  assign new_n3539_ = \i[1394]  & \i[1395] ;
  assign new_n3540_ = ~\i[850]  & ~\i[851] ;
  assign new_n3541_ = new_n3545_ ? new_n3542_ : (~new_n3546_ | (\i[754]  & \i[755] ));
  assign new_n3542_ = (\i[2523]  & (\i[2520]  | \i[2521]  | \i[2522] )) ? ~new_n3544_ : ~new_n3543_;
  assign new_n3543_ = \i[971]  & \i[970]  & \i[968]  & \i[969] ;
  assign new_n3544_ = ~\i[1627]  & ~\i[1625]  & ~\i[1626] ;
  assign new_n3545_ = ~\i[751]  & ~\i[749]  & ~\i[750] ;
  assign new_n3546_ = \i[2295]  & \i[2294]  & \i[2292]  & \i[2293] ;
  assign new_n3547_ = new_n3550_ & new_n3548_ & new_n3294_;
  assign new_n3548_ = new_n3549_ & ~\i[1508]  & ~\i[1509] ;
  assign new_n3549_ = ~\i[1510]  & ~\i[1511] ;
  assign new_n3550_ = ~\i[1174]  & ~\i[1175]  & (~\i[1173]  | ~\i[1172] );
  assign new_n3551_ = new_n3552_ ? (new_n3566_ ^ new_n3577_) : (~new_n3566_ ^ new_n3577_);
  assign new_n3552_ = ~new_n3558_ & (~new_n3563_ | (~new_n3561_ & ~new_n3553_ & ~\i[1214]  & ~\i[1215] ));
  assign new_n3553_ = new_n3554_ & (\i[2523]  | ~new_n3555_ | (\i[2522]  & (\i[2520]  | \i[2521] )));
  assign new_n3554_ = ~new_n3557_ & (new_n3555_ | \i[1588]  | \i[1589]  | \i[1590]  | \i[1591] );
  assign new_n3555_ = new_n3556_ & ~\i[1296]  & ~\i[1297] ;
  assign new_n3556_ = ~\i[1298]  & ~\i[1299] ;
  assign new_n3557_ = ~\i[1199]  & ~\i[1197]  & ~\i[1198] ;
  assign new_n3558_ = new_n3559_ & (\i[2620]  | \i[2621]  | \i[2622]  | \i[2623] );
  assign new_n3559_ = \i[1302]  & \i[1303]  & \i[1635]  & (~new_n3560_ | (~\i[1512]  & ~\i[1513] ));
  assign new_n3560_ = \i[1514]  & \i[1515] ;
  assign new_n3561_ = new_n3557_ & ((~new_n3562_ & ~new_n3462_) | (\i[1527]  & new_n3462_ & (\i[1526]  | \i[1525] )));
  assign new_n3562_ = \i[1534]  & \i[1535]  & (\i[1533]  | \i[1532] );
  assign new_n3563_ = ~\i[1635]  & ((~\i[1214]  & ~\i[1215] ) | \i[755]  | (new_n3564_ & ~new_n3565_));
  assign new_n3564_ = ~\i[1727]  & ~\i[1726]  & ~\i[1724]  & ~\i[1725] ;
  assign new_n3565_ = \i[1543]  & (\i[1542]  | \i[1541] );
  assign new_n3566_ = new_n3282_ & ((~new_n3571_ & ~new_n3576_) | (~new_n3567_ & new_n3310_ & new_n3576_));
  assign new_n3567_ = (~new_n3570_ & new_n3568_) | (~\i[1815]  & ~new_n3568_ & (~\i[1814]  | ~\i[1813] ));
  assign new_n3568_ = \i[949]  & new_n3569_ & \i[948] ;
  assign new_n3569_ = \i[950]  & \i[951] ;
  assign new_n3570_ = ~\i[1975]  & ~\i[1973]  & ~\i[1974] ;
  assign new_n3571_ = (new_n3534_ | new_n3572_ | ~new_n3523_) & (new_n3523_ | (new_n3574_ ? new_n3573_ : new_n3575_));
  assign new_n3572_ = ~\i[2295]  & ~\i[2294]  & ~\i[2292]  & ~\i[2293] ;
  assign new_n3573_ = ~\i[1935]  & ~\i[1933]  & ~\i[1934] ;
  assign new_n3574_ = ~\i[1947]  & ~\i[1945]  & ~\i[1946] ;
  assign new_n3575_ = \i[1630]  & \i[1631]  & (\i[1629]  | \i[1628] );
  assign new_n3576_ = ~\i[2283]  & ~\i[2281]  & ~\i[2282] ;
  assign new_n3577_ = new_n3586_ ? new_n3578_ : (new_n3588_ ? new_n3587_ : new_n3585_);
  assign new_n3578_ = (new_n3583_ | ~new_n3584_ | ~new_n3582_ | (~\i[835]  & ~\i[834] )) & (new_n3579_ | new_n3582_);
  assign new_n3579_ = (~new_n3580_ | new_n3515_) & (new_n3581_ | ~new_n3515_ | (\i[639]  & (\i[637]  | \i[638] )));
  assign new_n3580_ = ~\i[1955]  & (~\i[1485]  | ~\i[1486]  | ~\i[1487]  | ~\i[1484] );
  assign new_n3581_ = ~\i[1839]  & (~\i[1838]  | ~\i[1837] );
  assign new_n3582_ = ~\i[2395]  & ~\i[2393]  & ~\i[2394] ;
  assign new_n3583_ = \i[2078]  & \i[2079]  & (\i[2077]  | \i[2076] );
  assign new_n3584_ = \i[1059]  & \i[1058]  & \i[1056]  & \i[1057] ;
  assign new_n3585_ = new_n3504_ & ~\i[860]  & ~\i[861] ;
  assign new_n3586_ = ~\i[1663]  & (~\i[1662]  | (~\i[1661]  & ~\i[1660] ));
  assign new_n3587_ = ~\i[1327]  & ~\i[1326]  & ~\i[1324]  & ~\i[1325] ;
  assign new_n3588_ = ~\i[607]  & ~\i[605]  & ~\i[606] ;
  assign new_n3589_ = new_n3597_ ? new_n3590_ : (~new_n3596_ | (~\i[1820]  & ~\i[1821]  & ~\i[1822] ));
  assign new_n3590_ = (~new_n3593_ | ~new_n3594_) & (new_n3591_ | ~new_n3595_ | new_n3594_);
  assign new_n3591_ = ~\i[1658]  & ~\i[1659]  & new_n3592_ & (~\i[1657]  | ~\i[1656] );
  assign new_n3592_ = ~\i[1647]  & ~\i[1646]  & ~\i[1644]  & ~\i[1645] ;
  assign new_n3593_ = ~\i[1059]  & ~\i[1058]  & ~\i[1056]  & ~\i[1057] ;
  assign new_n3594_ = \i[1851]  & \i[1849]  & \i[1850] ;
  assign new_n3595_ = ~\i[411]  & ~\i[410]  & ~\i[408]  & ~\i[409] ;
  assign new_n3596_ = \i[1823]  & \i[2530]  & \i[2531]  & (\i[1995]  | (\i[1993]  & \i[1994] ));
  assign new_n3597_ = ~\i[711]  & ~\i[709]  & ~\i[710] ;
  assign new_n3598_ = new_n3473_ ? new_n3599_ : ((~new_n3610_ & new_n3278_) | (~new_n3612_ & ~new_n3617_ & ~new_n3278_));
  assign new_n3599_ = \i[2071]  ? new_n3600_ : ((~new_n3605_ & ~new_n3607_) | (~new_n3608_ & new_n3609_ & new_n3607_));
  assign new_n3600_ = new_n3253_ ? (~new_n3604_ & (~new_n3492_ | ~\i[940]  | ~\i[941] )) : new_n3601_;
  assign new_n3601_ = (~new_n3602_ & \i[1206]  & \i[1207]  & (\i[1204]  | \i[1205] )) | (new_n3603_ & (~\i[1206]  | ~\i[1207]  | (~\i[1204]  & ~\i[1205] )));
  assign new_n3602_ = \i[1175]  & (\i[1174]  | (\i[1173]  & \i[1172] ));
  assign new_n3603_ = \i[723]  & \i[722]  & \i[720]  & \i[721] ;
  assign new_n3604_ = \i[2743]  & (\i[2742]  | (\i[2741]  & \i[2740] ));
  assign new_n3605_ = new_n3303_ ? ~new_n3606_ : (\i[815]  & (\i[812]  | \i[813]  | \i[814] ));
  assign new_n3606_ = ~\i[1263]  & ~\i[1262]  & ~\i[1260]  & ~\i[1261] ;
  assign new_n3607_ = ~\i[599]  & ~\i[597]  & ~\i[598] ;
  assign new_n3608_ = \i[979]  & (\i[978]  | \i[977] );
  assign new_n3609_ = \i[1403]  & \i[1401]  & \i[1402] ;
  assign new_n3610_ = (~\i[1630]  | ~\i[1631]  | (~\i[718]  & ~\i[719] )) & \i[1287]  & (~new_n3611_ | \i[718]  | \i[719] );
  assign new_n3611_ = ~\i[851]  & (~\i[850]  | (~\i[849]  & ~\i[848] ));
  assign new_n3612_ = new_n3616_ & ((~new_n3615_ & ~new_n3613_) | (~\i[1843]  & new_n3613_ & (~\i[1840]  | ~new_n3614_)));
  assign new_n3613_ = ~\i[2419]  & ~\i[2418]  & ~\i[2416]  & ~\i[2417] ;
  assign new_n3614_ = \i[1841]  & \i[1842] ;
  assign new_n3615_ = ~\i[1158]  & ~\i[1159] ;
  assign new_n3616_ = \i[2047]  & (\i[2046]  | \i[2045] );
  assign new_n3617_ = new_n3618_ & ~new_n3616_ & ~new_n3619_;
  assign new_n3618_ = ~\i[1847]  & ~\i[1845]  & ~\i[1846] ;
  assign new_n3619_ = ~\i[2059]  & ~\i[2057]  & ~\i[2058] ;
  assign new_n3620_ = new_n3641_ ? new_n3621_ : ((~\i[1770]  & ~\i[1771]  & new_n3640_) | (~new_n3635_ & ~new_n3640_));
  assign new_n3621_ = ~new_n3622_ & (~new_n3626_ | (~new_n3629_ & ~new_n3634_) | (~new_n3632_ & new_n3634_));
  assign new_n3622_ = ~new_n3626_ & (new_n3627_ ? (~\i[1307]  | ~new_n3628_) : new_n3623_);
  assign new_n3623_ = new_n3513_ ? ~new_n3624_ : new_n3625_;
  assign new_n3624_ = ~\i[1955]  & ~\i[1953]  & ~\i[1954] ;
  assign new_n3625_ = ~\i[1970]  & ~\i[1971] ;
  assign new_n3626_ = ~\i[1875]  & (~\i[1874]  | (~\i[1873]  & ~\i[1872] ));
  assign new_n3627_ = ~\i[931]  & ~\i[930]  & ~\i[928]  & ~\i[929] ;
  assign new_n3628_ = ~\i[967]  & ~\i[966]  & ~\i[964]  & ~\i[965] ;
  assign new_n3629_ = (new_n3630_ | new_n3631_) & (\i[2514]  | \i[2515]  | ~new_n3631_ | (\i[2513]  & \i[2512] ));
  assign new_n3630_ = \i[2614]  & \i[2615]  & (\i[2613]  | \i[2612] );
  assign new_n3631_ = \i[731]  & (\i[729]  | \i[730]  | \i[728] );
  assign new_n3632_ = (new_n3633_ | new_n3241_) & (~\i[1978]  | ~\i[1979]  | ~new_n3241_);
  assign new_n3633_ = \i[1723]  & (\i[1722]  | \i[1721] );
  assign new_n3634_ = ~\i[2631]  & ~\i[2629]  & ~\i[2630] ;
  assign new_n3635_ = (new_n3636_ | (~\i[1975]  & (~\i[1972]  | ~\i[1974]  | ~\i[1973] ))) & (\i[1974]  | \i[1973]  | ~new_n3639_ | \i[1975] );
  assign new_n3636_ = ~new_n3637_ & ~new_n3638_;
  assign new_n3637_ = ~\i[1431]  & ~\i[1429]  & ~\i[1430] ;
  assign new_n3638_ = ~\i[2298]  & ~\i[2299] ;
  assign new_n3639_ = ~\i[823]  & ~\i[821]  & ~\i[822] ;
  assign new_n3640_ = new_n3438_ & (~\i[2049]  | ~\i[2048] );
  assign new_n3641_ = ~\i[1851]  & ~\i[1849]  & ~\i[1850] ;
  assign new_n3642_ = (new_n3641_ | (~new_n3643_ & (new_n3647_ | new_n3648_))) & (new_n3652_ | ~new_n3651_ | ~new_n3641_);
  assign new_n3643_ = new_n3647_ & (~new_n3646_ | ~new_n3644_) & (~\i[1701]  | ~\i[1702]  | ~\i[1703] );
  assign new_n3644_ = new_n3645_ & ~\i[1404]  & ~\i[1405] ;
  assign new_n3645_ = ~\i[1406]  & ~\i[1407] ;
  assign new_n3646_ = \i[1398]  & \i[1399] ;
  assign new_n3647_ = ~\i[2051]  & (~\i[2050]  | (~\i[2049]  & ~\i[2048] ));
  assign new_n3648_ = ~new_n3649_ & ((\i[2393]  & \i[2394]  & \i[2395] ) | ~\i[1315]  | new_n3650_);
  assign new_n3649_ = ~new_n3275_ & ~\i[1315]  & ((~\i[1320]  & ~\i[1321] ) | ~\i[1323]  | ~\i[1322] );
  assign new_n3650_ = ~\i[847]  & (~\i[846]  | (~\i[845]  & ~\i[844] ));
  assign new_n3651_ = ~\i[2643]  & ~\i[1543]  & ~\i[1542]  & ~\i[1331]  & ~\i[1329]  & ~\i[1330] ;
  assign new_n3652_ = ~\i[2543]  & ~\i[2542]  & ~\i[2540]  & ~\i[2541] ;
  assign new_n3653_ = new_n3654_ ? (~new_n3673_ ^ new_n3692_) : (new_n3673_ ^ new_n3692_);
  assign new_n3654_ = (\i[1703]  & (\i[1700]  | \i[1701]  | \i[1702] )) ? new_n3671_ : new_n3655_;
  assign new_n3655_ = new_n3670_ ? new_n3656_ : (new_n3669_ ? new_n3665_ : new_n3662_);
  assign new_n3656_ = (new_n3661_ | ~new_n3660_ | (\i[2042]  & \i[2043] )) & (~\i[2042]  | ~\i[2043]  | ~new_n3657_ | ~new_n3645_);
  assign new_n3657_ = ~new_n3658_ & new_n3659_ & (~\i[1405]  | ~\i[1404] );
  assign new_n3658_ = \i[612]  & \i[613] ;
  assign new_n3659_ = ~\i[614]  & ~\i[615] ;
  assign new_n3660_ = ~\i[2614]  & ~\i[2615]  & (~\i[2613]  | ~\i[2612] );
  assign new_n3661_ = ~\i[618]  & ~\i[619]  & (~\i[617]  | ~\i[616] );
  assign new_n3662_ = new_n3663_ ? ~new_n3630_ : ~new_n3664_;
  assign new_n3663_ = ~\i[991]  & ~\i[990]  & ~\i[988]  & ~\i[989] ;
  assign new_n3664_ = ~\i[1951]  & (~\i[1950]  | ~\i[1949] );
  assign new_n3665_ = new_n3666_ ? (\i[1071]  | (new_n3667_ & \i[1070] )) : ~new_n3668_;
  assign new_n3666_ = ~\i[2503]  & (~\i[2501]  | ~\i[2502]  | ~\i[2500] );
  assign new_n3667_ = \i[1068]  & \i[1069] ;
  assign new_n3668_ = ~\i[935]  & ~\i[933]  & ~\i[934] ;
  assign new_n3669_ = ~\i[2043]  & ~\i[2042]  & ~\i[2040]  & ~\i[2041] ;
  assign new_n3670_ = ~\i[1942]  & ~\i[1943] ;
  assign new_n3671_ = ~\i[1885]  & ~\i[1886]  & ~\i[1887]  & (new_n3672_ | new_n3606_);
  assign new_n3672_ = ~\i[2382]  & ~\i[2383]  & (~\i[2381]  | ~\i[2380] );
  assign new_n3673_ = new_n3691_ ? new_n3678_ : ((~new_n3674_ | ~new_n3690_) & (new_n3685_ | new_n3688_ | new_n3690_));
  assign new_n3674_ = (new_n3676_ | ~new_n3677_ | ~\i[2172]  | \i[1195] ) & (~new_n3312_ | ~new_n3675_ | ~\i[1195] );
  assign new_n3675_ = new_n3328_ & \i[2423] ;
  assign new_n3676_ = \i[1439]  & \i[1437]  & \i[1438] ;
  assign new_n3677_ = \i[2175]  & \i[2173]  & \i[2174] ;
  assign new_n3678_ = new_n3684_ ? new_n3679_ : ((~new_n3681_ & ~new_n3683_ & new_n3682_) | (~new_n3258_ & ~new_n3682_));
  assign new_n3679_ = (~\i[1206]  & ~\i[1207] ) ? new_n3680_ : ~\i[2163] ;
  assign new_n3680_ = \i[1518]  & \i[1519]  & (\i[1517]  | \i[1516] );
  assign new_n3681_ = \i[863]  & (\i[862]  | \i[861] );
  assign new_n3682_ = \i[1603]  & \i[1602]  & \i[1600]  & \i[1601] ;
  assign new_n3683_ = ~\i[1614]  & ~\i[1615] ;
  assign new_n3684_ = \i[975]  & \i[974]  & \i[972]  & \i[973] ;
  assign new_n3685_ = ~new_n3686_ & ~\i[2059]  & new_n3687_ & (~\i[2058]  | ~\i[2057]  | ~\i[2056] );
  assign new_n3686_ = \i[1971]  & (\i[1970]  | (\i[1969]  & \i[1968] ));
  assign new_n3687_ = ~\i[1931]  & ~\i[1930]  & ~\i[1928]  & ~\i[1929] ;
  assign new_n3688_ = new_n3686_ & (~new_n3689_ | new_n3234_) & (~\i[2381]  | ~\i[2382]  | ~\i[2383]  | ~new_n3234_);
  assign new_n3689_ = ~\i[1743]  & ~\i[1741]  & ~\i[1742] ;
  assign new_n3690_ = \i[962]  & \i[963]  & (\i[961]  | \i[960] );
  assign new_n3691_ = \i[1519]  & (\i[1517]  | \i[1518]  | \i[1516] );
  assign new_n3692_ = (\i[1511]  & (\i[1508]  | \i[1509]  | \i[1510] )) ? ~new_n3698_ : new_n3693_;
  assign new_n3693_ = ~new_n3694_ & (~new_n3697_ | ~new_n3437_ | ~new_n3696_ | (~\i[2519]  & ~\i[2518] ));
  assign new_n3694_ = ~new_n3437_ & ~new_n3695_ & (\i[1652]  | \i[1653]  | \i[1654]  | \i[1655] );
  assign new_n3695_ = ~\i[1195]  & (~\i[1193]  | ~\i[1194]  | ~\i[1192] );
  assign new_n3696_ = ~\i[2071]  & ~\i[2070]  & ~\i[2068]  & ~\i[2069] ;
  assign new_n3697_ = ~\i[599]  & ~\i[598]  & ~\i[596]  & ~\i[597] ;
  assign new_n3698_ = \i[863]  & \i[862]  & \i[2279]  & (~\i[1519]  | ~\i[1518]  | ~\i[1517] );
  assign new_n3699_ = (~new_n3691_ & (new_n3607_ ? new_n3706_ : new_n3700_)) | (~new_n3712_ & ~new_n3718_ & new_n3691_);
  assign new_n3700_ = (new_n3701_ | new_n3704_) & (new_n3702_ | new_n3705_ | ~new_n3704_);
  assign new_n3701_ = (~\i[1891]  | ~new_n3540_ | (~\i[1890]  & (~\i[1888]  | ~\i[1889] ))) & (new_n3392_ | new_n3540_);
  assign new_n3702_ = ~new_n3703_ & ~\i[2099]  & (~\i[2098]  | ~\i[2097] );
  assign new_n3703_ = ~\i[1167]  & ~\i[1165]  & ~\i[1166] ;
  assign new_n3704_ = \i[839]  & (\i[838]  | (\i[837]  & \i[836] ));
  assign new_n3705_ = (~\i[1379]  | ~\i[1377]  | ~\i[1378] ) & (\i[2099]  | (\i[2098]  & \i[2097] ));
  assign new_n3706_ = new_n3707_ ? new_n3709_ : new_n3711_;
  assign new_n3707_ = ~\i[1963]  & (~\i[1962]  | ~new_n3708_);
  assign new_n3708_ = \i[1960]  & \i[1961] ;
  assign new_n3709_ = (~\i[2659]  & (~\i[2656]  | ~\i[2657]  | ~\i[2658] )) ? ~new_n3710_ : new_n3362_;
  assign new_n3710_ = ~\i[2863]  & ~\i[2862]  & ~\i[2860]  & ~\i[2861] ;
  assign new_n3711_ = ~\i[2275]  & ~\i[2273]  & ~\i[2274] ;
  assign new_n3712_ = \i[1713]  & \i[1714]  & \i[1715]  & (new_n3716_ ? new_n3713_ : new_n3717_);
  assign new_n3713_ = (new_n3714_ | new_n3715_) & (\i[1662]  | \i[1663]  | ~new_n3715_);
  assign new_n3714_ = \i[730]  & \i[731]  & (\i[729]  | \i[728] );
  assign new_n3715_ = ~\i[2626]  & ~\i[2627]  & (~\i[2625]  | ~\i[2624] );
  assign new_n3716_ = \i[2051]  & (\i[2049]  | \i[2050]  | \i[2048] );
  assign new_n3717_ = \i[1283]  & \i[1281]  & \i[1282] ;
  assign new_n3718_ = new_n3721_ & (new_n3719_ | ~new_n3684_ | (\i[1767]  & (\i[1765]  | \i[1766] )));
  assign new_n3719_ = new_n3720_ & \i[1183] ;
  assign new_n3720_ = \i[1181]  & \i[1182] ;
  assign new_n3721_ = (~\i[1713]  | ~\i[1714]  | ~\i[1715] ) & (new_n3258_ | new_n3684_ | new_n3722_);
  assign new_n3722_ = \i[1547]  & \i[1546]  & \i[1544]  & \i[1545] ;
  assign new_n3723_ = (~new_n3724_ & ~new_n3745_) | (~new_n3732_ & ~new_n3738_ & new_n3745_);
  assign new_n3724_ = new_n3729_ ? ((~new_n3727_ | ~new_n3730_) & (new_n3731_ | ~new_n3327_ | new_n3730_)) : ~new_n3725_;
  assign new_n3725_ = new_n3677_ & new_n3726_ & ~\i[1631]  & ~\i[1629]  & ~\i[1630] ;
  assign new_n3726_ = \i[958]  & \i[959]  & (\i[957]  | \i[956] );
  assign new_n3727_ = \i[2275]  & \i[2274]  & new_n3728_ & \i[2273] ;
  assign new_n3728_ = \i[1482]  & \i[1483] ;
  assign new_n3729_ = \i[2395]  & (\i[2394]  | (\i[2393]  & \i[2392] ));
  assign new_n3730_ = ~\i[1831]  & ~\i[1829]  & ~\i[1830] ;
  assign new_n3731_ = \i[1627]  & \i[1625]  & \i[1626] ;
  assign new_n3732_ = new_n3310_ & (new_n3737_ ? new_n3733_ : (~new_n3735_ | (~\i[1066]  & ~\i[1067] )));
  assign new_n3733_ = ~\i[2635]  & new_n3734_ & (~\i[2634]  | ~\i[2633] );
  assign new_n3734_ = ~\i[2658]  & ~\i[2659]  & (~\i[2657]  | ~\i[2656] );
  assign new_n3735_ = new_n3736_ & ~\i[516]  & ~\i[517] ;
  assign new_n3736_ = ~\i[518]  & ~\i[519] ;
  assign new_n3737_ = ~\i[1295]  & (~\i[1294]  | ~\i[1293] );
  assign new_n3738_ = ~new_n3310_ & (new_n3741_ ? ~new_n3739_ : (new_n3743_ ? new_n3744_ : new_n3742_));
  assign new_n3739_ = new_n3740_ & (\i[1667]  | (\i[1666]  & (\i[1665]  | \i[1664] )));
  assign new_n3740_ = \i[1167]  & (\i[1166]  | (\i[1165]  & \i[1164] ));
  assign new_n3741_ = ~\i[1287]  & (~\i[1286]  | ~\i[1285] );
  assign new_n3742_ = ~\i[2503]  & (~\i[2502]  | (~\i[2501]  & ~\i[2500] ));
  assign new_n3743_ = \i[1495]  & (\i[1493]  | \i[1494]  | \i[1492] );
  assign new_n3744_ = ~\i[1319]  & ~\i[1317]  & ~\i[1318] ;
  assign new_n3745_ = ~\i[1635]  & ~\i[1633]  & ~\i[1634] ;
  assign new_n3746_ = new_n3641_ ? (new_n3763_ ? new_n3758_ : new_n3752_) : new_n3747_;
  assign new_n3747_ = (~new_n3750_ | ~new_n3748_ | new_n3647_) & (new_n3751_ | ~new_n3293_ | ~new_n3539_ | ~new_n3647_);
  assign new_n3748_ = new_n3749_ & \i[1435]  & (\i[1434]  | \i[1433]  | \i[1432] );
  assign new_n3749_ = \i[746]  & \i[747]  & (\i[745]  | \i[744] );
  assign new_n3750_ = ~\i[1071]  & (~\i[1070]  | (~\i[1069]  & ~\i[1068] ));
  assign new_n3751_ = \i[1775]  & \i[1774]  & \i[1772]  & \i[1773] ;
  assign new_n3752_ = (~new_n3755_ | ~new_n3753_) & (new_n3756_ | ~new_n3757_ | new_n3753_);
  assign new_n3753_ = new_n3754_ & (\i[1069]  | \i[1068] );
  assign new_n3754_ = \i[1070]  & \i[1071] ;
  assign new_n3755_ = ~\i[602]  & ~\i[603]  & new_n3244_ & (~\i[601]  | ~\i[600] );
  assign new_n3756_ = ~\i[1503]  & ~\i[1501]  & ~\i[1502] ;
  assign new_n3757_ = \i[539]  & \i[538]  & \i[536]  & \i[537] ;
  assign new_n3758_ = (~new_n3762_ | ~\i[2070]  | ~\i[2071]  | ~new_n3759_) & (new_n3759_ | (new_n3761_ & ~new_n3760_));
  assign new_n3759_ = \i[1723]  & (\i[1721]  | \i[1722]  | \i[1720] );
  assign new_n3760_ = ~\i[1182]  & ~\i[1183]  & (~\i[1181]  | ~\i[1180] );
  assign new_n3761_ = ~\i[1711]  & ~\i[1710]  & ~\i[1708]  & ~\i[1709] ;
  assign new_n3762_ = \i[1763]  & (\i[1761]  | \i[1762]  | \i[1760] );
  assign new_n3763_ = ~\i[1515]  & ~\i[1513]  & ~\i[1514] ;
  assign new_n3764_ = new_n3432_ ? (new_n3763_ ? new_n3774_ : new_n3780_) : new_n3765_;
  assign new_n3765_ = (new_n3769_ | new_n3766_ | ~new_n3454_) & (new_n3749_ | new_n3772_ | ~new_n3773_ | new_n3454_);
  assign new_n3766_ = new_n3767_ & (~\i[1552]  | ~\i[1553]  | ~\i[1554]  | ~\i[1555] );
  assign new_n3767_ = ~new_n3768_ & ((~\i[2365]  & ~\i[2364] ) | ~\i[2367]  | ~\i[2366] );
  assign new_n3768_ = \i[2165]  & new_n3431_ & \i[2164] ;
  assign new_n3769_ = new_n3768_ & (new_n3770_ | ~\i[1601]  | ~\i[1602]  | ~\i[1603] );
  assign new_n3770_ = \i[1285]  & new_n3771_ & \i[1284] ;
  assign new_n3771_ = \i[1286]  & \i[1287] ;
  assign new_n3772_ = \i[1479]  & (\i[1478]  | (\i[1477]  & \i[1476] ));
  assign new_n3773_ = \i[2155]  & \i[2154]  & \i[2152]  & \i[2153] ;
  assign new_n3774_ = (new_n3777_ | new_n3778_ | new_n3696_) & (~new_n3696_ | (\i[1291]  ? new_n3779_ : ~new_n3775_));
  assign new_n3775_ = new_n3776_ & ~\i[2514]  & ~\i[2515] ;
  assign new_n3776_ = ~\i[2512]  & ~\i[2513] ;
  assign new_n3777_ = ~\i[1283]  & (~\i[1282]  | (~\i[1281]  & ~\i[1280] ));
  assign new_n3778_ = ~\i[2287]  & ~\i[2285]  & ~\i[2286] ;
  assign new_n3779_ = ~\i[975]  & ~\i[973]  & ~\i[974] ;
  assign new_n3780_ = (\i[991]  | ~new_n3676_ | new_n3781_) & (~new_n3781_ | (new_n3744_ ? \i[1519]  : ~new_n3782_));
  assign new_n3781_ = new_n3667_ & new_n3754_;
  assign new_n3782_ = ~\i[843]  & ~\i[841]  & ~\i[842] ;
  assign new_n3783_ = (new_n3784_ | new_n3445_) & (new_n3794_ | ~new_n3801_ | ~new_n3445_);
  assign new_n3784_ = (new_n3785_ | new_n3793_) & (new_n3792_ | ~new_n3793_ | (~new_n3791_ & (~\i[526]  | ~\i[527] )));
  assign new_n3785_ = (new_n3786_ | new_n3770_) & (new_n3790_ | ~new_n3789_ | ~new_n3770_);
  assign new_n3786_ = (new_n3787_ | ~new_n3788_) & (\i[1733]  | \i[1734]  | \i[1735]  | new_n3788_);
  assign new_n3787_ = ~\i[2459]  & ~\i[2458]  & ~\i[2456]  & ~\i[2457] ;
  assign new_n3788_ = ~\i[1435]  & ~\i[1433]  & ~\i[1434] ;
  assign new_n3789_ = ~\i[1738]  & ~\i[1739]  & (~\i[1737]  | ~\i[1736] );
  assign new_n3790_ = \i[1423]  & \i[1422]  & \i[1420]  & \i[1421] ;
  assign new_n3791_ = \i[1095]  & \i[1094]  & \i[1092]  & \i[1093] ;
  assign new_n3792_ = \i[2039]  & \i[2037]  & \i[2038] ;
  assign new_n3793_ = \i[1435]  & \i[1433]  & \i[1434] ;
  assign new_n3794_ = (new_n3664_ | ~new_n3800_ | new_n3795_) & (~new_n3795_ | (new_n3798_ ? ~new_n3799_ : new_n3797_));
  assign new_n3795_ = new_n3796_ & ~\i[2508]  & ~\i[2509] ;
  assign new_n3796_ = ~\i[2510]  & ~\i[2511] ;
  assign new_n3797_ = ~\i[1391]  & (~\i[1390]  | (~\i[1389]  & ~\i[1388] ));
  assign new_n3798_ = ~\i[1862]  & ~\i[1863] ;
  assign new_n3799_ = ~\i[1774]  & ~\i[1775] ;
  assign new_n3800_ = ~\i[1963]  & ~\i[1961]  & ~\i[1962] ;
  assign new_n3801_ = ~\i[1407]  & ~\i[1405]  & ~\i[1406] ;
  assign \o[1]  = new_n3803_ ? (new_n3804_ ^ new_n3805_) : (~new_n3804_ ^ new_n3805_);
  assign new_n3803_ = (~new_n3764_ & ~new_n3783_) | (~new_n3209_ & (~new_n3764_ | ~new_n3783_));
  assign new_n3804_ = (~new_n3723_ & ~new_n3746_) | (~new_n3210_ & (~new_n3723_ | ~new_n3746_));
  assign new_n3805_ = new_n3806_ ? (~new_n3807_ ^ new_n3910_) : (new_n3807_ ^ new_n3910_);
  assign new_n3806_ = (~new_n3653_ & ~new_n3699_) | (~new_n3211_ & (~new_n3653_ | ~new_n3699_));
  assign new_n3807_ = new_n3808_ ? (new_n3809_ ^ new_n3907_) : (~new_n3809_ ^ new_n3907_);
  assign new_n3808_ = (~new_n3481_ & new_n3642_) | (~new_n3212_ & (~new_n3481_ | new_n3642_));
  assign new_n3809_ = new_n3810_ ? (new_n3835_ ^ new_n3836_) : (~new_n3835_ ^ new_n3836_);
  assign new_n3810_ = new_n3811_ ? (~new_n3812_ ^ new_n3813_) : (new_n3812_ ^ new_n3813_);
  assign new_n3811_ = (~new_n3296_ & ~new_n3315_) | (~new_n3214_ & (~new_n3296_ | ~new_n3315_));
  assign new_n3812_ = (~new_n3551_ & ~new_n3589_) | (~new_n3483_ & (~new_n3551_ | ~new_n3589_));
  assign new_n3813_ = new_n3814_ ? (new_n3815_ ^ new_n3830_) : (~new_n3815_ ^ new_n3830_);
  assign new_n3814_ = (~new_n3507_ & ~new_n3529_) | (~new_n3484_ & (~new_n3507_ | ~new_n3529_));
  assign new_n3815_ = new_n3816_ ? (~new_n3822_ ^ new_n3826_) : (new_n3822_ ^ new_n3826_);
  assign new_n3816_ = new_n3356_ ? ((~\i[2518]  & ~\i[2519] ) ? ~new_n3818_ : ~new_n3817_) : new_n3819_;
  assign new_n3817_ = ~new_n3341_ & (new_n3338_ | (new_n3323_ & (~new_n3340_ | (\i[1828]  & \i[1829] ))));
  assign new_n3818_ = ~new_n3334_ & (new_n3344_ | new_n3336_);
  assign new_n3819_ = (new_n3820_ | ~new_n3352_) & (new_n3354_ | \i[1531]  | ~new_n3355_ | new_n3352_);
  assign new_n3820_ = (~new_n3821_ | ~new_n3348_) & (new_n3350_ | ~new_n3351_ | new_n3348_);
  assign new_n3821_ = \i[1775]  & \i[1774]  & ~\i[607]  & \i[1773] ;
  assign new_n3822_ = (new_n3823_ | ~new_n3290_) & (~new_n3824_ | ~new_n3277_ | ~\i[1175]  | new_n3290_);
  assign new_n3823_ = (~new_n3280_ | \i[1607] ) & (~new_n3288_ | ~new_n3287_ | ~\i[1163]  | ~\i[1607] );
  assign new_n3824_ = new_n3825_ & (\i[2511]  | (\i[2509]  & \i[2510] ));
  assign new_n3825_ = new_n3278_ & (\i[1172]  | \i[1173]  | \i[1174] );
  assign new_n3826_ = (new_n3827_ | new_n3691_) & (~new_n3829_ | ~\i[1713]  | ~\i[1714]  | ~\i[1715]  | ~new_n3691_);
  assign new_n3827_ = (~new_n3704_ | ~new_n3702_ | new_n3607_) & (new_n3707_ | ~new_n3711_ | ~new_n3828_ | ~new_n3607_);
  assign new_n3828_ = \i[1551]  & \i[1550]  & \i[1548]  & \i[1549] ;
  assign new_n3829_ = new_n3716_ & ~new_n3714_ & ~new_n3715_;
  assign new_n3830_ = new_n3831_ ^ new_n3833_;
  assign new_n3831_ = (\i[1503]  | ~new_n3248_ | ~new_n3250_ | new_n3253_) & (~new_n3269_ | ~new_n3832_ | ~new_n3253_);
  assign new_n3832_ = ~new_n3263_ & ~new_n3266_ & (~new_n3265_ | (\i[1268]  & \i[1269] ));
  assign new_n3833_ = new_n3243_ & new_n3229_ & ~new_n3834_ & ~new_n3227_ & ~new_n3228_;
  assign new_n3834_ = ~\i[2170]  & ~\i[2171]  & (~\i[2169]  | ~\i[2168] );
  assign new_n3835_ = (~new_n3329_ & new_n3464_) | (~new_n3213_ & (~new_n3329_ | new_n3464_));
  assign new_n3836_ = new_n3837_ ? (new_n3860_ ^ new_n3861_) : (~new_n3860_ ^ new_n3861_);
  assign new_n3837_ = new_n3838_ ? (~new_n3839_ ^ new_n3859_) : (new_n3839_ ^ new_n3859_);
  assign new_n3838_ = (~new_n3245_ & ~new_n3270_) | (~new_n3215_ & (~new_n3245_ | ~new_n3270_));
  assign new_n3839_ = new_n3840_ ? (~new_n3846_ ^ new_n3851_) : (new_n3846_ ^ new_n3851_);
  assign new_n3840_ = new_n3641_ ? new_n3841_ : (~new_n3844_ & (~new_n3647_ | ~new_n3751_ | ~new_n3845_));
  assign new_n3841_ = (new_n3842_ | new_n3763_) & (~new_n3843_ | ~new_n3759_ | ~new_n3763_ | (\i[2071]  & \i[2070] ));
  assign new_n3842_ = (~new_n3240_ | new_n3244_ | ~new_n3753_) & (~new_n3756_ | new_n3753_ | (~\i[1655]  & ~\i[1654] ));
  assign new_n3843_ = ~\i[814]  & ~\i[815]  & (~\i[813]  | ~\i[812] );
  assign new_n3844_ = ~new_n3750_ & ~new_n3647_ & ((~new_n3614_ & ~\i[1843] ) ? ~new_n3413_ : new_n3618_);
  assign new_n3845_ = \i[2038]  & \i[2039]  & (\i[2037]  | \i[2036] );
  assign new_n3846_ = new_n3745_ ? (new_n3310_ ? new_n3847_ : new_n3850_) : new_n3724_;
  assign new_n3847_ = (new_n3848_ | new_n3733_ | ~new_n3737_) & (~new_n3735_ | new_n3737_ | (~\i[1067]  & ~\i[1066] ));
  assign new_n3848_ = new_n3849_ & ~new_n3734_ & ~\i[2753] ;
  assign new_n3849_ = ~\i[2754]  & ~\i[2755] ;
  assign new_n3850_ = new_n3741_ ? ~new_n3739_ : (new_n3743_ ? new_n3744_ : new_n3742_);
  assign new_n3851_ = new_n3379_ ? new_n3852_ : ((~new_n3374_ | ~\i[2051] ) & (new_n3858_ | ~new_n3376_ | \i[2051] ));
  assign new_n3852_ = new_n3366_ ? ((new_n3856_ | new_n3367_) & (~new_n3854_ | ~new_n3368_ | ~new_n3367_)) : new_n3853_;
  assign new_n3853_ = (new_n3362_ | ~new_n3361_ | new_n3364_) & (new_n3311_ | new_n3365_ | ~new_n3364_);
  assign new_n3854_ = new_n3855_ & ~\i[1852]  & ~\i[1853] ;
  assign new_n3855_ = ~\i[1854]  & ~\i[1855] ;
  assign new_n3856_ = ~new_n3857_ & (~\i[1996]  | ~\i[1997]  | ~\i[1998]  | ~\i[1999] );
  assign new_n3857_ = \i[882]  & \i[883]  & (\i[881]  | \i[880] );
  assign new_n3858_ = ~\i[1431]  & ~\i[1430]  & ~\i[1428]  & ~\i[1429] ;
  assign new_n3859_ = (~new_n3357_ & ~new_n3380_) | (~new_n3331_ & (~new_n3357_ | ~new_n3380_));
  assign new_n3860_ = (~new_n3410_ & new_n3456_) | (~new_n3330_ & (~new_n3410_ | new_n3456_));
  assign new_n3861_ = new_n3862_ ? (~new_n3885_ ^ new_n3906_) : (new_n3885_ ^ new_n3906_);
  assign new_n3862_ = new_n3863_ ? (~new_n3870_ ^ new_n3876_) : (new_n3870_ ^ new_n3876_);
  assign new_n3863_ = new_n3408_ ? ((new_n3866_ | ~new_n3394_) & (new_n3398_ | new_n3868_ | new_n3394_)) : new_n3864_;
  assign new_n3864_ = ~new_n3865_ & ((~new_n3404_ & new_n3480_) | ~new_n3409_ | ~new_n3403_);
  assign new_n3865_ = \i[2391]  & \i[2390]  & \i[2389]  & new_n3388_ & ~new_n3409_ & ~new_n3389_;
  assign new_n3866_ = (\i[1863]  | ~new_n3235_ | new_n3392_) & (new_n3402_ | new_n3867_ | ~new_n3392_);
  assign new_n3867_ = ~\i[1306]  & ~\i[1307]  & (~\i[1305]  | ~\i[1304] );
  assign new_n3868_ = (~\i[1890]  | ~\i[1891]  | (\i[2498]  & \i[2499] )) & new_n3399_ & (new_n3869_ | ~\i[2498]  | ~\i[2499] );
  assign new_n3869_ = \i[1406]  & \i[1407] ;
  assign new_n3870_ = new_n3432_ ? new_n3871_ : (new_n3409_ ? ~new_n3430_ : new_n3874_);
  assign new_n3871_ = (new_n3872_ | ~new_n3325_) & (~\i[2059]  | ~new_n3422_ | new_n3325_ | (~\i[2627]  & ~\i[2626] ));
  assign new_n3872_ = (new_n3873_ | new_n3417_ | ~new_n3413_) & (new_n3413_ | (new_n3415_ ? new_n3313_ : ~new_n3710_));
  assign new_n3873_ = \i[1863]  & (\i[1861]  | \i[1862]  | \i[1860] );
  assign new_n3874_ = (new_n3427_ | ~new_n3428_ | ~new_n3383_) & (~new_n3425_ | new_n3875_);
  assign new_n3875_ = \i[1742]  & \i[1743]  & (\i[1740]  | \i[1741] ) & (\i[1642]  | \i[1643] );
  assign new_n3876_ = new_n3432_ ? (new_n3763_ ? new_n3883_ : new_n3884_) : new_n3877_;
  assign new_n3877_ = (new_n3878_ | new_n3454_) & (~new_n3770_ | ~new_n3768_ | ~new_n3882_ | ~new_n3454_);
  assign new_n3878_ = (~new_n3772_ | ~new_n3451_ | new_n3749_) & (~new_n3749_ | (new_n3879_ ? ~new_n3880_ : ~new_n3881_));
  assign new_n3879_ = ~\i[1639]  & ~\i[1638]  & ~\i[1636]  & ~\i[1637] ;
  assign new_n3880_ = ~\i[1971]  & (~\i[1969]  | ~\i[1970]  | ~\i[1968] );
  assign new_n3881_ = \i[1299]  & (\i[1298]  | (\i[1297]  & \i[1296] ));
  assign new_n3882_ = \i[2619]  & (\i[2618]  | \i[2617] );
  assign new_n3883_ = (~new_n3777_ | ~\i[1667]  | new_n3696_) & (new_n3775_ | \i[1291]  | ~new_n3696_);
  assign new_n3884_ = (~new_n3325_ | ~\i[991]  | new_n3781_) & (new_n3744_ | new_n3782_ | ~new_n3781_);
  assign new_n3885_ = ~new_n3886_ ^ new_n3900_;
  assign new_n3886_ = new_n3445_ ? new_n3887_ : ((new_n3895_ | ~new_n3793_) & (~new_n3894_ | ~new_n3790_ | new_n3793_));
  assign new_n3887_ = ~new_n3888_ & (new_n3801_ | ((new_n3891_ | new_n3889_) & (new_n3892_ | ~new_n3893_ | ~new_n3889_)));
  assign new_n3888_ = new_n3801_ & ((~new_n3799_ & new_n3798_ & new_n3795_) | (~new_n3795_ & (new_n3800_ | ~new_n3311_)));
  assign new_n3889_ = new_n3890_ & ~\i[1208]  & ~\i[1209] ;
  assign new_n3890_ = ~\i[1210]  & ~\i[1211] ;
  assign new_n3891_ = (\i[1692]  | \i[1693]  | \i[1694]  | \i[1695]  | ~new_n3754_) & (~new_n3373_ | new_n3754_);
  assign new_n3892_ = ~\i[1315]  & (~\i[1314]  | (~\i[1313]  & ~\i[1312] ));
  assign new_n3893_ = \i[1067]  & \i[1066]  & \i[1064]  & \i[1065] ;
  assign new_n3894_ = \i[1719]  & new_n3770_ & \i[1718] ;
  assign new_n3895_ = (~new_n3792_ | (new_n3897_ ? ~new_n3896_ : ~new_n3898_)) & (~new_n3791_ | new_n3899_ | new_n3792_);
  assign new_n3896_ = ~\i[2171]  & (~\i[2170]  | (~\i[2169]  & ~\i[2168] ));
  assign new_n3897_ = \i[2382]  & \i[2383] ;
  assign new_n3898_ = \i[1182]  & \i[1183] ;
  assign new_n3899_ = ~\i[635]  & ~\i[634]  & ~\i[632]  & ~\i[633] ;
  assign new_n3900_ = ~new_n3901_ & (new_n3454_ | new_n3903_);
  assign new_n3901_ = new_n3454_ & (~new_n3455_ | new_n3902_);
  assign new_n3902_ = (~new_n3437_ | new_n3436_ | new_n3438_) & (new_n3439_ | ~new_n3438_ | (~\i[1819]  & ~\i[1818] ));
  assign new_n3903_ = ~new_n3904_ & (~new_n3445_ | ((~new_n3446_ | ~new_n3447_) & (new_n3448_ | \i[1663]  | new_n3447_)));
  assign new_n3904_ = ~new_n3445_ & (~new_n3452_ | ~new_n3450_ | new_n3451_) & (~new_n3453_ | ~new_n3905_ | ~new_n3451_);
  assign new_n3905_ = ~\i[1967]  & ~\i[1966]  & ~\i[1964]  & ~\i[1965] ;
  assign new_n3906_ = new_n3411_ & new_n3433_;
  assign new_n3907_ = ~new_n3908_ ^ new_n3909_;
  assign new_n3908_ = (~new_n3598_ & ~new_n3620_) | (~new_n3482_ & (~new_n3598_ | ~new_n3620_));
  assign new_n3909_ = (~new_n3577_ & new_n3566_) | (~new_n3552_ & (~new_n3577_ | new_n3566_));
  assign new_n3910_ = (~new_n3673_ & ~new_n3692_) | (~new_n3654_ & (~new_n3673_ | ~new_n3692_));
  assign \o[2]  = ~new_n3912_ ^ new_n3913_;
  assign new_n3912_ = (~new_n3805_ & new_n3804_) | (new_n3803_ & (~new_n3805_ | new_n3804_));
  assign new_n3913_ = new_n3914_ ^ new_n3915_;
  assign new_n3914_ = (~new_n3807_ & new_n3910_) | (new_n3806_ & (~new_n3807_ | new_n3910_));
  assign new_n3915_ = new_n3916_ ? (~new_n3917_ ^ new_n3942_) : (new_n3917_ ^ new_n3942_);
  assign new_n3916_ = (~new_n3809_ & ~new_n3907_) | (new_n3808_ & (~new_n3809_ | ~new_n3907_));
  assign new_n3917_ = new_n3918_ ? (new_n3921_ ^ new_n3922_) : (~new_n3921_ ^ new_n3922_);
  assign new_n3918_ = ~new_n3919_ ^ new_n3920_;
  assign new_n3919_ = (~new_n3813_ & new_n3812_) | (new_n3811_ & (~new_n3813_ | new_n3812_));
  assign new_n3920_ = ~new_n3831_ & new_n3833_;
  assign new_n3921_ = (~new_n3836_ & new_n3835_) | (~new_n3810_ & (~new_n3836_ | new_n3835_));
  assign new_n3922_ = new_n3923_ ? (new_n3927_ ^ new_n3928_) : (~new_n3927_ ^ new_n3928_);
  assign new_n3923_ = new_n3924_ ? (new_n3925_ ^ new_n3926_) : (~new_n3925_ ^ new_n3926_);
  assign new_n3924_ = (~new_n3839_ & new_n3859_) | (new_n3838_ & (~new_n3839_ | new_n3859_));
  assign new_n3925_ = (~new_n3815_ & ~new_n3830_) | (new_n3814_ & (~new_n3815_ | ~new_n3830_));
  assign new_n3926_ = (~new_n3822_ & ~new_n3826_) | (~new_n3816_ & (~new_n3822_ | ~new_n3826_));
  assign new_n3927_ = (~new_n3861_ & new_n3860_) | (~new_n3837_ & (~new_n3861_ | new_n3860_));
  assign new_n3928_ = new_n3929_ ? (new_n3932_ ^ new_n3933_) : (~new_n3932_ ^ new_n3933_);
  assign new_n3929_ = ~new_n3930_ ^ new_n3931_;
  assign new_n3930_ = (~new_n3846_ & ~new_n3851_) | (~new_n3840_ & (~new_n3846_ | ~new_n3851_));
  assign new_n3931_ = (~new_n3870_ & ~new_n3876_) | (~new_n3863_ & (~new_n3870_ | ~new_n3876_));
  assign new_n3932_ = (~new_n3885_ & ~new_n3906_) | (~new_n3862_ & (~new_n3885_ | ~new_n3906_));
  assign new_n3933_ = ~new_n3934_ ^ new_n3935_;
  assign new_n3934_ = ~new_n3900_ & new_n3886_;
  assign new_n3935_ = ~new_n3936_ ^ new_n3941_;
  assign new_n3936_ = ~new_n3901_ & (new_n3939_ | new_n3454_ | (new_n3445_ & (new_n3938_ | new_n3937_)));
  assign new_n3937_ = new_n3447_ & (~\i[1535]  | new_n3446_) & (\i[2377]  | \i[2378]  | \i[2379]  | ~new_n3446_);
  assign new_n3938_ = new_n3448_ & ~new_n3447_ & ~\i[1415] ;
  assign new_n3939_ = ~new_n3453_ & ~new_n3445_ & new_n3451_ & (~\i[1843]  | (~\i[1840]  & new_n3940_));
  assign new_n3940_ = ~\i[1841]  & ~\i[1842] ;
  assign new_n3941_ = new_n3897_ & new_n3792_ & new_n3793_ & ~new_n3445_ & ~new_n3896_;
  assign new_n3942_ = new_n3908_ & new_n3909_;
  assign \o[3]  = ((new_n3944_ | new_n3945_) & (~new_n3946_ ^ ~new_n3947_)) | (~new_n3944_ & ~new_n3945_ & (~new_n3946_ ^ new_n3947_));
  assign new_n3944_ = ~new_n3913_ & new_n3912_;
  assign new_n3945_ = ~new_n3915_ & new_n3914_;
  assign new_n3946_ = (~new_n3917_ & new_n3942_) | (new_n3916_ & (~new_n3917_ | new_n3942_));
  assign new_n3947_ = new_n3948_ ? (~new_n3949_ ^ new_n3958_) : (new_n3949_ ^ new_n3958_);
  assign new_n3948_ = (~new_n3922_ & new_n3921_) | (~new_n3918_ & (~new_n3922_ | new_n3921_));
  assign new_n3949_ = new_n3950_ ? (~new_n3951_ ^ new_n3952_) : (new_n3951_ ^ new_n3952_);
  assign new_n3950_ = (~new_n3928_ & new_n3927_) | (~new_n3923_ & (~new_n3928_ | new_n3927_));
  assign new_n3951_ = (new_n3925_ & new_n3926_) | (new_n3924_ & (new_n3925_ | new_n3926_));
  assign new_n3952_ = new_n3953_ ? (~new_n3954_ ^ new_n3957_) : (new_n3954_ ^ new_n3957_);
  assign new_n3953_ = (~new_n3933_ & new_n3932_) | (~new_n3929_ & (~new_n3933_ | new_n3932_));
  assign new_n3954_ = new_n3955_ ^ new_n3956_;
  assign new_n3955_ = ~new_n3934_ & ~new_n3935_;
  assign new_n3956_ = new_n3936_ & new_n3941_;
  assign new_n3957_ = new_n3930_ & new_n3931_;
  assign new_n3958_ = new_n3919_ & new_n3920_;
  assign \o[4]  = ~new_n3960_ ^ new_n3961_;
  assign new_n3960_ = (new_n3946_ | (~new_n3947_ & (new_n3945_ | new_n3944_))) & (new_n3945_ | new_n3944_ | ~new_n3947_);
  assign new_n3961_ = new_n3962_ ^ new_n3963_;
  assign new_n3962_ = (~new_n3949_ & new_n3958_) | (new_n3948_ & (~new_n3949_ | new_n3958_));
  assign new_n3963_ = new_n3964_ ^ new_n3965_;
  assign new_n3964_ = (~new_n3952_ & new_n3951_) | (new_n3950_ & (~new_n3952_ | new_n3951_));
  assign new_n3965_ = new_n3966_ ^ new_n3967_;
  assign new_n3966_ = (~new_n3954_ & new_n3957_) | (new_n3953_ & (~new_n3954_ | new_n3957_));
  assign new_n3967_ = ~new_n3955_ & ~new_n3956_;
  assign \o[5]  = ((new_n3969_ | new_n3970_) & (~new_n3971_ ^ new_n3972_)) | (~new_n3969_ & ~new_n3970_ & (~new_n3971_ ^ ~new_n3972_));
  assign new_n3969_ = ~new_n3961_ & new_n3960_;
  assign new_n3970_ = ~new_n3963_ & new_n3962_;
  assign new_n3971_ = ~new_n3965_ & new_n3964_;
  assign new_n3972_ = ~new_n3967_ & new_n3966_;
  assign \o[6]  = (new_n3972_ | new_n3969_ | new_n3970_) & (new_n3971_ | (new_n3972_ & (new_n3969_ | new_n3970_)));
  assign \o[7]  = new_n3975_ ^ new_n4455_;
  assign new_n3975_ = new_n3976_ ? (new_n4420_ ^ new_n4438_) : (~new_n4420_ ^ new_n4438_);
  assign new_n3976_ = new_n3977_ ? (new_n4346_ ^ new_n4404_) : (~new_n4346_ ^ new_n4404_);
  assign new_n3977_ = new_n3978_ ? (new_n4200_ ^ new_n4319_) : (~new_n4200_ ^ new_n4319_);
  assign new_n3978_ = new_n3979_ ? (new_n4114_ ^ new_n4182_) : (~new_n4114_ ^ new_n4182_);
  assign new_n3979_ = new_n3980_ ? (new_n4051_ ^ new_n4106_) : (~new_n4051_ ^ new_n4106_);
  assign new_n3980_ = new_n3981_ ? (~new_n4003_ ^ new_n4026_) : (new_n4003_ ^ new_n4026_);
  assign new_n3981_ = (new_n3982_ & \i[1531] ) | (~new_n3991_ & ~\i[1531]  & (~new_n4001_ | new_n3999_));
  assign new_n3982_ = (\i[2497]  & \i[2498]  & \i[2499] ) ? (new_n3986_ | new_n3989_) : new_n3983_;
  assign new_n3983_ = ~new_n3984_ & (~\i[877]  | ~\i[878]  | ~\i[879] );
  assign new_n3984_ = \i[1403]  & \i[1402]  & \i[1401]  & ~new_n3985_ & \i[1400] ;
  assign new_n3985_ = new_n3798_ & ~\i[1860]  & ~\i[1861] ;
  assign new_n3986_ = ~new_n3987_ & ~new_n3988_ & ~\i[654]  & ~\i[655]  & (~\i[653]  | ~\i[652] );
  assign new_n3987_ = \i[2839]  & (\i[2838]  | \i[2837] );
  assign new_n3988_ = ~\i[735]  & ~\i[734]  & ~\i[732]  & ~\i[733] ;
  assign new_n3989_ = new_n3990_ & new_n3988_ & (\i[2379]  | \i[2378]  | \i[2377] );
  assign new_n3990_ = \i[1307]  & \i[1306]  & \i[1304]  & \i[1305] ;
  assign new_n3991_ = ~new_n3992_ & new_n3998_ & (new_n3997_ | \i[1962]  | \i[1963]  | ~new_n3993_);
  assign new_n3992_ = ~new_n3993_ & ((new_n3995_ & \i[1509] ) ? ~new_n3756_ : new_n3996_);
  assign new_n3993_ = new_n3994_ & ~\i[1836]  & ~\i[1837] ;
  assign new_n3994_ = ~\i[1838]  & ~\i[1839] ;
  assign new_n3995_ = \i[1510]  & \i[1511] ;
  assign new_n3996_ = ~\i[523]  & ~\i[522]  & ~\i[520]  & ~\i[521] ;
  assign new_n3997_ = ~\i[2631]  & ~\i[2630]  & ~\i[2628]  & ~\i[2629] ;
  assign new_n3998_ = ~\i[1199]  & ~\i[1198]  & ~\i[1196]  & ~\i[1197] ;
  assign new_n3999_ = ~\i[627]  & ~\i[626]  & ~new_n4000_ & ~\i[625] ;
  assign new_n4000_ = ~\i[754]  & ~\i[755] ;
  assign new_n4001_ = ~new_n3998_ & new_n4002_ & (~new_n4000_ | (\i[1955]  & (\i[1954]  | \i[1953] )));
  assign new_n4002_ = ~\i[951]  & ~\i[950]  & ~\i[948]  & ~\i[949] ;
  assign new_n4003_ = ~new_n4004_ & (~new_n3259_ | (~new_n4014_ & (~new_n4022_ | (~new_n4023_ & ~new_n3546_))));
  assign new_n4004_ = ~new_n3259_ & (new_n4005_ | new_n4012_) & (new_n4011_ | new_n4009_ | ~new_n4013_ | ~new_n4012_);
  assign new_n4005_ = new_n4006_ & (new_n4007_ | ~\i[2767]  | (~\i[2766]  & (~\i[2764]  | ~\i[2765] )));
  assign new_n4006_ = ~new_n4008_ & (\i[1531]  | ~new_n4007_ | (\i[1530]  & (\i[1528]  | \i[1529] )));
  assign new_n4007_ = \i[1403]  & (\i[1402]  | (\i[1401]  & \i[1400] ));
  assign new_n4008_ = \i[2483]  & \i[2482]  & \i[2480]  & \i[2481] ;
  assign new_n4009_ = ~\i[763]  & new_n4010_;
  assign new_n4010_ = \i[1943]  & (\i[1941]  | \i[1942]  | \i[1940] );
  assign new_n4011_ = ~new_n4010_ & (~\i[1643]  | (~\i[1642]  & (~\i[1641]  | ~\i[1640] )));
  assign new_n4012_ = \i[1950]  & \i[1951]  & (\i[1949]  | \i[1948] );
  assign new_n4013_ = ~\i[1055]  & ~\i[1054]  & ~\i[1052]  & ~\i[1053] ;
  assign new_n4014_ = new_n4020_ & (new_n4015_ | (~new_n4018_ & (new_n4019_ ? new_n4021_ : ~new_n3781_)));
  assign new_n4015_ = new_n4018_ & (~new_n4016_ | new_n4017_) & (new_n3708_ | \i[1962]  | \i[1963]  | ~new_n4017_);
  assign new_n4016_ = ~\i[2519]  & (~\i[2517]  | ~\i[2518]  | ~\i[2516] );
  assign new_n4017_ = ~\i[755]  & ~\i[753]  & ~\i[754] ;
  assign new_n4018_ = ~\i[1195]  & ~\i[1194]  & ~\i[1192]  & ~\i[1193] ;
  assign new_n4019_ = ~\i[839]  & ~\i[838]  & ~\i[836]  & ~\i[837] ;
  assign new_n4020_ = ~\i[1867]  & ~\i[1866]  & ~\i[1864]  & ~\i[1865] ;
  assign new_n4021_ = \i[1411]  & \i[1409]  & \i[1410] ;
  assign new_n4022_ = ~new_n4020_ & (~new_n3546_ | ((new_n3415_ | ~new_n3349_) & (~\i[394]  | ~\i[395]  | new_n3349_)));
  assign new_n4023_ = (new_n4024_ | new_n4025_) & (~\i[524]  | ~\i[525]  | ~\i[526]  | ~\i[527]  | ~new_n4025_);
  assign new_n4024_ = \i[819]  & \i[818]  & \i[816]  & \i[817] ;
  assign new_n4025_ = ~\i[587]  & (~\i[586]  | (~\i[585]  & ~\i[584] ));
  assign new_n4026_ = \i[1531]  ? ((~new_n4027_ | new_n4048_) & (new_n4045_ | ~new_n4050_ | ~new_n4048_)) : new_n4032_;
  assign new_n4027_ = (~new_n4028_ | new_n4031_) & (\i[651]  | ~new_n4030_ | ~new_n4031_);
  assign new_n4028_ = new_n4029_ & ~\i[1060]  & ~\i[1061] ;
  assign new_n4029_ = ~\i[1062]  & ~\i[1063] ;
  assign new_n4030_ = ~\i[506]  & ~\i[507]  & (~\i[505]  | ~\i[504] );
  assign new_n4031_ = ~\i[766]  & ~\i[767] ;
  assign new_n4032_ = (new_n4038_ | new_n4042_ | new_n4044_) & (new_n4033_ | new_n4037_ | ~new_n4044_);
  assign new_n4033_ = ~new_n4036_ & ((~new_n4035_ & ~new_n4034_) | (\i[851]  & new_n4034_ & (\i[850]  | \i[849] )));
  assign new_n4034_ = ~\i[2423]  & (~\i[2422]  | (~\i[2421]  & ~\i[2420] ));
  assign new_n4035_ = ~\i[2175]  & ~\i[2173]  & ~\i[2174] ;
  assign new_n4036_ = ~\i[831]  & ~\i[829]  & ~\i[830] ;
  assign new_n4037_ = new_n4036_ & new_n3428_ & new_n4017_;
  assign new_n4038_ = ~new_n4040_ & (~new_n4041_ | ~new_n4039_) & (~\i[597]  | ~\i[598]  | ~\i[599]  | new_n4039_);
  assign new_n4039_ = \i[1067]  & \i[1065]  & \i[1066] ;
  assign new_n4040_ = \i[2311]  & \i[2310]  & \i[2308]  & \i[2309] ;
  assign new_n4041_ = \i[2630]  & \i[2631]  & (\i[2629]  | \i[2628] );
  assign new_n4042_ = ~new_n4043_ & ~\i[2439]  & new_n4040_ & (~\i[2438]  | ~\i[2437] );
  assign new_n4043_ = \i[2079]  & (\i[2078]  | (\i[2077]  & \i[2076] ));
  assign new_n4044_ = ~\i[1975]  & (~\i[1974]  | ~\i[1973] );
  assign new_n4045_ = new_n3666_ ? ~new_n4046_ : ~new_n4047_;
  assign new_n4046_ = \i[2067]  & \i[2066]  & \i[2064]  & \i[2065] ;
  assign new_n4047_ = \i[1315]  & (\i[1313]  | \i[1314]  | \i[1312] );
  assign new_n4048_ = \i[1081]  & new_n4049_ & \i[1080] ;
  assign new_n4049_ = \i[1082]  & \i[1083] ;
  assign new_n4050_ = ~\i[727]  & ~\i[725]  & ~\i[726] ;
  assign new_n4051_ = new_n4052_ ? (~new_n4081_ ^ new_n4095_) : (new_n4081_ ^ new_n4095_);
  assign new_n4052_ = new_n4007_ ? ((new_n4064_ | ~new_n3221_) & (new_n4073_ | new_n4076_ | new_n3221_)) : new_n4053_;
  assign new_n4053_ = new_n4058_ ? ((~new_n4059_ | ~new_n4061_) & (new_n4063_ | ~new_n4062_ | new_n4061_)) : new_n4054_;
  assign new_n4054_ = (~new_n4019_ | ~new_n4055_) & (~new_n4056_ | ~new_n3646_ | ~\i[1396]  | ~\i[1397]  | new_n4055_);
  assign new_n4055_ = new_n3869_ & (\i[1405]  | \i[1404] );
  assign new_n4056_ = new_n4057_ & ~\i[1388]  & ~\i[1389] ;
  assign new_n4057_ = ~\i[1390]  & ~\i[1391] ;
  assign new_n4058_ = \i[1405]  & new_n3869_ & \i[1404] ;
  assign new_n4059_ = ~new_n4060_ & ~\i[1734]  & ~\i[1735]  & (~\i[1733]  | ~\i[1732] );
  assign new_n4060_ = ~\i[2195]  & ~\i[2194]  & ~\i[2192]  & ~\i[2193] ;
  assign new_n4061_ = ~\i[835]  & ~\i[834]  & ~\i[832]  & ~\i[833] ;
  assign new_n4062_ = ~\i[1303]  & ~\i[1302]  & ~\i[1300]  & ~\i[1301] ;
  assign new_n4063_ = ~\i[507]  & ~\i[506]  & ~\i[504]  & ~\i[505] ;
  assign new_n4064_ = (new_n4070_ | ~new_n4071_ | new_n4069_) & (~new_n4069_ | (new_n4072_ ? ~new_n4067_ : ~new_n4065_));
  assign new_n4065_ = \i[1849]  & new_n4066_ & \i[1848] ;
  assign new_n4066_ = \i[1850]  & \i[1851] ;
  assign new_n4067_ = new_n4068_ & ~\i[1200]  & ~\i[1201] ;
  assign new_n4068_ = ~\i[1202]  & ~\i[1203] ;
  assign new_n4069_ = ~\i[2203]  & ~\i[2202]  & ~\i[2200]  & ~\i[2201] ;
  assign new_n4070_ = \i[1967]  & \i[1966]  & \i[1964]  & \i[1965] ;
  assign new_n4071_ = \i[2075]  & \i[2074]  & \i[2072]  & \i[2073] ;
  assign new_n4072_ = ~\i[1863]  & ~\i[1861]  & ~\i[1862] ;
  assign new_n4073_ = (~new_n4062_ | ~new_n4074_) & (~\i[1959]  | ((~\i[1958]  | new_n4074_) & (~\i[1957]  | (new_n4074_ & (~\i[1956]  | ~\i[1958] )))));
  assign new_n4074_ = new_n3708_ & new_n4075_;
  assign new_n4075_ = \i[1962]  & \i[1963] ;
  assign new_n4076_ = new_n4077_ & ((~new_n4079_ & ~new_n4080_) | (~\i[2090]  & ~\i[2091]  & new_n4080_));
  assign new_n4077_ = \i[1957]  & new_n4078_ & \i[1956] ;
  assign new_n4078_ = \i[1958]  & \i[1959] ;
  assign new_n4079_ = \i[1178]  & \i[1179]  & (\i[1177]  | \i[1176] );
  assign new_n4080_ = ~\i[1499]  & ~\i[1498]  & ~\i[1496]  & ~\i[1497] ;
  assign new_n4081_ = (new_n4082_ | ~new_n3351_) & (~new_n4092_ | (~new_n4065_ & new_n4093_ & new_n4094_));
  assign new_n4082_ = (new_n4085_ | new_n4083_ | ~new_n4087_) & (new_n4088_ | new_n4087_ | (new_n4091_ & ~new_n4090_));
  assign new_n4083_ = new_n3288_ & new_n4084_ & \i[2515]  & (\i[2514]  | \i[2513] );
  assign new_n4084_ = ~\i[2735]  & ~\i[2734]  & ~\i[2732]  & ~\i[2733] ;
  assign new_n4085_ = new_n4086_ & ~new_n4019_ & ~new_n4084_;
  assign new_n4086_ = \i[1179]  & \i[1178]  & \i[1176]  & \i[1177] ;
  assign new_n4087_ = new_n3615_ & ~\i[1156]  & ~\i[1157] ;
  assign new_n4088_ = ~new_n4089_ & new_n4090_ & (\i[2119]  | (\i[2117]  & \i[2118] ));
  assign new_n4089_ = \i[391]  & (\i[389]  | \i[390]  | \i[388] );
  assign new_n4090_ = ~\i[402]  & ~\i[403]  & (~\i[401]  | ~\i[400] );
  assign new_n4091_ = ~\i[719]  & ~\i[718]  & ~\i[716]  & ~\i[717] ;
  assign new_n4092_ = ~new_n3351_ & (~\i[278]  | ~\i[279] ) & (~new_n4008_ | new_n4093_);
  assign new_n4093_ = \i[1511]  & \i[1510]  & \i[1508]  & \i[1509] ;
  assign new_n4094_ = ~\i[1519]  & ~\i[1517]  & ~\i[1518] ;
  assign new_n4095_ = ~new_n4101_ & (~new_n3257_ | (~new_n4096_ & (~new_n4104_ | ~new_n4100_ | ~new_n4105_)));
  assign new_n4096_ = new_n4097_ & new_n4099_ & ~new_n4098_ & ~new_n4100_;
  assign new_n4097_ = \i[1513]  & new_n3560_ & \i[1512] ;
  assign new_n4098_ = \i[398]  & \i[399] ;
  assign new_n4099_ = \i[1175]  & \i[1174]  & \i[1172]  & \i[1173] ;
  assign new_n4100_ = ~\i[1051]  & ~\i[1050]  & ~\i[1048]  & ~\i[1049] ;
  assign new_n4101_ = ~new_n3677_ & ~new_n3257_ & new_n4103_ & (new_n4102_ | (new_n4007_ & new_n4080_));
  assign new_n4102_ = \i[427]  & \i[426]  & ~new_n4080_ & \i[425] ;
  assign new_n4103_ = new_n3798_ & (~\i[1861]  | ~\i[1860] );
  assign new_n4104_ = (new_n3669_ | ~new_n4020_) & (\i[274]  | \i[275]  | new_n4020_ | (\i[273]  & \i[272] ));
  assign new_n4105_ = ~\i[711]  & ~\i[710]  & ~\i[708]  & ~\i[709] ;
  assign new_n4106_ = ~new_n4110_ & ((new_n4107_ & new_n4111_ & new_n4112_) | (new_n4108_ & new_n4113_ & ~new_n4112_));
  assign new_n4107_ = ~new_n3383_ & \i[1287]  & (\i[1286]  | \i[1285]  | \i[1284] );
  assign new_n4108_ = new_n4109_ & (\i[515]  | (\i[513]  & \i[514] ));
  assign new_n4109_ = ~\i[1842]  & ~\i[1843] ;
  assign new_n4110_ = ~\i[2519]  & ~\i[2517]  & ~\i[2518] ;
  assign new_n4111_ = ~\i[2395]  & ~\i[2394]  & ~\i[2392]  & ~\i[2393] ;
  assign new_n4112_ = \i[1179]  & (\i[1177]  | \i[1178]  | \i[1176] );
  assign new_n4113_ = ~\i[1399]  & ~\i[1398]  & ~\i[1396]  & ~\i[1397] ;
  assign new_n4114_ = new_n4115_ ? (~new_n4106_ ^ new_n4169_) : (new_n4106_ ^ new_n4169_);
  assign new_n4115_ = new_n4116_ ? (new_n4137_ ^ new_n4155_) : (~new_n4137_ ^ new_n4155_);
  assign new_n4116_ = new_n3873_ ? ((~new_n4117_ & ~new_n4135_) | (new_n4133_ & new_n4136_ & new_n4135_)) : new_n4123_;
  assign new_n4117_ = ~new_n4118_ & (~new_n4122_ | (\i[2636]  & \i[2637]  & \i[2638]  & \i[2639] ));
  assign new_n4118_ = new_n4121_ & new_n4119_ & new_n3603_;
  assign new_n4119_ = new_n4120_ & ~\i[824]  & ~\i[825] ;
  assign new_n4120_ = ~\i[826]  & ~\i[827] ;
  assign new_n4121_ = \i[2179]  & \i[2178]  & \i[2176]  & \i[2177] ;
  assign new_n4122_ = ~new_n3603_ & (~\i[2735]  | (~\i[2733]  & ~\i[2734] ));
  assign new_n4123_ = new_n4131_ ? new_n4127_ : ((~new_n4124_ & new_n3770_) | (~new_n4132_ & \i[2743]  & ~new_n3770_));
  assign new_n4124_ = ~new_n4125_ & (~new_n4126_ | ~new_n3228_);
  assign new_n4125_ = ~new_n4126_ & (~\i[1523]  | (~\i[1522]  & (~\i[1521]  | ~\i[1520] )));
  assign new_n4126_ = \i[751]  & (\i[749]  | \i[750]  | \i[748] );
  assign new_n4127_ = ~new_n4128_ & (~\i[1727]  | (~\i[1725]  & ~\i[1726] ));
  assign new_n4128_ = new_n4129_ ? ~new_n4130_ : (~\i[2303]  & (~\i[2300]  | ~\i[2301]  | ~\i[2302] ));
  assign new_n4129_ = ~\i[1519]  & (~\i[1518]  | (~\i[1517]  & ~\i[1516] ));
  assign new_n4130_ = \i[2415]  & \i[2414]  & \i[2412]  & \i[2413] ;
  assign new_n4131_ = new_n3549_ & (~\i[1509]  | ~\i[1508] );
  assign new_n4132_ = ~\i[723]  & ~\i[722]  & ~\i[720]  & ~\i[721] ;
  assign new_n4133_ = \i[2307]  & new_n4134_ & \i[2306] ;
  assign new_n4134_ = new_n3670_ & ~\i[1940]  & ~\i[1941] ;
  assign new_n4135_ = \i[2535]  & (\i[2534]  | (\i[2533]  & \i[2532] ));
  assign new_n4136_ = \i[1174]  & \i[1175]  & (\i[1173]  | \i[1172] );
  assign new_n4137_ = ~new_n4144_ & (new_n4151_ | ~new_n4138_);
  assign new_n4138_ = new_n4143_ & (new_n4139_ | ~\i[2314]  | ~\i[2315] );
  assign new_n4139_ = ~new_n4140_ & (~new_n3555_ | ~new_n4142_ | ~\i[1734]  | ~\i[1735] );
  assign new_n4140_ = ~new_n4142_ & ~\i[1955]  & new_n4141_ & (~\i[1954]  | ~\i[1953]  | ~\i[1952] );
  assign new_n4141_ = ~\i[2646]  & ~\i[2647]  & (~\i[2645]  | ~\i[2644] );
  assign new_n4142_ = ~\i[1855]  & (~\i[1854]  | ~\i[1853] );
  assign new_n4143_ = ~\i[1863]  & (~\i[1862]  | ~\i[1861] );
  assign new_n4144_ = ~new_n4143_ & (new_n4146_ | (new_n4145_ & (~new_n4150_ | ~new_n4149_)));
  assign new_n4145_ = ~new_n3517_ & ~\i[699]  & (~\i[698]  | (~\i[696]  & ~\i[697] ));
  assign new_n4146_ = new_n3517_ & (~new_n3451_ | ~new_n4147_ | ~new_n4148_);
  assign new_n4147_ = \i[1295]  & \i[1293]  & \i[1294] ;
  assign new_n4148_ = ~\i[1867]  & (~\i[1866]  | ~\i[1865] );
  assign new_n4149_ = \i[627]  & \i[625]  & \i[626] ;
  assign new_n4150_ = \i[2627]  & \i[2625]  & \i[2626] ;
  assign new_n4151_ = (~\i[2314]  | ~\i[2315] ) & ((new_n4152_ & new_n4154_) | (~\i[1171]  & new_n4120_ & ~new_n4154_));
  assign new_n4152_ = new_n4013_ & \i[2431]  & (\i[2430]  | new_n4153_);
  assign new_n4153_ = \i[2428]  & \i[2429] ;
  assign new_n4154_ = ~\i[711]  & (~\i[710]  | (~\i[709]  & ~\i[708] ));
  assign new_n4155_ = (~\i[2338]  & ~\i[2339] ) ? (new_n4156_ | new_n4163_) : new_n4168_;
  assign new_n4156_ = new_n4157_ & ((~new_n4159_ & \i[743] ) | (~new_n3897_ & new_n4162_ & ~\i[743] ));
  assign new_n4157_ = new_n4158_ & (~\i[1265]  | ~\i[1264] );
  assign new_n4158_ = ~\i[1266]  & ~\i[1267] ;
  assign new_n4159_ = (~new_n4161_ | new_n4160_) & (\i[506]  | \i[507]  | ~new_n4160_);
  assign new_n4160_ = \i[1075]  & (\i[1074]  | (\i[1073]  & \i[1072] ));
  assign new_n4161_ = \i[599]  & (\i[598]  | (\i[597]  & \i[596] ));
  assign new_n4162_ = ~\i[1191]  & ~\i[1190]  & ~\i[1188]  & ~\i[1189] ;
  assign new_n4163_ = ~new_n4157_ & (new_n4165_ ? new_n4167_ : (new_n4166_ | new_n4164_));
  assign new_n4164_ = \i[499]  & \i[497]  & \i[498] ;
  assign new_n4165_ = \i[2287]  & \i[2285]  & \i[2286] ;
  assign new_n4166_ = \i[510]  & \i[511] ;
  assign new_n4167_ = ~\i[1490]  & ~\i[1491] ;
  assign new_n4168_ = ~\i[1735]  & (~\i[1734]  | (~\i[1733]  & ~\i[1732] ));
  assign new_n4169_ = (new_n4180_ | ~new_n4181_) & (new_n4173_ | new_n4181_ | (new_n4013_ & (new_n4178_ | new_n4170_)));
  assign new_n4170_ = new_n4132_ & ~new_n4171_ & ~new_n4172_;
  assign new_n4171_ = \i[1071]  & (\i[1070]  | new_n3667_);
  assign new_n4172_ = ~\i[739]  & (~\i[737]  | ~\i[738]  | ~\i[736] );
  assign new_n4173_ = ~new_n4013_ & (new_n4174_ | new_n4177_) & (~\i[2537]  | ~\i[2538]  | ~\i[2539]  | ~new_n4177_);
  assign new_n4174_ = new_n4175_ ? ~new_n4176_ : (~\i[2515]  | (~\i[2514]  & new_n3776_));
  assign new_n4175_ = ~\i[1078]  & ~\i[1079]  & (~\i[1077]  | ~\i[1076] );
  assign new_n4176_ = \i[2295]  & (\i[2294]  | \i[2293] );
  assign new_n4177_ = ~\i[2415]  & (~\i[2414]  | ~\i[2413] );
  assign new_n4178_ = ~new_n4132_ & (new_n3422_ ? (\i[739]  | (\i[737]  & \i[738] )) : new_n4179_);
  assign new_n4179_ = ~\i[519]  & ~\i[517]  & ~\i[518] ;
  assign new_n4180_ = ~\i[763]  & (~\i[762]  | (~\i[761]  & ~\i[760] ));
  assign new_n4181_ = \i[1090]  & \i[1091]  & (\i[1089]  | \i[1088] );
  assign new_n4182_ = ~new_n4183_ & (~new_n4197_ | (new_n4196_ & (~new_n4199_ | (\i[2060]  & \i[2061] ))));
  assign new_n4183_ = new_n4195_ & (new_n4184_ | (new_n4191_ & (new_n4190_ | new_n4194_ | ~new_n4192_)));
  assign new_n4184_ = ~new_n4187_ & (new_n4188_ ? ~new_n4185_ : (new_n3524_ ? new_n3745_ : new_n4189_));
  assign new_n4185_ = (~new_n4186_ | ~new_n3273_) & (\i[600]  | \i[601]  | \i[602]  | \i[603]  | new_n3273_);
  assign new_n4186_ = \i[1739]  & \i[1737]  & \i[1738] ;
  assign new_n4187_ = \i[1078]  & \i[1079]  & (\i[1077]  | \i[1076] );
  assign new_n4188_ = ~\i[747]  & (~\i[746]  | ~\i[745] );
  assign new_n4189_ = ~\i[1067]  & ~\i[1065]  & ~\i[1066] ;
  assign new_n4190_ = new_n3384_ & ~\i[1524]  & ~\i[1525] ;
  assign new_n4191_ = new_n4187_ & (new_n4192_ | new_n4193_ | ~\i[1963]  | (~\i[1962]  & ~new_n3708_));
  assign new_n4192_ = \i[1631]  & \i[1630]  & \i[1628]  & \i[1629] ;
  assign new_n4193_ = \i[2627]  & \i[2626]  & \i[2624]  & \i[2625] ;
  assign new_n4194_ = \i[1411]  & \i[1410]  & \i[1408]  & \i[1409] ;
  assign new_n4195_ = ~\i[1054]  & ~\i[1055]  & (~\i[1053]  | ~\i[1052] );
  assign new_n4196_ = (\i[2425]  | \i[2426]  | \i[2427] ) & (~new_n3658_ | ~\i[614]  | ~\i[615] );
  assign new_n4197_ = ~new_n4195_ & (~new_n4198_ | (\i[724]  & \i[725]  & \i[726]  & \i[727] ));
  assign new_n4198_ = ~\i[2426]  & ~\i[2427]  & ~\i[719]  & ~\i[2425]  & (~\i[2859]  | ~\i[2858] );
  assign new_n4199_ = ~\i[2062]  & ~\i[2063] ;
  assign new_n4200_ = new_n4201_ ? (new_n4295_ ^ new_n4311_) : (~new_n4295_ ^ new_n4311_);
  assign new_n4201_ = new_n4202_ ? (new_n4252_ ^ new_n4280_) : (~new_n4252_ ^ new_n4280_);
  assign new_n4202_ = new_n4203_ ? (new_n4227_ ^ new_n4242_) : (~new_n4227_ ^ new_n4242_);
  assign new_n4203_ = new_n4226_ ? new_n4204_ : ((new_n4212_ | ~new_n4220_) & (new_n4221_ | new_n4224_ | new_n4220_));
  assign new_n4204_ = \i[2523]  ? ((new_n4208_ & ~new_n4210_) | (~new_n4211_ & new_n4060_ & new_n4210_)) : new_n4205_;
  assign new_n4205_ = (\i[1402]  & \i[1403] ) ? new_n4207_ : ~new_n4206_;
  assign new_n4206_ = new_n4109_ & ~\i[1840]  & ~\i[1841] ;
  assign new_n4207_ = ~\i[2207]  & ~\i[2205]  & ~\i[2206] ;
  assign new_n4208_ = ~new_n4209_ & \i[2171]  & (\i[2170]  | \i[2169] );
  assign new_n4209_ = ~\i[2418]  & ~\i[2419]  & (~\i[2417]  | ~\i[2416] );
  assign new_n4210_ = \i[2747]  & (\i[2746]  | (\i[2745]  & \i[2744] ));
  assign new_n4211_ = \i[2855]  & \i[2854]  & \i[2852]  & \i[2853] ;
  assign new_n4212_ = (new_n4213_ | new_n4218_) & (~new_n4217_ | ~new_n4219_ | ~new_n4218_);
  assign new_n4213_ = (~new_n4216_ | ~new_n4214_) & (~\i[627]  | new_n4214_ | (~\i[626]  & (~\i[624]  | ~\i[625] )));
  assign new_n4214_ = new_n4215_ & ~\i[840]  & ~\i[841] ;
  assign new_n4215_ = ~\i[842]  & ~\i[843] ;
  assign new_n4216_ = ~\i[619]  & ~\i[618]  & ~\i[616]  & ~\i[617] ;
  assign new_n4217_ = new_n3269_ & (~\i[1609]  | ~\i[1608] );
  assign new_n4218_ = \i[1955]  & (\i[1954]  | (\i[1953]  & \i[1952] ));
  assign new_n4219_ = ~\i[2083]  & ~\i[2081]  & ~\i[2082] ;
  assign new_n4220_ = new_n3638_ & ~\i[2296]  & ~\i[2297] ;
  assign new_n4221_ = ~new_n4222_ & (~new_n4223_ | (~\i[823]  & \i[822]  & (\i[821]  | \i[820] )));
  assign new_n4222_ = \i[1187]  & (\i[1185]  | \i[1186]  | \i[1184] );
  assign new_n4223_ = ~\i[823]  & ~\i[1307]  & (~\i[1306]  | (~\i[1304]  & ~\i[1305] ));
  assign new_n4224_ = new_n4222_ & (~new_n4225_ | ~\i[624]  | ~\i[625]  | ~\i[626]  | ~\i[627] );
  assign new_n4225_ = \i[2294]  & \i[2295]  & (\i[2293]  | \i[2292] );
  assign new_n4226_ = \i[2299]  & \i[2298]  & \i[2296]  & \i[2297] ;
  assign new_n4227_ = new_n4241_ ? ((~new_n4239_ & ~\i[2427]  & new_n4240_) | (~new_n3543_ & ~new_n4240_)) : new_n4228_;
  assign new_n4228_ = (new_n4229_ | new_n4238_) & (new_n4233_ | new_n4237_ | ~new_n4238_);
  assign new_n4229_ = new_n3646_ ? (~new_n4232_ & (\i[945]  | \i[946]  | \i[947] )) : new_n4230_;
  assign new_n4230_ = (~new_n4029_ | ~new_n4231_) & (\i[1626]  | \i[1627]  | new_n4231_ | (\i[1625]  & \i[1624] ));
  assign new_n4231_ = \i[2063]  & (\i[2061]  | \i[2062]  | \i[2060] );
  assign new_n4232_ = ~\i[2750]  & ~\i[2751]  & (~\i[2749]  | ~\i[2748] );
  assign new_n4233_ = new_n4235_ & (new_n4234_ ? ~new_n4236_ : ~new_n3520_);
  assign new_n4234_ = ~\i[615]  & (~\i[614]  | (~\i[613]  & ~\i[612] ));
  assign new_n4235_ = ~\i[1286]  & ~\i[1287] ;
  assign new_n4236_ = ~\i[1835]  & ~\i[1833]  & ~\i[1834] ;
  assign new_n4237_ = ~new_n4235_ & ~\i[1502]  & ~\i[1503]  & (\i[1299]  | \i[1298]  | \i[1297] );
  assign new_n4238_ = ~\i[1618]  & ~\i[1619]  & (~\i[1617]  | ~\i[1616] );
  assign new_n4239_ = \i[1735]  & \i[1734]  & \i[1732]  & \i[1733] ;
  assign new_n4240_ = \i[2195]  & (\i[2194]  | \i[2193] );
  assign new_n4241_ = \i[1751]  & (\i[1749]  | \i[1750]  | \i[1748] );
  assign new_n4242_ = new_n4250_ ? (~new_n3669_ | (~new_n4243_ & ~new_n4248_)) : ~new_n4251_;
  assign new_n4243_ = new_n4246_ & (new_n4028_ ? new_n4247_ : new_n4244_);
  assign new_n4244_ = \i[1061]  & new_n4245_ & \i[1060] ;
  assign new_n4245_ = \i[1062]  & \i[1063] ;
  assign new_n4246_ = ~\i[735]  & (~\i[734]  | (~\i[733]  & ~\i[732] ));
  assign new_n4247_ = \i[1627]  & (\i[1625]  | \i[1626]  | \i[1624] );
  assign new_n4248_ = ~new_n4246_ & (new_n3442_ ? ~new_n3741_ : new_n4249_);
  assign new_n4249_ = ~\i[1739]  & (~\i[1738]  | ~\i[1737] );
  assign new_n4250_ = ~\i[2223]  & (~\i[2222]  | (~\i[2221]  & ~\i[2220] ));
  assign new_n4251_ = \i[2159]  & \i[2158]  & \i[2156]  & \i[2157] ;
  assign new_n4252_ = new_n4253_ ? (new_n4260_ ^ new_n4270_) : (~new_n4260_ ^ new_n4270_);
  assign new_n4253_ = new_n4044_ ? (~new_n4254_ & (new_n3597_ | new_n4257_ | \i[2311] )) : new_n4258_;
  assign new_n4254_ = new_n4257_ & (new_n3564_ ? new_n4255_ : (\i[1963]  | \i[1962] ));
  assign new_n4255_ = (~\i[838]  & ~\i[839] ) ? new_n3467_ : ~new_n4256_;
  assign new_n4256_ = \i[627]  & (\i[625]  | \i[626]  | \i[624] );
  assign new_n4257_ = ~\i[1403]  & ~\i[1402]  & ~\i[1400]  & ~\i[1401] ;
  assign new_n4258_ = ~new_n4259_ & \i[2082]  & \i[2083]  & (\i[2081]  | \i[2080] );
  assign new_n4259_ = ~new_n3431_ & ~\i[2537]  & ~\i[2538]  & ~\i[2539]  & (~\i[839]  | ~\i[838] );
  assign new_n4260_ = new_n4157_ ? ((new_n4261_ | new_n4269_ | ~new_n3373_) & (new_n4263_ | new_n3373_)) : ~new_n4267_;
  assign new_n4261_ = new_n3290_ & (~\i[1632]  | ~\i[1633] ) & (new_n3301_ ? ~new_n3545_ : new_n4262_);
  assign new_n4262_ = \i[747]  & (\i[745]  | \i[746]  | \i[744] );
  assign new_n4263_ = ~new_n4264_ & ((new_n4214_ & (\i[2490]  | \i[2491] )) | ~\i[1415]  | (new_n4265_ & ~\i[2490]  & ~\i[2491] ));
  assign new_n4264_ = ~new_n4175_ & ~\i[1415]  & (\i[2224]  | \i[2225]  | \i[2226]  | \i[2227] );
  assign new_n4265_ = \i[2521]  & new_n4266_ & \i[2520] ;
  assign new_n4266_ = \i[2522]  & \i[2523] ;
  assign new_n4267_ = ~\i[506]  & ~\i[507]  & ~\i[505]  & new_n4268_ & (~\i[2325]  | ~\i[2324] );
  assign new_n4268_ = ~\i[2326]  & ~\i[2327] ;
  assign new_n4269_ = (new_n4036_ | (~\i[1082]  & ~\i[1083] )) & (~new_n3290_ | (\i[1632]  & \i[1633] ));
  assign new_n4270_ = (~new_n3546_ | new_n4278_) & (new_n4276_ | new_n4271_ | ~new_n4279_ | ~new_n4278_);
  assign new_n4271_ = new_n4275_ & (new_n4274_ ? new_n4272_ : ~new_n3719_);
  assign new_n4272_ = new_n4273_ & (\i[1501]  | \i[1500] );
  assign new_n4273_ = \i[1502]  & \i[1503] ;
  assign new_n4274_ = ~\i[2747]  & (~\i[2746]  | (~\i[2745]  & ~\i[2744] ));
  assign new_n4275_ = ~\i[1495]  & ~\i[1494]  & ~\i[1492]  & ~\i[1493] ;
  assign new_n4276_ = ~new_n4275_ & (\i[1410]  | \i[1411] ) & (~new_n4277_ | (\i[1728]  & \i[1729] ));
  assign new_n4277_ = ~\i[1730]  & ~\i[1731] ;
  assign new_n4278_ = ~\i[1491]  & (~\i[1490]  | (~\i[1489]  & ~\i[1488] ));
  assign new_n4279_ = ~\i[2847]  & (~\i[2846]  | (~\i[2845]  & ~\i[2844] ));
  assign new_n4280_ = (new_n4290_ | ~new_n4281_) & (new_n4283_ | (~new_n4284_ & (~new_n4292_ | ~new_n4294_)));
  assign new_n4281_ = new_n4283_ & (~new_n4048_ | new_n4282_);
  assign new_n4282_ = (~new_n4097_ | ~new_n4017_) & (\i[730]  | \i[731]  | new_n4017_ | (\i[729]  & \i[728] ));
  assign new_n4283_ = \i[1419]  & (\i[1418]  | (\i[1417]  & \i[1416] ));
  assign new_n4284_ = ~new_n4287_ & (~new_n4288_ | (~new_n4285_ & ~new_n4289_));
  assign new_n4285_ = new_n4286_ & ~\i[2520]  & ~\i[2521] ;
  assign new_n4286_ = ~\i[2522]  & ~\i[2523] ;
  assign new_n4287_ = ~\i[707]  & ~\i[705]  & ~\i[706] ;
  assign new_n4288_ = ~\i[1067]  & ~\i[1066]  & ~\i[1064]  & ~\i[1065] ;
  assign new_n4289_ = \i[846]  & \i[847] ;
  assign new_n4290_ = ~new_n4048_ & \i[2171]  & ((new_n4291_ & \i[2170] ) | (\i[2168]  & \i[2169]  & ~\i[2170] ));
  assign new_n4291_ = \i[1083]  & (\i[1081]  | \i[1082]  | \i[1080] );
  assign new_n4292_ = ~new_n3669_ & ~new_n4293_;
  assign new_n4293_ = \i[1415]  & (\i[1413]  | \i[1414]  | \i[1412] );
  assign new_n4294_ = new_n4287_ & ((~\i[2001]  & ~\i[2000] ) | ~\i[2003]  | ~\i[2002] );
  assign new_n4295_ = new_n4110_ ? (new_n4305_ | (~new_n4272_ & ~new_n4307_)) : new_n4296_;
  assign new_n4296_ = new_n4112_ ? new_n4297_ : ((~new_n4302_ & new_n4113_) | (~new_n3238_ & ~new_n4304_ & ~new_n4113_));
  assign new_n4297_ = new_n4111_ ? new_n4298_ : (new_n4300_ ? new_n4069_ : ~new_n4301_);
  assign new_n4298_ = (\i[1287]  & (\i[1284]  | \i[1285]  | \i[1286] )) ? ~new_n3383_ : ~new_n4299_;
  assign new_n4299_ = ~\i[1278]  & ~\i[1279] ;
  assign new_n4300_ = \i[2083]  & \i[2081]  & \i[2082] ;
  assign new_n4301_ = \i[2403]  & \i[2401]  & \i[2402] ;
  assign new_n4302_ = ~new_n4108_ & (new_n4303_ | new_n4109_);
  assign new_n4303_ = ~\i[2527]  & ~\i[2526]  & ~\i[2524]  & ~\i[2525] ;
  assign new_n4304_ = \i[2175]  & (\i[2174]  | (\i[2173]  & \i[2172] ));
  assign new_n4305_ = new_n4306_ & (~new_n3534_ | (~\i[2192]  & ~\i[2193] ));
  assign new_n4306_ = new_n4272_ & ((~\i[2269]  & ~\i[2268] ) | ~\i[2271]  | ~\i[2270] );
  assign new_n4307_ = (new_n4308_ | new_n4309_) & (~new_n4310_ | ~new_n4309_ | (\i[1951]  & (\i[1949]  | \i[1950] )));
  assign new_n4308_ = \i[2202]  & \i[2203]  & (\i[2201]  | \i[2200] );
  assign new_n4309_ = ~\i[931]  & ~\i[929]  & ~\i[930] ;
  assign new_n4310_ = \i[1639]  & (\i[1638]  | (\i[1637]  & \i[1636] ));
  assign new_n4311_ = new_n3987_ ? new_n4317_ : (new_n3557_ ? new_n4318_ : new_n4312_);
  assign new_n4312_ = \i[2187]  ? (new_n4314_ | (new_n4315_ & new_n4316_)) : new_n4313_;
  assign new_n4313_ = new_n3988_ & (\i[2063]  | (\i[2061]  & \i[2062] ));
  assign new_n4314_ = ~new_n4315_ & \i[535]  & (\i[534]  | \i[533] );
  assign new_n4315_ = ~\i[1639]  & (~\i[1638]  | ~\i[1637] );
  assign new_n4316_ = ~\i[1199]  & (~\i[1198]  | (~\i[1197]  & ~\i[1196] ));
  assign new_n4317_ = ~\i[1619]  & ~\i[1618]  & ~\i[1616]  & ~\i[1617] ;
  assign new_n4318_ = ~\i[1306]  & ~\i[1307]  & \i[1531]  & (\i[1530]  | \i[1529] );
  assign new_n4319_ = new_n4345_ ? (~new_n4332_ & (new_n4341_ | new_n4344_ | new_n4340_)) : new_n4320_;
  assign new_n4320_ = new_n4219_ ? new_n4321_ : ((~new_n4327_ & new_n4265_) | (~new_n4331_ & new_n3993_ & ~new_n4265_));
  assign new_n4321_ = new_n4325_ ? new_n4322_ : (new_n3741_ ? new_n4078_ : new_n4326_);
  assign new_n4322_ = new_n4324_ ? (\i[2535]  | (\i[2533]  & \i[2534] )) : new_n4323_;
  assign new_n4323_ = ~\i[1386]  & ~\i[1387] ;
  assign new_n4324_ = \i[1058]  & \i[1059]  & (\i[1057]  | \i[1056] );
  assign new_n4325_ = ~\i[607]  & ~\i[606]  & ~\i[604]  & ~\i[605] ;
  assign new_n4326_ = \i[1963]  & (\i[1962]  | \i[1961] );
  assign new_n4327_ = new_n4329_ ? ~new_n4328_ : ~new_n4330_;
  assign new_n4328_ = ~\i[2290]  & ~\i[2291]  & (~\i[2289]  | ~\i[2288] );
  assign new_n4329_ = \i[2187]  & \i[2186]  & \i[2184]  & \i[2185] ;
  assign new_n4330_ = \i[1498]  & \i[1499] ;
  assign new_n4331_ = ~\i[2203]  & ~\i[2201]  & ~\i[2202] ;
  assign new_n4332_ = new_n4340_ & ~new_n4333_ & ~new_n4339_;
  assign new_n4333_ = new_n4336_ ? new_n4334_ : new_n4338_;
  assign new_n4334_ = new_n4335_ & ~\i[704]  & ~\i[705] ;
  assign new_n4335_ = ~\i[706]  & ~\i[707] ;
  assign new_n4336_ = new_n4337_ & ~\i[2064]  & ~\i[2065] ;
  assign new_n4337_ = ~\i[2066]  & ~\i[2067] ;
  assign new_n4338_ = \i[1283]  & \i[1282]  & \i[1280]  & \i[1281] ;
  assign new_n4339_ = \i[2331]  & (\i[2329]  | \i[2330]  | \i[2328] );
  assign new_n4340_ = ~\i[1622]  & ~\i[1623]  & (~\i[1621]  | ~\i[1620] );
  assign new_n4341_ = ~new_n4111_ & ((~new_n4343_ & ~new_n4342_) | (\i[2071]  & new_n4342_ & (\i[2070]  | \i[2069] )));
  assign new_n4342_ = \i[842]  & \i[843] ;
  assign new_n4343_ = ~\i[1063]  & (~\i[1061]  | ~\i[1062]  | ~\i[1060] );
  assign new_n4344_ = ~\i[2743]  & new_n4111_ & new_n4066_ & (~\i[2742]  | ~\i[2741] );
  assign new_n4345_ = \i[2303]  & \i[2302]  & \i[2300]  & \i[2301] ;
  assign new_n4346_ = new_n4347_ ? (new_n4383_ ^ new_n4399_) : (~new_n4383_ ^ new_n4399_);
  assign new_n4347_ = new_n4280_ ? (new_n4348_ ^ new_n4374_) : (~new_n4348_ ^ new_n4374_);
  assign new_n4348_ = new_n4349_ ? (new_n4358_ ^ new_n4365_) : (~new_n4358_ ^ new_n4365_);
  assign new_n4349_ = new_n4157_ & ((\i[2302]  & \i[2303] ) ? ~new_n4354_ : ~new_n4350_);
  assign new_n4350_ = (new_n4351_ | (\i[2187]  & (\i[2185]  | \i[2186] ))) & (~new_n3703_ | ~new_n4353_ | ~\i[2187]  | (~\i[2185]  & ~\i[2186] ));
  assign new_n4351_ = (~\i[2414]  & ~\i[2415] ) ? ~new_n4132_ : ~new_n4352_;
  assign new_n4352_ = \i[1959]  & (\i[1958]  | (\i[1957]  & \i[1956] ));
  assign new_n4353_ = \i[1295]  & \i[1294]  & \i[1292]  & \i[1293] ;
  assign new_n4354_ = (~new_n4357_ & new_n4356_ & new_n4355_) | (~new_n4355_ & (~new_n3546_ | ~new_n3583_));
  assign new_n4355_ = new_n4199_ & ~\i[2060]  & ~\i[2061] ;
  assign new_n4356_ = ~\i[2187]  & (~\i[2186]  | (~\i[2185]  & ~\i[2184] ));
  assign new_n4357_ = \i[1283]  & (\i[1282]  | (\i[1281]  & \i[1280] ));
  assign new_n4358_ = new_n4279_ & ~new_n4359_ & new_n3396_;
  assign new_n4359_ = (new_n4360_ & \i[2502]  & \i[2503]  & (\i[2500]  | \i[2501] )) | (new_n4363_ & (~\i[2502]  | ~\i[2503]  | (~\i[2500]  & ~\i[2501] )));
  assign new_n4360_ = (~new_n4361_ | ~new_n4362_) & (~new_n3287_ | ~\i[2056]  | ~\i[2057]  | new_n4362_);
  assign new_n4361_ = ~\i[838]  & ~\i[839]  & (~\i[837]  | ~\i[836] );
  assign new_n4362_ = ~\i[1291]  & ~\i[1289]  & ~\i[1290] ;
  assign new_n4363_ = (~\i[2321]  | ~\i[2322]  | ~\i[2323]  | new_n4364_) & (~new_n4364_ | (~\i[1291]  & ~\i[1290] ));
  assign new_n4364_ = ~\i[819]  & ~\i[818]  & ~\i[816]  & ~\i[817] ;
  assign new_n4365_ = new_n3858_ & ((~new_n4366_ & new_n4371_) | (new_n4370_ & new_n4373_ & ~new_n4371_));
  assign new_n4366_ = (~new_n4367_ | new_n4369_) & (new_n3990_ | ~new_n3703_ | ~new_n4369_);
  assign new_n4367_ = new_n4368_ & (\i[2311]  | (\i[2309]  & \i[2310] ));
  assign new_n4368_ = ~\i[2067]  & ~\i[2065]  & ~\i[2066] ;
  assign new_n4369_ = ~\i[603]  & ~\i[601]  & ~\i[602] ;
  assign new_n4370_ = new_n4097_ & (~\i[1723]  | ~\i[1722] );
  assign new_n4371_ = new_n4372_ & ~\i[1748]  & ~\i[1749] ;
  assign new_n4372_ = ~\i[1750]  & ~\i[1751] ;
  assign new_n4373_ = \i[1855]  & \i[1854]  & \i[1852]  & \i[1853] ;
  assign new_n4374_ = (new_n3372_ | new_n4381_ | ~new_n4382_ | ~\i[2087] ) & (~new_n4380_ | new_n4375_ | \i[2087] );
  assign new_n4375_ = (~new_n4376_ & new_n4241_) | (~new_n4378_ & ~new_n4241_ & (\i[411]  | (\i[409]  & \i[410] )));
  assign new_n4376_ = new_n4377_ & \i[2627]  & (\i[2626]  | (\i[2624]  & \i[2625] ));
  assign new_n4377_ = \i[2403]  & \i[2402]  & \i[2400]  & \i[2401] ;
  assign new_n4378_ = new_n4379_ & (\i[1073]  | \i[1072] );
  assign new_n4379_ = \i[1074]  & \i[1075] ;
  assign new_n4380_ = ~\i[883]  & ~\i[882]  & ~\i[880]  & ~\i[881] ;
  assign new_n4381_ = \i[1839]  & (\i[1837]  | \i[1838]  | \i[1836] );
  assign new_n4382_ = \i[2079]  & (\i[2077]  | \i[2078]  | \i[2076] );
  assign new_n4383_ = new_n4157_ ? new_n4384_ : new_n4394_;
  assign new_n4384_ = new_n4393_ ? new_n4387_ : (new_n4385_ | (~new_n4132_ & new_n4392_ & new_n3735_));
  assign new_n4385_ = (~\i[1186]  | (~new_n4386_ & (~\i[1187]  | ~\i[1185]  | ~\i[1184] ))) & (~new_n4386_ | (~\i[1187]  & (~\i[1185]  | ~\i[1184] ))) & (~new_n3854_ | new_n4386_);
  assign new_n4386_ = ~\i[1511]  & ~\i[1509]  & ~\i[1510] ;
  assign new_n4387_ = (new_n4388_ | ~new_n4391_) & (~new_n3322_ | new_n4391_ | (\i[2623]  & (\i[2621]  | \i[2622] )));
  assign new_n4388_ = (\i[1068]  | \i[1069]  | \i[1070]  | \i[1071]  | ~new_n4390_) & (~new_n4389_ | new_n4390_);
  assign new_n4389_ = ~\i[2171]  & ~\i[2170]  & ~\i[2168]  & ~\i[2169] ;
  assign new_n4390_ = ~\i[623]  & (~\i[622]  | ~\i[621] );
  assign new_n4391_ = \i[1186]  & \i[1187] ;
  assign new_n4392_ = \i[1185]  & new_n4391_ & \i[1184] ;
  assign new_n4393_ = ~\i[855]  & ~\i[854]  & ~\i[852]  & ~\i[853] ;
  assign new_n4394_ = (new_n4395_ & (\i[396]  | \i[397]  | \i[398]  | \i[399] )) | (new_n4397_ & ~\i[396]  & ~\i[397]  & ~\i[398]  & ~\i[399] );
  assign new_n4395_ = \i[953]  & new_n4396_ & \i[952] ;
  assign new_n4396_ = \i[954]  & \i[955] ;
  assign new_n4397_ = ~new_n4398_ & ((~\i[2489]  & ~\i[2488] ) | ~\i[2491]  | ~\i[2490] );
  assign new_n4398_ = \i[502]  & \i[503] ;
  assign new_n4399_ = (~new_n4281_ | new_n4400_) & (new_n4403_ | new_n4283_ | (new_n4294_ & ~new_n4292_));
  assign new_n4400_ = ~new_n4048_ & ((~new_n4401_ & new_n4402_) | (new_n4058_ & new_n3581_ & ~new_n4402_));
  assign new_n4401_ = \i[2171]  & ~new_n4291_ & \i[2170] ;
  assign new_n4402_ = \i[2171]  & (\i[2170]  | (\i[2169]  & \i[2168] ));
  assign new_n4403_ = ~new_n4287_ & ((new_n4119_ & ~new_n4288_) | (~new_n4285_ & new_n4289_ & new_n4288_));
  assign new_n4404_ = (~new_n4405_ & ~new_n4020_) | (~new_n4415_ & new_n4020_ & (~new_n4084_ | ~new_n4410_));
  assign new_n4405_ = ~new_n4406_ & ~new_n4408_ & ~\i[279]  & (~\i[278]  | ~\i[277] );
  assign new_n4406_ = new_n3770_ & ((~\i[1871]  & new_n4192_) | (\i[2731]  & ~new_n4192_ & (\i[2728]  | ~new_n4407_)));
  assign new_n4407_ = ~\i[2729]  & ~\i[2730] ;
  assign new_n4408_ = ~new_n3770_ & new_n4409_ & (\i[1891]  | (\i[1889]  & \i[1890] ));
  assign new_n4409_ = ~\i[1302]  & ~\i[1303]  & (~\i[1301]  | ~\i[1300] );
  assign new_n4410_ = new_n4219_ ? new_n4411_ : (~new_n4206_ | (~\i[2422]  & ~\i[2423] ));
  assign new_n4411_ = new_n4412_ ? ~new_n4413_ : (~new_n4414_ | (~\i[732]  & ~\i[733] ));
  assign new_n4412_ = new_n4299_ & (~\i[1277]  | ~\i[1276] );
  assign new_n4413_ = ~\i[718]  & ~\i[719]  & (~\i[717]  | ~\i[716] );
  assign new_n4414_ = \i[734]  & \i[735] ;
  assign new_n4415_ = ~new_n4084_ & (new_n4132_ ? (new_n4417_ ? ~new_n4418_ : ~new_n4419_) : ~new_n4416_);
  assign new_n4416_ = \i[1743]  & new_n3281_ & \i[1742] ;
  assign new_n4417_ = ~\i[1058]  & ~\i[1059]  & (~\i[1057]  | ~\i[1056] );
  assign new_n4418_ = ~\i[2079]  & (~\i[2077]  | ~\i[2078]  | ~\i[2076] );
  assign new_n4419_ = \i[1603]  & (\i[1602]  | (\i[1601]  & \i[1600] ));
  assign new_n4420_ = (new_n4421_ | ~new_n4437_) & (new_n4432_ | new_n4437_ | (\i[1175]  & (new_n4436_ | new_n4429_)));
  assign new_n4421_ = new_n4428_ ? ~new_n4422_ : ((~new_n4427_ & new_n3781_) | (~\i[739]  & new_n4093_ & ~new_n3781_));
  assign new_n4422_ = new_n3394_ ? ((~new_n4426_ | new_n4272_) & (~\i[2306]  | ~\i[2307]  | ~new_n4272_)) : new_n4423_;
  assign new_n4423_ = (~new_n4424_ | ~new_n4425_) & (~\i[2524]  | ~\i[2525]  | ~\i[2526]  | ~\i[2527]  | new_n4425_);
  assign new_n4424_ = \i[1299]  & \i[1298]  & \i[1296]  & \i[1297] ;
  assign new_n4425_ = \i[2499]  & \i[2498]  & \i[2496]  & \i[2497] ;
  assign new_n4426_ = ~\i[927]  & (~\i[926]  | (~\i[925]  & ~\i[924] ));
  assign new_n4427_ = new_n3597_ & (~\i[623]  | (~\i[620]  & ~\i[621]  & ~\i[622] ));
  assign new_n4428_ = ~\i[2519]  & ~\i[2518]  & ~\i[2516]  & ~\i[2517] ;
  assign new_n4429_ = new_n4431_ & ~new_n4430_ & new_n4226_;
  assign new_n4430_ = new_n3683_ & (~\i[1613]  | ~\i[1612] );
  assign new_n4431_ = \i[2755]  & \i[2754]  & \i[2752]  & \i[2753] ;
  assign new_n4432_ = new_n4435_ & new_n4433_ & (\i[2390]  | (\i[2388]  & \i[2389] ));
  assign new_n4433_ = new_n4434_ & ~\i[1528]  & ~\i[1529] ;
  assign new_n4434_ = ~\i[1530]  & ~\i[1531] ;
  assign new_n4435_ = ~\i[1175]  & \i[2391]  & (\i[1963]  | (\i[1961]  & \i[1962] ));
  assign new_n4436_ = \i[755]  & \i[754]  & \i[753]  & \i[752]  & ~new_n4226_ & new_n4338_;
  assign new_n4437_ = new_n3265_ & ~\i[1268]  & ~\i[1269] ;
  assign new_n4438_ = (~new_n3351_ & (new_n4449_ ? ~new_n4439_ : new_n4450_)) | (~new_n4443_ & ~new_n4452_ & new_n3351_);
  assign new_n4439_ = (new_n4442_ | \i[539]  | (\i[1290]  & \i[1291] )) & (~\i[1290]  | ~\i[1291]  | new_n4440_ | new_n3628_);
  assign new_n4440_ = \i[1413]  & new_n4441_ & \i[1412] ;
  assign new_n4441_ = \i[1414]  & \i[1415] ;
  assign new_n4442_ = \i[415]  & (\i[414]  | (\i[413]  & \i[412] ));
  assign new_n4443_ = ~new_n4444_ & ~new_n4446_ & (new_n4445_ | (new_n4019_ & ~new_n4447_) | (new_n4448_ & new_n4447_));
  assign new_n4444_ = new_n4445_ & (~new_n4219_ | new_n3564_) & (\i[1081]  | \i[1082]  | \i[1083]  | ~new_n3564_);
  assign new_n4445_ = ~\i[1419]  & ~\i[1417]  & ~\i[1418] ;
  assign new_n4446_ = \i[1739]  & \i[1738]  & \i[1736]  & \i[1737] ;
  assign new_n4447_ = ~\i[2482]  & ~\i[2483]  & (~\i[2481]  | ~\i[2480] );
  assign new_n4448_ = \i[651]  & \i[649]  & \i[650] ;
  assign new_n4449_ = new_n3220_ & ~\i[1756]  & ~\i[1757] ;
  assign new_n4450_ = new_n4451_ & ((~\i[277]  & ~\i[276] ) | ~\i[279]  | ~\i[278] );
  assign new_n4451_ = ~\i[1675]  & ~\i[1674]  & ~\i[1672]  & ~\i[1673] ;
  assign new_n4452_ = new_n4446_ & ((~new_n4453_ & ~new_n4454_ & ~new_n3242_) | (~new_n3988_ & new_n3898_ & new_n3242_));
  assign new_n4453_ = ~\i[1410]  & ~\i[1411]  & (~\i[1409]  | ~\i[1408] );
  assign new_n4454_ = ~\i[407]  & ~\i[405]  & ~\i[406] ;
  assign new_n4455_ = new_n3257_ ? (new_n4470_ ? new_n4460_ : new_n4466_) : new_n4456_;
  assign new_n4456_ = (~new_n3990_ | ~new_n4275_ | ~new_n4459_) & (new_n4459_ | (new_n4046_ ? new_n4458_ : ~new_n4457_));
  assign new_n4457_ = \i[583]  & \i[582]  & \i[581]  & ~new_n4103_ & \i[580] ;
  assign new_n4458_ = (~new_n3592_ | ~new_n4424_) & (~\i[277]  | ~\i[278]  | ~\i[279]  | new_n4424_);
  assign new_n4459_ = \i[650]  & \i[651]  & (\i[649]  | \i[648] );
  assign new_n4460_ = (~new_n4463_ | (new_n4462_ ? new_n3775_ : ~new_n4461_)) & (~new_n4464_ | ~new_n4465_ | new_n4463_);
  assign new_n4461_ = ~\i[2083]  & ~\i[2082]  & ~\i[2080]  & ~\i[2081] ;
  assign new_n4462_ = \i[1739]  & (\i[1737]  | \i[1738]  | \i[1736] );
  assign new_n4463_ = ~\i[823]  & ~\i[822]  & ~\i[820]  & ~\i[821] ;
  assign new_n4464_ = ~\i[398]  & ~\i[399]  & (~\i[397]  | ~\i[396] );
  assign new_n4465_ = \i[1170]  & \i[1171]  & (\i[1169]  | \i[1168] );
  assign new_n4466_ = (~new_n4467_ | ~\i[487]  | new_n4468_) & (~new_n4192_ | ~new_n4469_ | ~new_n4468_);
  assign new_n4467_ = \i[1055]  & \i[1054]  & \i[1052]  & \i[1053] ;
  assign new_n4468_ = \i[1290]  & \i[1291]  & (\i[1289]  | \i[1288] );
  assign new_n4469_ = ~\i[395]  & ~\i[393]  & ~\i[394] ;
  assign new_n4470_ = new_n4471_ & ~\i[1272]  & ~\i[1273] ;
  assign new_n4471_ = ~\i[1274]  & ~\i[1275] ;
  assign \o[8]  = new_n4473_ ? (new_n4474_ ^ new_n4475_) : (~new_n4474_ ^ new_n4475_);
  assign new_n4473_ = ~new_n3975_ & ~new_n4455_;
  assign new_n4474_ = (~new_n4420_ & ~new_n4438_) | (new_n3976_ & (~new_n4420_ | ~new_n4438_));
  assign new_n4475_ = new_n4476_ ? (~new_n4477_ ^ new_n4568_) : (new_n4477_ ^ new_n4568_);
  assign new_n4476_ = (~new_n4404_ & new_n4346_) | (new_n3977_ & (~new_n4404_ | new_n4346_));
  assign new_n4477_ = new_n4478_ ? (new_n4479_ ^ new_n4559_) : (~new_n4479_ ^ new_n4559_);
  assign new_n4478_ = (~new_n4319_ & new_n4200_) | (new_n3978_ & (~new_n4319_ | new_n4200_));
  assign new_n4479_ = new_n4480_ ? (new_n4481_ ^ new_n4537_) : (~new_n4481_ ^ new_n4537_);
  assign new_n4480_ = (~new_n4182_ & new_n4114_) | (new_n3979_ & (~new_n4182_ | new_n4114_));
  assign new_n4481_ = new_n4482_ ? (new_n4496_ ^ new_n4497_) : (~new_n4496_ ^ new_n4497_);
  assign new_n4482_ = new_n4483_ ? (~new_n4484_ ^ new_n4485_) : (new_n4484_ ^ new_n4485_);
  assign new_n4483_ = (~new_n4026_ & new_n4003_) | (~new_n3981_ & (~new_n4026_ | new_n4003_));
  assign new_n4484_ = (~new_n4137_ & new_n4155_) | (~new_n4116_ & (~new_n4137_ | new_n4155_));
  assign new_n4485_ = new_n4486_ ? (~new_n4488_ ^ new_n4492_) : (new_n4488_ ^ new_n4492_);
  assign new_n4486_ = new_n4020_ ? ((new_n4410_ | ~new_n4084_) & (new_n4487_ | ~new_n4132_ | new_n4084_)) : new_n4405_;
  assign new_n4487_ = new_n4417_ ? ~new_n4418_ : ~new_n4419_;
  assign new_n4488_ = (new_n4489_ | \i[1531] ) & (~new_n3989_ | ~\i[2497]  | ~\i[2498]  | ~\i[2499]  | ~\i[1531] );
  assign new_n4489_ = ~new_n4490_ & (new_n3998_ | ((~new_n3999_ | ~new_n4002_) & (new_n4331_ | ~new_n4491_ | new_n4002_)));
  assign new_n4490_ = \i[1511]  & \i[1510]  & \i[1509]  & new_n3998_ & ~new_n3993_ & ~new_n3756_;
  assign new_n4491_ = ~\i[2087]  & ~\i[2086]  & ~\i[2084]  & ~\i[2085] ;
  assign new_n4492_ = (new_n4437_ & (new_n4428_ ? new_n4422_ : new_n4493_)) | (~new_n4495_ & ~new_n4432_ & ~new_n4437_);
  assign new_n4493_ = (new_n3300_ | ~new_n4494_ | ~\i[623]  | ~new_n3781_) & (~new_n4093_ | \i[739]  | new_n3781_);
  assign new_n4494_ = \i[959]  & \i[957]  & \i[958] ;
  assign new_n4495_ = \i[1175]  & (new_n4436_ | (new_n4226_ & (new_n4430_ ? new_n3592_ : new_n4431_)));
  assign new_n4496_ = (~new_n4051_ & new_n4106_) | (new_n3980_ & (~new_n4051_ | new_n4106_));
  assign new_n4497_ = new_n4498_ ? (new_n4514_ ^ new_n4515_) : (~new_n4514_ ^ new_n4515_);
  assign new_n4498_ = new_n4499_ ? (~new_n4503_ ^ new_n4507_) : (new_n4503_ ^ new_n4507_);
  assign new_n4499_ = (new_n4500_ | ~new_n3259_) & (~new_n4011_ | ~new_n4012_ | ~new_n4013_ | new_n3259_);
  assign new_n4500_ = new_n4020_ ? ((~new_n4502_ | ~new_n4018_) & (~new_n4019_ | ~new_n4021_ | new_n4018_)) : new_n4501_;
  assign new_n4501_ = (~new_n3415_ | ~new_n3349_ | ~new_n3546_) & (new_n4025_ | ~new_n4024_ | new_n3546_);
  assign new_n4502_ = new_n4017_ & (new_n3708_ | \i[1962]  | \i[1963] );
  assign new_n4503_ = ~new_n4504_ & (~new_n3351_ | ((new_n4506_ | ~new_n4446_) & (new_n4445_ | ~new_n4505_ | new_n4446_)));
  assign new_n4504_ = \i[1291]  & \i[1290]  & new_n3628_ & new_n3568_ & ~new_n3351_ & new_n4449_;
  assign new_n4505_ = ~new_n4447_ & new_n4019_;
  assign new_n4506_ = (~new_n4040_ | ~new_n4453_ | new_n3242_) & (~new_n4080_ | ~new_n3988_ | ~new_n3242_);
  assign new_n4507_ = ~new_n4510_ & (~new_n3351_ | ((new_n4508_ | new_n4513_ | ~new_n4087_) & (new_n4511_ | new_n4087_)));
  assign new_n4508_ = new_n4084_ & ((new_n4509_ & ~new_n3288_) | (\i[2515]  & new_n3288_ & (\i[2514]  | \i[2513] )));
  assign new_n4509_ = ~\i[2598]  & ~\i[2599]  & (~\i[2597]  | ~\i[2596] );
  assign new_n4510_ = ~new_n3351_ & new_n4093_ & new_n4058_ & new_n4065_ & (~\i[279]  | ~\i[278] );
  assign new_n4511_ = (~new_n4089_ | ~new_n3893_ | ~new_n4090_) & (new_n4512_ | \i[1383]  | ~new_n4091_ | new_n4090_);
  assign new_n4512_ = \i[1382]  & (\i[1381]  | \i[1380] );
  assign new_n4513_ = ~new_n4084_ & (~new_n4019_ | (~\i[1075]  & (~\i[1074]  | (~\i[1072]  & ~\i[1073] ))));
  assign new_n4514_ = (new_n4081_ & new_n4095_) | (~new_n4052_ & (new_n4081_ | new_n4095_));
  assign new_n4515_ = new_n4516_ ? (~new_n4524_ ^ new_n4530_) : (new_n4524_ ^ new_n4530_);
  assign new_n4516_ = new_n4007_ ? (~new_n4522_ & (new_n3221_ | ~new_n4523_ | ~new_n4062_)) : new_n4517_;
  assign new_n4517_ = (new_n4518_ | ~new_n4058_) & (new_n4019_ | ~new_n4055_ | ~new_n4453_ | new_n4058_);
  assign new_n4518_ = (new_n4519_ | new_n4061_) & (~new_n4520_ | ~new_n4060_ | ~new_n4061_);
  assign new_n4519_ = new_n4062_ ? new_n4063_ : (~\i[411]  | (~\i[409]  & ~\i[410] ));
  assign new_n4520_ = new_n4521_ & ~\i[1720]  & ~\i[1721] ;
  assign new_n4521_ = ~\i[1722]  & ~\i[1723] ;
  assign new_n4522_ = new_n4069_ & new_n3221_ & (new_n4072_ | new_n4065_);
  assign new_n4523_ = ~new_n4077_ & new_n4074_;
  assign new_n4524_ = (new_n4525_ | ~new_n3257_) & (\i[1831]  | ~new_n3990_ | ~new_n4529_ | new_n3257_);
  assign new_n4525_ = (new_n4526_ | new_n4470_) & (~new_n3775_ | ~new_n4463_ | ~new_n4528_ | ~new_n4470_);
  assign new_n4526_ = new_n4468_ ? ~new_n4527_ : ((~new_n4467_ | ~\i[487] ) & (~\i[278]  | ~\i[279]  | \i[487] ));
  assign new_n4527_ = ~new_n4192_ & new_n4098_ & (\i[397]  | \i[396] );
  assign new_n4528_ = \i[1739]  & (\i[1737]  | \i[1738]  | \i[1736] );
  assign new_n4529_ = new_n4459_ & new_n4275_ & (~\i[1830]  | ~\i[1829]  | ~\i[1828] );
  assign new_n4530_ = new_n3257_ ? new_n4531_ : ((new_n4534_ | ~new_n3677_) & (~new_n4102_ | ~new_n4103_ | new_n3677_));
  assign new_n4531_ = ~new_n4096_ & (~new_n4100_ | (~new_n4532_ & (~new_n4105_ | ~new_n4104_)));
  assign new_n4532_ = ~new_n4105_ & (new_n3782_ | new_n4533_) & (\i[413]  | \i[414]  | \i[415]  | ~new_n4533_);
  assign new_n4533_ = ~\i[1055]  & (~\i[1054]  | ~\i[1053] );
  assign new_n4534_ = ~new_n4535_ & (~new_n4424_ | ~new_n4061_ | (\i[1755]  & (\i[1753]  | \i[1754] )));
  assign new_n4535_ = \i[651]  & \i[650]  & \i[649]  & \i[648]  & ~new_n4424_ & new_n4536_;
  assign new_n4536_ = ~\i[2179]  & (~\i[2178]  | ~\i[2177] );
  assign new_n4537_ = new_n4538_ ? (~new_n4539_ ^ new_n4558_) : (new_n4539_ ^ new_n4558_);
  assign new_n4538_ = (new_n4252_ & new_n4280_) | (new_n4202_ & (new_n4252_ | new_n4280_));
  assign new_n4539_ = new_n4540_ ? (new_n4549_ ^ new_n4550_) : (~new_n4549_ ^ new_n4550_);
  assign new_n4540_ = new_n4541_ ? (new_n4542_ ^ new_n4547_) : (~new_n4542_ ^ new_n4547_);
  assign new_n4541_ = ~new_n4138_ & ~new_n4144_;
  assign new_n4542_ = new_n4345_ ? ((new_n4546_ | new_n4340_) & (new_n4339_ | ~new_n4333_ | ~new_n4340_)) : new_n4543_;
  assign new_n4543_ = new_n4219_ ? ((new_n4545_ | ~new_n4325_) & (new_n3741_ | ~new_n4326_ | new_n4325_)) : new_n4544_;
  assign new_n4544_ = (~new_n4329_ & ~new_n4330_ & new_n4265_) | (~new_n4265_ & (new_n4331_ | ~new_n3993_));
  assign new_n4545_ = (~new_n4323_ & ~new_n4324_) | (~\i[2535]  & new_n4324_ & (~\i[2534]  | ~\i[2533] ));
  assign new_n4546_ = ~new_n4344_ & (new_n4111_ | ~new_n4342_ | ~\i[2071]  | (~\i[2070]  & ~\i[2069] ));
  assign new_n4547_ = new_n3873_ ? new_n4548_ : ((~new_n4127_ | ~new_n4131_) & (~new_n3770_ | ~new_n4125_ | new_n4131_));
  assign new_n4548_ = (~new_n4118_ | new_n4135_) & (~new_n4133_ | ~new_n4136_ | ~new_n4135_);
  assign new_n4549_ = (~new_n4270_ & new_n4260_) | (new_n4253_ & (~new_n4270_ | new_n4260_));
  assign new_n4550_ = new_n4551_ ? (new_n4555_ ^ new_n4557_) : (~new_n4555_ ^ new_n4557_);
  assign new_n4551_ = (new_n4554_ & \i[1531] ) | (~new_n4552_ & ~\i[1531]  & (~new_n4044_ | ~new_n4037_));
  assign new_n4552_ = new_n4553_ & (\i[1527]  | (\i[1526]  & (\i[1525]  | \i[1524] )));
  assign new_n4553_ = ~new_n4044_ & new_n4040_ & (\i[2439]  | (\i[2437]  & \i[2438] ));
  assign new_n4554_ = (new_n3666_ | new_n4047_ | ~new_n4050_ | ~new_n4048_) & (~new_n4028_ | new_n4031_ | new_n4048_);
  assign new_n4555_ = (~new_n4168_ | (~\i[2338]  & ~\i[2339] )) & (~new_n4157_ | ~new_n4556_ | ~new_n3897_ | \i[2338]  | \i[2339] );
  assign new_n4556_ = new_n4029_ & ~\i[743]  & ~\i[1061] ;
  assign new_n4557_ = ~new_n4157_ & new_n4395_ & (\i[396]  | \i[397]  | \i[398]  | \i[399] );
  assign new_n4558_ = (~new_n4169_ & new_n4106_) | (~new_n4115_ & (~new_n4169_ | new_n4106_));
  assign new_n4559_ = new_n4560_ ? (~new_n4561_ ^ new_n4567_) : (new_n4561_ ^ new_n4567_);
  assign new_n4560_ = (~new_n4295_ & ~new_n4311_) | (~new_n4201_ & (~new_n4295_ | ~new_n4311_));
  assign new_n4561_ = new_n4562_ ? (~new_n4563_ ^ new_n4564_) : (new_n4563_ ^ new_n4564_);
  assign new_n4562_ = (~new_n4227_ & ~new_n4242_) | (~new_n4203_ & (~new_n4227_ | ~new_n4242_));
  assign new_n4563_ = (new_n4358_ & new_n4365_) | (new_n4349_ & (new_n4358_ | new_n4365_));
  assign new_n4564_ = ((new_n3373_ | ~new_n4157_ | ~new_n4264_) & (~new_n4565_ ^ ~new_n4566_)) | (~new_n3373_ & new_n4157_ & new_n4264_ & (~new_n4565_ ^ new_n4566_));
  assign new_n4565_ = new_n3564_ & new_n3467_ & new_n4257_ & new_n4044_ & ~\i[838]  & ~\i[839] ;
  assign new_n4566_ = (~new_n4317_ | ~new_n3987_) & (new_n3557_ | new_n3987_ | (\i[2187]  ? ~new_n4314_ : ~new_n4313_));
  assign new_n4567_ = (~new_n4348_ & ~new_n4374_) | (new_n4280_ & (~new_n4348_ | ~new_n4374_));
  assign new_n4568_ = (~new_n4383_ & ~new_n4399_) | (~new_n4347_ & (~new_n4383_ | ~new_n4399_));
  assign \o[9]  = ~new_n4570_ ^ new_n4571_;
  assign new_n4570_ = (~new_n4475_ & new_n4474_) | (new_n4473_ & (~new_n4475_ | new_n4474_));
  assign new_n4571_ = new_n4572_ ^ new_n4573_;
  assign new_n4572_ = (~new_n4477_ & new_n4568_) | (new_n4476_ & (~new_n4477_ | new_n4568_));
  assign new_n4573_ = new_n4574_ ? (~new_n4575_ ^ new_n4605_) : (new_n4575_ ^ new_n4605_);
  assign new_n4574_ = (~new_n4479_ & ~new_n4559_) | (new_n4478_ & (~new_n4479_ | ~new_n4559_));
  assign new_n4575_ = new_n4576_ ? (new_n4577_ ^ new_n4599_) : (~new_n4577_ ^ new_n4599_);
  assign new_n4576_ = (~new_n4481_ & ~new_n4537_) | (new_n4480_ & (~new_n4481_ | ~new_n4537_));
  assign new_n4577_ = new_n4578_ ? (new_n4582_ ^ new_n4583_) : (~new_n4582_ ^ new_n4583_);
  assign new_n4578_ = new_n4579_ ? (new_n4580_ ^ new_n4581_) : (~new_n4580_ ^ new_n4581_);
  assign new_n4579_ = (~new_n4485_ & new_n4484_) | (new_n4483_ & (~new_n4485_ | new_n4484_));
  assign new_n4580_ = (~new_n4550_ & new_n4549_) | (~new_n4540_ & (~new_n4550_ | new_n4549_));
  assign new_n4581_ = (~new_n4555_ & new_n4557_) | (~new_n4551_ & (~new_n4555_ | new_n4557_));
  assign new_n4582_ = (~new_n4497_ & new_n4496_) | (~new_n4482_ & (~new_n4497_ | new_n4496_));
  assign new_n4583_ = new_n4584_ ? (new_n4587_ ^ new_n4588_) : (~new_n4587_ ^ new_n4588_);
  assign new_n4584_ = ~new_n4585_ ^ new_n4586_;
  assign new_n4585_ = (~new_n4488_ & ~new_n4492_) | (~new_n4486_ & (~new_n4488_ | ~new_n4492_));
  assign new_n4586_ = (~new_n4503_ & ~new_n4507_) | (~new_n4499_ & (~new_n4503_ | ~new_n4507_));
  assign new_n4587_ = (~new_n4515_ & new_n4514_) | (~new_n4498_ & (~new_n4515_ | new_n4514_));
  assign new_n4588_ = new_n4589_ ? (new_n4590_ ^ new_n4596_) : (~new_n4590_ ^ new_n4596_);
  assign new_n4589_ = (~new_n4524_ & ~new_n4530_) | (~new_n4516_ & (~new_n4524_ | ~new_n4530_));
  assign new_n4590_ = (~new_n4591_ & (new_n4100_ | ~new_n4134_ | ~new_n3257_ | ~new_n4098_ | ~\i[843] )) | (~new_n4100_ & new_n4134_ & new_n3257_ & new_n4098_ & \i[843]  & new_n4591_);
  assign new_n4591_ = new_n4007_ ? new_n4592_ : (~new_n4595_ & (~new_n4594_ | ~new_n4055_ | ~new_n4019_));
  assign new_n4592_ = (new_n4593_ | ~new_n3221_) & (~new_n4080_ | ~new_n4077_ | new_n3221_ | \i[2090]  | \i[2091] );
  assign new_n4593_ = (~new_n4070_ | ~new_n4162_ | new_n4069_) & (~new_n4067_ | ~new_n4072_ | ~new_n4069_);
  assign new_n4594_ = ~new_n4058_ & (\i[640]  | \i[641]  | \i[642]  | \i[643] );
  assign new_n4595_ = new_n4060_ & new_n4061_ & new_n4058_ & new_n4520_;
  assign new_n4596_ = (~new_n4597_ & (~new_n4345_ | ~new_n4339_ | ~new_n4340_)) | (new_n4345_ & new_n4339_ & new_n4340_ & new_n4597_);
  assign new_n4597_ = new_n3257_ & (new_n4598_ | (~new_n4463_ & ~new_n4464_ & new_n4206_ & new_n4470_));
  assign new_n4598_ = new_n4192_ & new_n4468_ & ~new_n4470_ & ~new_n4469_;
  assign new_n4599_ = new_n4600_ ? (~new_n4601_ ^ new_n4602_) : (new_n4601_ ^ new_n4602_);
  assign new_n4600_ = (~new_n4539_ & new_n4558_) | (new_n4538_ & (~new_n4539_ | new_n4558_));
  assign new_n4601_ = (~new_n4564_ & new_n4563_) | (new_n4562_ & (~new_n4564_ | new_n4563_));
  assign new_n4602_ = new_n4603_ ^ new_n4604_;
  assign new_n4603_ = (~new_n4542_ & ~new_n4547_) | (new_n4541_ & (~new_n4542_ | ~new_n4547_));
  assign new_n4604_ = (~new_n4565_ | (new_n4566_ & (new_n3373_ | ~new_n4264_ | ~new_n4157_))) & (new_n4566_ | new_n3373_ | ~new_n4264_ | ~new_n4157_);
  assign new_n4605_ = (~new_n4561_ & new_n4567_) | (new_n4560_ & (~new_n4561_ | new_n4567_));
  assign \o[10]  = ((new_n4607_ | new_n4608_) & (~new_n4609_ ^ ~new_n4610_)) | (~new_n4607_ & ~new_n4608_ & (~new_n4609_ ^ new_n4610_));
  assign new_n4607_ = ~new_n4571_ & new_n4570_;
  assign new_n4608_ = ~new_n4573_ & new_n4572_;
  assign new_n4609_ = (~new_n4575_ & new_n4605_) | (new_n4574_ & (~new_n4575_ | new_n4605_));
  assign new_n4610_ = new_n4611_ ? (~new_n4612_ ^ new_n4624_) : (new_n4612_ ^ new_n4624_);
  assign new_n4611_ = (~new_n4577_ & ~new_n4599_) | (new_n4576_ & (~new_n4577_ | ~new_n4599_));
  assign new_n4612_ = new_n4613_ ? (new_n4616_ ^ new_n4617_) : (~new_n4616_ ^ new_n4617_);
  assign new_n4613_ = ~new_n4614_ ^ new_n4615_;
  assign new_n4614_ = (new_n4580_ & new_n4581_) | (new_n4579_ & (new_n4580_ | new_n4581_));
  assign new_n4615_ = ~new_n4604_ & new_n4603_;
  assign new_n4616_ = (~new_n4583_ & new_n4582_) | (~new_n4578_ & (~new_n4583_ | new_n4582_));
  assign new_n4617_ = new_n4618_ ? (~new_n4619_ ^ new_n4623_) : (new_n4619_ ^ new_n4623_);
  assign new_n4618_ = (~new_n4588_ & new_n4587_) | (~new_n4584_ & (~new_n4588_ | new_n4587_));
  assign new_n4619_ = new_n4620_ ? (~new_n4621_ ^ new_n4622_) : (new_n4621_ ^ new_n4622_);
  assign new_n4620_ = (~new_n4590_ & ~new_n4596_) | (new_n4589_ & (~new_n4590_ | ~new_n4596_));
  assign new_n4621_ = new_n4591_ & (new_n4100_ | ~new_n3257_ | ~new_n4098_ | ~new_n4134_ | ~\i[843] );
  assign new_n4622_ = new_n4340_ & new_n4339_ & new_n4597_ & new_n4345_;
  assign new_n4623_ = new_n4585_ & new_n4586_;
  assign new_n4624_ = (~new_n4602_ & new_n4601_) | (new_n4600_ & (~new_n4602_ | new_n4601_));
  assign \o[11]  = ~new_n4626_ ^ new_n4627_;
  assign new_n4626_ = (new_n4609_ | (~new_n4610_ & (new_n4608_ | new_n4607_))) & (new_n4608_ | new_n4607_ | ~new_n4610_);
  assign new_n4627_ = new_n4628_ ^ new_n4629_;
  assign new_n4628_ = (~new_n4612_ & new_n4624_) | (new_n4611_ & (~new_n4612_ | new_n4624_));
  assign new_n4629_ = new_n4630_ ? (~new_n4631_ ^ new_n4634_) : (new_n4631_ ^ new_n4634_);
  assign new_n4630_ = (~new_n4617_ & new_n4616_) | (~new_n4613_ & (~new_n4617_ | new_n4616_));
  assign new_n4631_ = ~new_n4632_ ^ new_n4633_;
  assign new_n4632_ = (~new_n4619_ & new_n4623_) | (new_n4618_ & (~new_n4619_ | new_n4623_));
  assign new_n4633_ = (~new_n4621_ & new_n4622_) | (new_n4620_ & (~new_n4621_ | new_n4622_));
  assign new_n4634_ = new_n4614_ & new_n4615_;
  assign \o[12]  = ((new_n4636_ | new_n4637_) & (~new_n4638_ ^ new_n4639_)) | (~new_n4636_ & ~new_n4637_ & (~new_n4638_ ^ ~new_n4639_));
  assign new_n4636_ = ~new_n4627_ & new_n4626_;
  assign new_n4637_ = ~new_n4629_ & new_n4628_;
  assign new_n4638_ = (~new_n4631_ & new_n4634_) | (new_n4630_ & (~new_n4631_ | new_n4634_));
  assign new_n4639_ = new_n4632_ & new_n4633_;
  assign \o[13]  = (new_n4639_ | new_n4636_ | new_n4637_) & (new_n4638_ | (new_n4639_ & (new_n4636_ | new_n4637_)));
  assign \o[14]  = new_n4642_ ^ new_n5145_;
  assign new_n4642_ = new_n4643_ ? (~new_n4795_ ^ new_n5130_) : (new_n4795_ ^ new_n5130_);
  assign new_n4643_ = new_n4644_ ? (~new_n4751_ ^ new_n4775_) : (new_n4751_ ^ new_n4775_);
  assign new_n4644_ = new_n4645_ ? (~new_n4728_ ^ new_n4743_) : (new_n4728_ ^ new_n4743_);
  assign new_n4645_ = new_n4646_ ? (~new_n4706_ ^ new_n4712_) : (new_n4706_ ^ new_n4712_);
  assign new_n4646_ = new_n4647_ ? (~new_n4669_ ^ new_n4686_) : (new_n4669_ ^ new_n4686_);
  assign new_n4647_ = new_n4667_ ? new_n4648_ : ((new_n4658_ | new_n4665_ | ~new_n4668_) & (new_n4663_ | new_n4668_));
  assign new_n4648_ = new_n4055_ ? (new_n4657_ ? new_n4652_ : new_n4655_) : new_n4649_;
  assign new_n4649_ = new_n4651_ ? new_n4650_ : ((~\i[1191]  | ~\i[2399] ) & (~\i[2270]  | ~\i[2271]  | \i[2399] ));
  assign new_n4650_ = ~new_n3268_ & (~\i[871]  | (~\i[868]  & ~\i[869]  & ~\i[870] ));
  assign new_n4651_ = ~\i[1047]  & ~\i[1046]  & ~\i[1044]  & ~\i[1045] ;
  assign new_n4652_ = (~\i[1607]  & (~\i[1605]  | ~\i[1606] )) ? new_n4653_ : new_n4654_;
  assign new_n4653_ = ~\i[2651]  & ~\i[2650]  & ~\i[2648]  & ~\i[2649] ;
  assign new_n4654_ = ~\i[515]  & (~\i[513]  | ~\i[514]  | ~\i[512] );
  assign new_n4655_ = (new_n4656_ | ~new_n4389_) & (\i[644]  | \i[645]  | \i[646]  | \i[647]  | new_n4389_);
  assign new_n4656_ = \i[1519]  & \i[1518]  & \i[1516]  & \i[1517] ;
  assign new_n4657_ = ~\i[1950]  & ~\i[1951] ;
  assign new_n4658_ = ~new_n4660_ & (new_n4662_ ? new_n4661_ : new_n4659_);
  assign new_n4659_ = new_n4299_ & ~\i[1276]  & ~\i[1277] ;
  assign new_n4660_ = ~\i[2195]  & ~\i[2193]  & ~\i[2194] ;
  assign new_n4661_ = ~\i[2219]  & ~\i[2218]  & ~\i[2216]  & ~\i[2217] ;
  assign new_n4662_ = ~\i[2615]  & ~\i[2614]  & ~\i[2612]  & ~\i[2613] ;
  assign new_n4663_ = new_n4664_ & (~\i[2327]  | (~\i[2324]  & ~\i[2325]  & ~\i[2326] ));
  assign new_n4664_ = ~\i[2763]  & ~\i[2762]  & ~\i[2760]  & ~\i[2761] ;
  assign new_n4665_ = new_n4660_ & (~new_n3399_ | ~new_n4666_) & (\i[1957]  | \i[1958]  | \i[1959]  | new_n4666_);
  assign new_n4666_ = ~\i[2291]  & ~\i[2289]  & ~\i[2290] ;
  assign new_n4667_ = ~\i[1175]  & ~\i[1173]  & ~\i[1174] ;
  assign new_n4668_ = ~\i[2635]  & (~\i[2633]  | ~\i[2634]  | ~\i[2632] );
  assign new_n4669_ = new_n4685_ ? new_n4670_ : ((~new_n4684_ & new_n4682_) | (~new_n4683_ & ~new_n4680_ & ~new_n4682_));
  assign new_n4670_ = new_n4679_ ? new_n4671_ : ~new_n4675_;
  assign new_n4671_ = new_n4674_ ? (~new_n3313_ | (~\i[2070]  & ~\i[2071] )) : new_n4672_;
  assign new_n4672_ = new_n3686_ ? new_n4673_ : ~new_n3259_;
  assign new_n4673_ = ~\i[1759]  & (~\i[1758]  | ~\i[1757] );
  assign new_n4674_ = ~\i[2410]  & ~\i[2411] ;
  assign new_n4675_ = ~new_n4676_ & ~\i[1055]  & new_n4678_ & (~\i[1054]  | ~\i[1053]  | ~\i[1052] );
  assign new_n4676_ = new_n4677_ & ~\i[1664]  & ~\i[1665] ;
  assign new_n4677_ = ~\i[1666]  & ~\i[1667] ;
  assign new_n4678_ = ~\i[1379]  & ~\i[1378]  & ~\i[1376]  & ~\i[1377] ;
  assign new_n4679_ = ~\i[1751]  & (~\i[1750]  | (~\i[1749]  & ~\i[1748] ));
  assign new_n4680_ = ~new_n4681_ & \i[2379]  & (\i[2378]  | \i[2377]  | \i[2376] );
  assign new_n4681_ = ~\i[1399]  & (~\i[1398]  | ~\i[1397] );
  assign new_n4682_ = ~\i[1967]  & (~\i[1966]  | (~\i[1965]  & ~\i[1964] ));
  assign new_n4683_ = ~\i[2391]  & (~\i[2389]  | ~\i[2390]  | ~\i[2388] );
  assign new_n4684_ = ~\i[1531]  & (~\i[1530]  | ~\i[1529] );
  assign new_n4685_ = ~\i[2034]  & ~\i[2035]  & (~\i[2033]  | ~\i[2032] );
  assign new_n4686_ = (~new_n4687_ & ~new_n4691_ & new_n4696_) | (~new_n4696_ & (new_n4702_ | (~new_n4698_ & ~\i[2399] )));
  assign new_n4687_ = ~new_n4690_ & (~new_n4689_ | new_n4055_ | ~new_n4688_) & (\i[1735]  | ~new_n3339_ | new_n4688_);
  assign new_n4688_ = ~\i[1951]  & (~\i[1949]  | ~\i[1950]  | ~\i[1948] );
  assign new_n4689_ = ~\i[1939]  & ~\i[1937]  & ~\i[1938] ;
  assign new_n4690_ = \i[610]  & \i[611] ;
  assign new_n4691_ = new_n4690_ & (new_n4695_ ? ~new_n4692_ : (~new_n4694_ | new_n3376_));
  assign new_n4692_ = new_n4693_ & (\i[1615]  | (\i[1613]  & \i[1614] ));
  assign new_n4693_ = ~\i[2051]  & ~\i[2049]  & ~\i[2050] ;
  assign new_n4694_ = ~\i[2435]  & ~\i[2434]  & ~\i[2432]  & ~\i[2433] ;
  assign new_n4695_ = \i[1079]  & (\i[1078]  | \i[1077] );
  assign new_n4696_ = new_n4697_ & (\i[1841]  | \i[1840] );
  assign new_n4697_ = \i[1842]  & \i[1843] ;
  assign new_n4698_ = (new_n4701_ | ~new_n4700_ | (~\i[2203]  & ~\i[2202] )) & (new_n4699_ | new_n3244_ | new_n4700_);
  assign new_n4699_ = \i[1851]  & (\i[1850]  | (\i[1849]  & \i[1848] ));
  assign new_n4700_ = \i[715]  & \i[714]  & \i[712]  & \i[713] ;
  assign new_n4701_ = ~\i[1851]  & ~\i[1850]  & ~\i[1848]  & ~\i[1849] ;
  assign new_n4702_ = \i[2409]  & \i[2399]  & new_n4705_ & new_n4703_ & new_n4704_;
  assign new_n4703_ = \i[1307]  & (\i[1306]  | (\i[1305]  & \i[1304] ));
  assign new_n4704_ = ~\i[2307]  & ~\i[2306]  & ~\i[2304]  & ~\i[2305] ;
  assign new_n4705_ = \i[2410]  & \i[2411] ;
  assign new_n4706_ = (~new_n4711_ & \i[593]  & \i[594]  & \i[595] ) | (new_n4707_ & (~\i[593]  | ~\i[594]  | ~\i[595] ));
  assign new_n4707_ = new_n4667_ ? ~new_n4708_ : ((new_n4080_ | new_n4710_ | ~new_n4398_) & (~new_n4709_ | new_n4398_));
  assign new_n4708_ = \i[1387]  & \i[1386]  & ~\i[1275]  & new_n4437_;
  assign new_n4709_ = (~new_n3467_ | (~\i[1555]  & (~\i[1553]  | ~\i[1554] ))) & (\i[2006]  | \i[2007]  | \i[1555]  | (\i[1553]  & \i[1554] ));
  assign new_n4710_ = \i[947]  & (\i[946]  | \i[945] );
  assign new_n4711_ = new_n4087_ & ~\i[1531]  & ~\i[2215] ;
  assign new_n4712_ = new_n4726_ ? (~new_n4720_ & (new_n4725_ | new_n4727_ | ~new_n3473_)) : new_n4713_;
  assign new_n4713_ = (new_n4714_ | new_n4718_) & (\i[2087]  | ~new_n4719_ | ~new_n4718_ | (\i[2086]  & \i[2085] ));
  assign new_n4714_ = (new_n4715_ & ~new_n4716_) | (new_n4717_ & new_n4716_ & (~\i[2165]  | ~new_n3431_));
  assign new_n4715_ = ~\i[1713]  & ~\i[1714]  & ~\i[1715]  & \i[1619]  & (\i[1618]  | \i[1617] );
  assign new_n4716_ = \i[1946]  & \i[1947]  & (\i[1945]  | \i[1944] );
  assign new_n4717_ = ~\i[1839]  & (~\i[1837]  | ~\i[1838]  | ~\i[1836] );
  assign new_n4718_ = \i[2758]  & \i[2759]  & (\i[2757]  | \i[2756] );
  assign new_n4719_ = ~\i[959]  & (~\i[958]  | ~\i[957] );
  assign new_n4720_ = ~new_n4721_ & new_n4725_ & (new_n4724_ | ~new_n4723_ | ~new_n4722_);
  assign new_n4721_ = ~new_n4722_ & (new_n4047_ ? (~new_n3890_ | (\i[1208]  & \i[1209] )) : ~new_n3229_);
  assign new_n4722_ = ~\i[959]  & ~\i[958]  & ~\i[956]  & ~\i[957] ;
  assign new_n4723_ = \i[1303]  & (\i[1302]  | \i[1301] );
  assign new_n4724_ = ~\i[831]  & ~\i[830]  & ~\i[828]  & ~\i[829] ;
  assign new_n4725_ = ~\i[2647]  & ~\i[2646]  & ~\i[2644]  & ~\i[2645] ;
  assign new_n4726_ = \i[1867]  & (\i[1866]  | (\i[1865]  & \i[1864] ));
  assign new_n4727_ = ~\i[923]  & ~\i[922]  & ~\i[920]  & ~\i[921] ;
  assign new_n4728_ = new_n4742_ ? new_n4729_ : new_n4738_;
  assign new_n4729_ = (\i[1043]  | ~new_n3274_ | ~new_n4734_ | new_n4737_) & (~new_n4737_ | (~new_n4736_ & ~new_n4730_));
  assign new_n4730_ = new_n4733_ & (new_n4732_ | new_n4731_) & (\i[1545]  | \i[1546]  | \i[1547]  | ~new_n4731_);
  assign new_n4731_ = new_n4268_ & ~\i[2324]  & ~\i[2325] ;
  assign new_n4732_ = ~\i[487]  & ~\i[486]  & ~\i[484]  & ~\i[485] ;
  assign new_n4733_ = ~\i[2555]  & ~\i[2554]  & ~\i[2552]  & ~\i[2553] ;
  assign new_n4734_ = new_n4735_ & ~\i[2532]  & ~\i[2533] ;
  assign new_n4735_ = ~\i[2534]  & ~\i[2535] ;
  assign new_n4736_ = ~new_n4733_ & ~new_n4091_ & (\i[835]  | (\i[833]  & \i[834] ));
  assign new_n4737_ = ~\i[1995]  & ~\i[1993]  & ~\i[1994] ;
  assign new_n4738_ = (~new_n4739_ & new_n4741_) | (~\i[495]  & ~new_n4741_ & (~\i[494]  | ~\i[493] ));
  assign new_n4739_ = new_n4740_ & (~\i[2101]  | ~\i[2100] );
  assign new_n4740_ = ~\i[2102]  & ~\i[2103] ;
  assign new_n4741_ = \i[2535]  & (\i[2534]  | \i[2533] );
  assign new_n4742_ = ~\i[486]  & ~\i[487]  & (~\i[485]  | ~\i[484] );
  assign new_n4743_ = (\i[593]  & \i[594]  & \i[595] ) ? (new_n4749_ | ~new_n4087_) : new_n4744_;
  assign new_n4744_ = (new_n4667_ | (~new_n4748_ & (new_n4398_ | new_n4709_))) & (new_n4745_ | new_n4747_ | ~new_n4667_);
  assign new_n4745_ = new_n4437_ & ((~new_n4746_ & \i[1275] ) | (\i[1386]  & \i[1387]  & ~\i[1275] ));
  assign new_n4746_ = \i[2498]  & \i[2499]  & (\i[2497]  | \i[2496] );
  assign new_n4747_ = ~new_n3546_ & ~new_n4437_ & ~\i[511]  & (~\i[510]  | (~\i[508]  & ~\i[509] ));
  assign new_n4748_ = \i[2431]  & \i[2430]  & new_n4398_ & new_n4080_ & new_n4153_;
  assign new_n4749_ = (~\i[1531]  & ~\i[2215] ) | (~new_n4750_ & ~new_n3513_ & \i[2215] );
  assign new_n4750_ = \i[2187]  & (\i[2186]  | (\i[2185]  & \i[2184] ));
  assign new_n4751_ = new_n4774_ ? ((~new_n4765_ | ~new_n4219_) & (new_n4770_ | new_n4773_ | new_n4219_)) : new_n4752_;
  assign new_n4752_ = new_n3275_ ? new_n4753_ : ((new_n4758_ | ~new_n4764_) & (new_n4761_ | new_n4763_ | new_n4764_));
  assign new_n4753_ = (~new_n4754_ | new_n4756_) & (~new_n4755_ | (new_n4757_ ? new_n4021_ : ~new_n4207_));
  assign new_n4754_ = ~new_n4755_ & ~\i[1615]  & (~\i[1614]  | ~\i[1613] );
  assign new_n4755_ = ~\i[2610]  & ~\i[2611] ;
  assign new_n4756_ = ~\i[2735]  & ~\i[2733]  & ~\i[2734] ;
  assign new_n4757_ = ~\i[1163]  & ~\i[1162]  & ~\i[1160]  & ~\i[1161] ;
  assign new_n4758_ = new_n4760_ ? ~new_n4759_ : ~new_n4676_;
  assign new_n4759_ = ~\i[1155]  & ~\i[1154]  & ~\i[1152]  & ~\i[1153] ;
  assign new_n4760_ = \i[1483]  & (\i[1482]  | \i[1481] );
  assign new_n4761_ = ~new_n4762_ & ~\i[2647]  & (~\i[2646]  | ~\i[2645]  | ~\i[2644] );
  assign new_n4762_ = \i[1051]  & (\i[1049]  | \i[1050]  | \i[1048] );
  assign new_n4763_ = new_n4762_ & \i[747]  & (\i[746]  | \i[745]  | \i[744] );
  assign new_n4764_ = ~\i[2722]  & ~\i[2723] ;
  assign new_n4765_ = new_n4769_ ? new_n4766_ : (new_n3310_ ? \i[483]  : ~new_n4091_);
  assign new_n4766_ = new_n4767_ ? (\i[1635]  | (\i[1633]  & \i[1634] )) : new_n4768_;
  assign new_n4767_ = \i[1835]  & (\i[1833]  | \i[1834]  | \i[1832] );
  assign new_n4768_ = ~\i[2279]  & ~\i[2277]  & ~\i[2278] ;
  assign new_n4769_ = ~\i[1531]  & ~\i[1529]  & ~\i[1530] ;
  assign new_n4770_ = new_n4772_ & (~new_n4771_ | ~\i[2074]  | ~\i[2075]  | (~\i[2073]  & ~\i[2072] ));
  assign new_n4771_ = ~\i[2330]  & ~\i[2331]  & (~\i[2329]  | ~\i[2328] );
  assign new_n4772_ = \i[1410]  & \i[1411]  & (\i[1409]  | \i[1408] );
  assign new_n4773_ = ~new_n4772_ & new_n3736_ & \i[1279]  & (\i[1278]  | \i[1277]  | \i[1276] );
  assign new_n4774_ = ~\i[2063]  & ~\i[2061]  & ~\i[2062] ;
  assign new_n4775_ = (new_n4776_ & new_n3736_) | (~new_n4786_ & ~new_n3736_ & (~new_n4793_ | new_n4791_));
  assign new_n4776_ = new_n3697_ ? ((new_n4785_ & ~new_n4784_) | (~new_n3258_ & new_n4783_ & new_n4784_)) : new_n4777_;
  assign new_n4777_ = (new_n4778_ | ~new_n3615_) & (new_n3365_ | ~new_n4781_ | ~new_n4782_ | new_n3615_);
  assign new_n4778_ = (~new_n4779_ | ~new_n4780_) & (~\i[2626]  | ~\i[2627]  | new_n4780_ | (~\i[2625]  & ~\i[2624] ));
  assign new_n4779_ = ~\i[2183]  & ~\i[2182]  & ~\i[2180]  & ~\i[2181] ;
  assign new_n4780_ = ~\i[1371]  & ~\i[1370]  & ~\i[1368]  & ~\i[1369] ;
  assign new_n4781_ = \i[966]  & \i[967] ;
  assign new_n4782_ = \i[964]  & \i[965] ;
  assign new_n4783_ = ~\i[2107]  & ~\i[2106]  & ~\i[2104]  & ~\i[2105] ;
  assign new_n4784_ = ~\i[1559]  & ~\i[1558]  & ~\i[1556]  & ~\i[1557] ;
  assign new_n4785_ = ~\i[1179]  & ~\i[1177]  & ~\i[1178] ;
  assign new_n4786_ = ~new_n4787_ & new_n4788_ & (new_n3585_ | (new_n4790_ & ~new_n4789_) | (new_n3257_ & new_n4789_));
  assign new_n4787_ = ~new_n4757_ & new_n3585_ & ((~\i[2436]  & ~\i[2437] ) | ~\i[2439]  | ~\i[2438] );
  assign new_n4788_ = ~\i[1291]  & (~\i[1289]  | ~\i[1290]  | ~\i[1288] );
  assign new_n4789_ = \i[2635]  & (\i[2633]  | \i[2634]  | \i[2632] );
  assign new_n4790_ = \i[1183]  & (\i[1182]  | \i[1181] );
  assign new_n4791_ = ~new_n4190_ & (new_n4792_ | ~\i[2427]  | (~\i[2426]  & (~\i[2424]  | ~\i[2425] )));
  assign new_n4792_ = \i[1427]  & \i[1426]  & \i[1424]  & \i[1425] ;
  assign new_n4793_ = ~new_n4788_ & (new_n4794_ | \i[2089]  | \i[2090]  | \i[2091]  | ~new_n4190_);
  assign new_n4794_ = \i[2423]  & (\i[2421]  | \i[2422]  | \i[2420] );
  assign new_n4795_ = new_n4796_ ? (~new_n4922_ ^ new_n5111_) : (new_n4922_ ^ new_n5111_);
  assign new_n4796_ = new_n4797_ ? (~new_n4886_ ^ new_n4909_) : (new_n4886_ ^ new_n4909_);
  assign new_n4797_ = new_n4798_ ? (~new_n4852_ ^ new_n4706_) : (new_n4852_ ^ new_n4706_);
  assign new_n4798_ = new_n4799_ ? (~new_n4825_ ^ new_n4838_) : (new_n4825_ ^ new_n4838_);
  assign new_n4799_ = new_n3258_ ? new_n4800_ : ((new_n4811_ | ~new_n4821_) & (new_n4815_ | new_n4822_ | new_n4821_));
  assign new_n4800_ = new_n4165_ ? ((new_n4807_ | ~new_n4809_) & (\i[1299]  | ~new_n4810_ | new_n4809_)) : new_n4801_;
  assign new_n4801_ = (new_n4802_ | (new_n4806_ ? ~new_n4805_ : new_n4206_)) & (new_n3349_ | ~new_n4804_ | ~new_n4802_);
  assign new_n4802_ = \i[2749]  & new_n4803_ & \i[2748] ;
  assign new_n4803_ = \i[2750]  & \i[2751] ;
  assign new_n4804_ = ~\i[1835]  & ~\i[1834]  & ~\i[1832]  & ~\i[1833] ;
  assign new_n4805_ = ~\i[963]  & ~\i[962]  & ~\i[960]  & ~\i[961] ;
  assign new_n4806_ = ~\i[2274]  & ~\i[2275] ;
  assign new_n4807_ = (new_n3613_ & (\i[2726]  | \i[2727] )) | (\i[1603]  & ~\i[2726]  & ~\i[2727]  & (\i[1602]  | ~new_n4808_));
  assign new_n4808_ = ~\i[1600]  & ~\i[1601] ;
  assign new_n4809_ = ~\i[403]  & ~\i[402]  & ~\i[400]  & ~\i[401] ;
  assign new_n4810_ = ~\i[1651]  & ~\i[1650]  & ~\i[1648]  & ~\i[1649] ;
  assign new_n4811_ = new_n4814_ ? (new_n4813_ ? new_n4315_ : ~new_n4078_) : new_n4812_;
  assign new_n4812_ = (~\i[845]  | ~new_n4289_ | ~\i[844] ) & (\i[1183]  | \i[1182] );
  assign new_n4813_ = ~\i[623]  & (~\i[621]  | ~\i[622]  | ~\i[620] );
  assign new_n4814_ = \i[1959]  & (\i[1957]  | \i[1958]  | \i[1956] );
  assign new_n4815_ = new_n4818_ & (new_n4816_ ? new_n4819_ : new_n4820_);
  assign new_n4816_ = \i[1719]  & (\i[1718]  | new_n4817_);
  assign new_n4817_ = \i[1716]  & \i[1717] ;
  assign new_n4818_ = ~\i[958]  & ~\i[959]  & (~\i[957]  | ~\i[956] );
  assign new_n4819_ = ~\i[2159]  & ~\i[2157]  & ~\i[2158] ;
  assign new_n4820_ = \i[1639]  & (\i[1637]  | \i[1638]  | \i[1636] );
  assign new_n4821_ = \i[1073]  & new_n4379_ & \i[1072] ;
  assign new_n4822_ = ~new_n4818_ & ((~new_n4824_ & new_n4823_) | (~\i[2441]  & ~\i[2442]  & ~\i[2443]  & ~new_n4823_));
  assign new_n4823_ = \i[2103]  & (\i[2102]  | \i[2101] );
  assign new_n4824_ = ~\i[2431]  & (~\i[2430]  | ~\i[2429] );
  assign new_n4825_ = new_n4836_ ? ((new_n4826_ & new_n4837_) | (~new_n4829_ & ~new_n4834_ & ~new_n4837_)) : ~new_n4832_;
  assign new_n4826_ = (\i[1482]  | \i[1483]  | (~\i[1773]  & new_n3799_)) & (new_n4827_ | new_n4828_ | \i[1773]  | ~new_n3799_);
  assign new_n4827_ = ~\i[2094]  & ~\i[2095]  & (~new_n3855_ | (\i[1852]  & \i[1853] ));
  assign new_n4828_ = new_n3855_ & \i[1981]  & \i[1982]  & \i[1983]  & (~\i[1853]  | ~\i[1852] );
  assign new_n4829_ = ~new_n4830_ & (~\i[1599]  | (~\i[1597]  & ~\i[1598] ));
  assign new_n4830_ = (~new_n4831_ | ~\i[507] ) & (~\i[2101]  | ~\i[2102]  | ~\i[2103]  | \i[507] );
  assign new_n4831_ = ~\i[1275]  & ~\i[1273]  & ~\i[1274] ;
  assign new_n4832_ = ~\i[1818]  & ~\i[1819]  & new_n4833_ & (~\i[1817]  | ~\i[1816] );
  assign new_n4833_ = \i[1854]  & \i[1855]  & (\i[1853]  | \i[1852] );
  assign new_n4834_ = \i[1599]  & (\i[1597]  | \i[1598] ) & (new_n3422_ ? ~new_n4386_ : ~new_n4835_);
  assign new_n4835_ = ~\i[1858]  & ~\i[1859]  & (~\i[1857]  | ~\i[1856] );
  assign new_n4836_ = ~\i[1479]  & (~\i[1477]  | ~\i[1478]  | ~\i[1476] );
  assign new_n4837_ = ~\i[1499]  & (~\i[1497]  | ~\i[1498]  | ~\i[1496] );
  assign new_n4838_ = new_n4850_ ? new_n4839_ : ((new_n4844_ | ~new_n3479_) & (new_n4846_ | new_n4849_ | new_n3479_));
  assign new_n4839_ = new_n4841_ ? ((~new_n4843_ & ~new_n4842_) | (~new_n4681_ & new_n4694_ & new_n4842_)) : new_n4840_;
  assign new_n4840_ = ~new_n3606_ & ((~\i[2617]  & ~\i[2616] ) | ~\i[2619]  | ~\i[2618] );
  assign new_n4841_ = ~\i[1487]  & (~\i[1485]  | ~\i[1486]  | ~\i[1484] );
  assign new_n4842_ = ~\i[1887]  & ~\i[1886]  & ~\i[1884]  & ~\i[1885] ;
  assign new_n4843_ = ~\i[1591]  & (~\i[1590]  | (~\i[1589]  & ~\i[1588] ));
  assign new_n4844_ = (\i[1055]  | new_n3548_ | ~new_n4845_) & (~\i[1711]  | new_n4845_ | (~\i[1710]  & ~new_n3397_));
  assign new_n4845_ = \i[1823]  & (\i[1822]  | \i[1821] );
  assign new_n4846_ = ~new_n4847_ & (new_n4848_ ? (\i[2753]  | ~new_n3849_) : ~new_n4100_);
  assign new_n4847_ = \i[1841]  & new_n4697_ & \i[1840] ;
  assign new_n4848_ = \i[2407]  & \i[2405]  & \i[2406] ;
  assign new_n4849_ = new_n4847_ & (~new_n3392_ | (\i[1611]  & (\i[1608]  | \i[1609]  | \i[1610] )));
  assign new_n4850_ = new_n4851_ & (~\i[1381]  | ~\i[1380] );
  assign new_n4851_ = ~\i[1382]  & ~\i[1383] ;
  assign new_n4852_ = new_n4853_ ? (new_n4866_ ^ new_n4882_) : (~new_n4866_ ^ new_n4882_);
  assign new_n4853_ = new_n4865_ ? new_n4854_ : ~new_n4864_;
  assign new_n4854_ = ~new_n4855_ & (~\i[1378]  | ~\i[1379]  | (new_n4862_ ? ~new_n4863_ : new_n4860_));
  assign new_n4855_ = new_n4857_ & (new_n4858_ | (~\i[2114]  & ~\i[2115]  & new_n4856_) | (\i[2211]  & ~new_n4856_));
  assign new_n4856_ = new_n3510_ & (~\i[2529]  | ~\i[2528] );
  assign new_n4857_ = (~\i[1379]  | ~\i[1378] ) & (\i[743]  | new_n4859_ | ~new_n4858_);
  assign new_n4858_ = ~\i[1886]  & ~\i[1887]  & (~\i[1885]  | ~\i[1884] );
  assign new_n4859_ = ~\i[1087]  & (~\i[1086]  | (~\i[1085]  & ~\i[1084] ));
  assign new_n4860_ = (~\i[1539]  & (~\i[1538]  | (~\i[1536]  & ~\i[1537] ))) ? ~\i[943]  : ~new_n4861_;
  assign new_n4861_ = \i[866]  & \i[867] ;
  assign new_n4862_ = ~\i[1279]  & (~\i[1278]  | ~\i[1277] );
  assign new_n4863_ = ~\i[1267]  & (~\i[1266]  | (~\i[1265]  & ~\i[1264] ));
  assign new_n4864_ = \i[1966]  & \i[1967]  & (\i[1965]  | \i[1964] );
  assign new_n4865_ = ~\i[1474]  & ~\i[1475]  & (~\i[1473]  | ~\i[1472] );
  assign new_n4866_ = new_n4881_ ? (new_n4392_ ? new_n4873_ : new_n4876_) : new_n4867_;
  assign new_n4867_ = (~new_n4275_ & (\i[1554]  | \i[1555] )) | (~\i[1554]  & ~\i[1555]  & (new_n4268_ ? new_n4868_ : new_n4871_));
  assign new_n4868_ = new_n4869_ ? (~\i[979]  | (~\i[976]  & ~\i[977]  & ~\i[978] )) : ~new_n4870_;
  assign new_n4869_ = \i[1095]  & (\i[1094]  | (\i[1093]  & \i[1092] ));
  assign new_n4870_ = \i[1991]  & (\i[1990]  | \i[1989] );
  assign new_n4871_ = (~\i[1991]  & (~\i[1990]  | (~\i[1988]  & ~\i[1989] ))) ? ~new_n4872_ : ~new_n4446_;
  assign new_n4872_ = ~\i[2655]  & ~\i[2654]  & ~\i[2652]  & ~\i[2653] ;
  assign new_n4873_ = new_n4875_ ? ((~\i[1419]  | \i[511] ) & (~\i[2066]  | ~\i[2067]  | ~\i[511] )) : new_n4874_;
  assign new_n4874_ = (new_n4818_ | ~new_n4654_) & (\i[2203]  | new_n4654_ | (\i[2202]  & (\i[2200]  | \i[2201] )));
  assign new_n4875_ = \i[855]  & \i[853]  & \i[854] ;
  assign new_n4876_ = (~new_n4878_ | ~new_n4879_ | new_n4877_) & (~new_n4877_ | (new_n4880_ ? new_n4657_ : new_n3585_));
  assign new_n4877_ = \i[635]  & (\i[634]  | \i[633] );
  assign new_n4878_ = ~\i[979]  & ~\i[977]  & ~\i[978] ;
  assign new_n4879_ = \i[2179]  & \i[2177]  & \i[2178] ;
  assign new_n4880_ = \i[1523]  & \i[1522]  & \i[1520]  & \i[1521] ;
  assign new_n4881_ = ~\i[1179]  & (~\i[1177]  | ~\i[1178]  | ~\i[1176] );
  assign new_n4882_ = (\i[381]  | \i[382]  | ~\i[383] ) & (new_n4883_ | new_n4885_ | \i[383] );
  assign new_n4883_ = new_n4884_ & new_n3728_ & (\i[2087]  | (\i[2086]  & (\i[2085]  | \i[2084] )));
  assign new_n4884_ = ~\i[1827]  & (~\i[1826]  | ~\i[1825] );
  assign new_n4885_ = ~new_n3728_ & ((\i[1051]  & \i[1050] ) | (~\i[2709]  & ~\i[2710]  & ~\i[2711] ));
  assign new_n4886_ = (new_n4887_ & \i[628]  & \i[629]  & \i[630]  & \i[631] ) | (new_n4897_ & (~\i[628]  | ~\i[629]  | ~\i[630]  | ~\i[631] ));
  assign new_n4887_ = (\i[2499]  & (\i[2497]  | \i[2498] )) ? new_n4888_ : new_n4893_;
  assign new_n4888_ = (~new_n3940_ & \i[1843] ) ? new_n4892_ : new_n4889_;
  assign new_n4889_ = (new_n4058_ | ~new_n4890_) & (\i[1189]  | \i[1190]  | \i[1191]  | new_n4890_);
  assign new_n4890_ = \i[2285]  & new_n4891_ & \i[2284] ;
  assign new_n4891_ = \i[2286]  & \i[2287] ;
  assign new_n4892_ = \i[1398]  & \i[1399]  & \i[1397]  & (~\i[2423]  | (~\i[2421]  & ~\i[2422] ));
  assign new_n4893_ = (new_n4894_ & (~new_n4705_ | ~\i[2408]  | ~\i[2409] )) | (new_n4896_ & new_n4705_ & \i[2408]  & \i[2409] );
  assign new_n4894_ = (new_n3770_ | new_n4895_) & (~\i[862]  | ~\i[863]  | ~new_n4895_ | (~\i[861]  & ~\i[860] ));
  assign new_n4895_ = ~\i[855]  & ~\i[853]  & ~\i[854] ;
  assign new_n4896_ = new_n3281_ ? ~\i[1511]  : (~\i[1039]  | (~\i[1038]  & ~\i[1037] ));
  assign new_n4897_ = ~new_n4898_ & (~new_n3416_ | (~new_n4906_ & ~new_n4905_) | (~new_n4329_ & new_n4440_ & new_n4905_));
  assign new_n4898_ = ~new_n4899_ & ~new_n3416_ & (new_n4900_ | (~new_n4904_ & new_n4902_) | (~new_n4903_ & ~new_n4902_));
  assign new_n4899_ = new_n4901_ & new_n4900_ & (~\i[2047]  | (~\i[2044]  & ~\i[2045]  & ~\i[2046] ));
  assign new_n4900_ = \i[739]  & \i[738]  & \i[736]  & \i[737] ;
  assign new_n4901_ = ~\i[2507]  & ~\i[2506]  & ~\i[2504]  & ~\i[2505] ;
  assign new_n4902_ = ~\i[1407]  & (~\i[1405]  | ~\i[1406]  | ~\i[1404] );
  assign new_n4903_ = ~\i[2859]  & (~\i[2857]  | ~\i[2858]  | ~\i[2856] );
  assign new_n4904_ = ~\i[2275]  & (~\i[2273]  | ~\i[2274]  | ~\i[2272] );
  assign new_n4905_ = new_n4075_ & (\i[1961]  | \i[1960] );
  assign new_n4906_ = (~new_n4907_ & ~\i[1310]  & ~\i[1311]  & (~\i[1308]  | ~\i[1309] )) | (new_n4908_ & (\i[1310]  | \i[1311]  | (\i[1308]  & \i[1309] )));
  assign new_n4907_ = \i[2311]  & (\i[2309]  | \i[2310]  | \i[2308] );
  assign new_n4908_ = \i[523]  & (\i[521]  | \i[522]  | \i[520] );
  assign new_n4909_ = new_n3728_ ? ((new_n4921_ | ~new_n3606_) & (~new_n4919_ | ~new_n4920_ | new_n3606_)) : new_n4910_;
  assign new_n4910_ = (new_n4911_ | new_n4918_) & (new_n4914_ | new_n4917_ | ~new_n4918_);
  assign new_n4911_ = (~new_n3606_ | new_n3497_ | new_n4913_) & (~new_n4913_ | (new_n4704_ ? new_n4912_ : new_n3896_));
  assign new_n4912_ = ~\i[2518]  & ~\i[2519]  & (~\i[2517]  | ~\i[2516] );
  assign new_n4913_ = ~\i[1491]  & (~\i[1490]  | ~\i[1489] );
  assign new_n4914_ = ~new_n4694_ & (new_n4915_ ? new_n4916_ : (~\i[2199]  | ~\i[2198] ));
  assign new_n4915_ = ~\i[1991]  & ~\i[1990]  & ~\i[1988]  & ~\i[1989] ;
  assign new_n4916_ = \i[2655]  & (\i[2654]  | \i[2653] );
  assign new_n4917_ = ~\i[2103]  & new_n4694_ & new_n4872_ & (~\i[2102]  | (~\i[2100]  & ~\i[2101] ));
  assign new_n4918_ = ~\i[1779]  & (~\i[1778]  | ~\i[1777] );
  assign new_n4919_ = ~\i[1823]  & ~\i[1822]  & ~\i[1820]  & ~\i[1821] ;
  assign new_n4920_ = \i[1855]  & (\i[1854]  | \i[1853] );
  assign new_n4921_ = ~\i[2043]  & ~\i[2041]  & ~\i[2042] ;
  assign new_n4922_ = new_n4923_ ? (~new_n5000_ ^ new_n5103_) : (new_n5000_ ^ new_n5103_);
  assign new_n4923_ = new_n4924_ ? (new_n4988_ ^ new_n4999_) : (~new_n4988_ ^ new_n4999_);
  assign new_n4924_ = new_n4925_ ? (~new_n4943_ ^ new_n4969_) : (new_n4943_ ^ new_n4969_);
  assign new_n4925_ = new_n4837_ ? (\i[1519]  ? new_n4934_ : new_n4940_) : new_n4926_;
  assign new_n4926_ = (new_n4927_ | \i[1599]  | (\i[1597]  & \i[1598] )) & (new_n4931_ | new_n4933_ | (~\i[1599]  & (~\i[1597]  | ~\i[1598] )));
  assign new_n4927_ = (new_n4928_ & ~new_n4930_) | (new_n4732_ & new_n4930_ & (~\i[623]  | ~\i[622] ));
  assign new_n4928_ = new_n4929_ & ((~\i[1997]  & ~\i[1996] ) | ~\i[1999]  | ~\i[1998] );
  assign new_n4929_ = ~\i[419]  & ~\i[418]  & ~\i[416]  & ~\i[417] ;
  assign new_n4930_ = ~\i[1731]  & (~\i[1729]  | ~\i[1730]  | ~\i[1728] );
  assign new_n4931_ = ~\i[2109]  & ~\i[2110]  & ~\i[2111]  & \i[1167]  & (\i[1166]  | ~new_n4932_);
  assign new_n4932_ = ~\i[1164]  & ~\i[1165] ;
  assign new_n4933_ = (\i[1038]  | \i[1039]  | \i[1037] ) & (~\i[1167]  | (~\i[1166]  & new_n4932_));
  assign new_n4934_ = new_n3985_ ? new_n4935_ : (new_n4303_ ? new_n3219_ : new_n4939_);
  assign new_n4935_ = new_n4938_ ? new_n4936_ : ~new_n4461_;
  assign new_n4936_ = new_n4937_ & ~\i[2196]  & ~\i[2197] ;
  assign new_n4937_ = ~\i[2198]  & ~\i[2199] ;
  assign new_n4938_ = new_n3491_ & ~\i[2640]  & ~\i[2641] ;
  assign new_n4939_ = ~\i[2443]  & ~\i[2442]  & ~\i[2440]  & ~\i[2441] ;
  assign new_n4940_ = \i[1487]  ? new_n4941_ : (new_n4666_ ? new_n4134_ : ~new_n3849_);
  assign new_n4941_ = (~\i[1499]  & new_n4942_ & ~new_n3311_) | (new_n3311_ & (~new_n4891_ | (~\i[2285]  & ~\i[2284] )));
  assign new_n4942_ = ~\i[1497]  & ~\i[1498] ;
  assign new_n4943_ = (new_n4944_ | new_n4951_ | new_n4968_) & (~new_n4968_ | (~new_n4959_ & (new_n4964_ | ~new_n4967_)));
  assign new_n4944_ = ~new_n3275_ & ((~new_n4945_ & new_n4948_) | (~new_n4950_ & new_n3527_ & ~new_n4948_));
  assign new_n4945_ = (~\i[1203]  | ~new_n4946_) & (\i[2756]  | \i[2757]  | \i[2758]  | \i[2759]  | new_n4946_);
  assign new_n4946_ = new_n4947_ & ~\i[856]  & ~\i[857] ;
  assign new_n4947_ = ~\i[858]  & ~\i[859] ;
  assign new_n4948_ = new_n4949_ & ~\i[2312]  & ~\i[2313] ;
  assign new_n4949_ = ~\i[2314]  & ~\i[2315] ;
  assign new_n4950_ = ~\i[1979]  & ~\i[1978]  & ~\i[1976]  & ~\i[1977] ;
  assign new_n4951_ = new_n3275_ & (new_n4956_ ? new_n4952_ : (new_n4958_ | new_n4957_));
  assign new_n4952_ = new_n4954_ ? ~new_n4953_ : new_n4955_;
  assign new_n4953_ = ~\i[947]  & (~\i[945]  | ~\i[946]  | ~\i[944] );
  assign new_n4954_ = \i[1727]  & (\i[1725]  | \i[1726]  | \i[1724] );
  assign new_n4955_ = ~\i[1751]  & ~\i[1749]  & ~\i[1750] ;
  assign new_n4956_ = ~\i[2611]  & (~\i[2610]  | (~\i[2609]  & ~\i[2608] ));
  assign new_n4957_ = \i[2191]  & (\i[2189]  | \i[2190]  | \i[2188] );
  assign new_n4958_ = \i[1407]  & (\i[1406]  | \i[1405] );
  assign new_n4959_ = new_n4963_ & (new_n4962_ | new_n4961_) & (new_n4960_ | ~\i[862]  | ~\i[863]  | ~new_n4961_);
  assign new_n4960_ = new_n4000_ & (~\i[753]  | ~\i[752] );
  assign new_n4961_ = ~\i[1263]  & (~\i[1262]  | (~\i[1261]  & ~\i[1260] ));
  assign new_n4962_ = \i[1763]  & \i[1762]  & \i[1760]  & \i[1761] ;
  assign new_n4963_ = \i[2043]  & (\i[2042]  | (\i[2041]  & \i[2040] ));
  assign new_n4964_ = new_n4966_ & ((~new_n3303_ & new_n4965_) | (\i[859]  & ~new_n4965_ & (\i[858]  | \i[857] )));
  assign new_n4965_ = ~\i[715]  & (~\i[713]  | ~\i[714]  | ~\i[712] );
  assign new_n4966_ = ~\i[1843]  & (~\i[1842]  | (~\i[1841]  & ~\i[1840] ));
  assign new_n4967_ = ~new_n4963_ & (new_n4966_ | ((~new_n3669_ | ~new_n4289_) & (~\i[1634]  | ~\i[1635]  | new_n4289_)));
  assign new_n4968_ = ~\i[2171]  & ~\i[2169]  & ~\i[2170] ;
  assign new_n4969_ = (new_n4974_ | ~new_n4820_) & (new_n4970_ | new_n4984_ | new_n4820_);
  assign new_n4970_ = new_n4971_ & (new_n4973_ ? ~new_n3233_ : (~\i[1755]  | (~\i[1753]  & ~\i[1754] )));
  assign new_n4971_ = ~new_n4972_ & \i[1419]  & (\i[1418]  | \i[1417]  | \i[1416] );
  assign new_n4972_ = \i[1947]  & \i[1946]  & \i[1944]  & \i[1945] ;
  assign new_n4973_ = \i[1955]  & \i[1954]  & \i[1952]  & \i[1953] ;
  assign new_n4974_ = (new_n4982_ | new_n4978_ | new_n3905_) & (new_n4975_ | new_n4983_ | ~new_n3905_);
  assign new_n4975_ = new_n4976_ ? ~new_n4977_ : ~new_n4300_;
  assign new_n4976_ = \i[1543]  & (\i[1541]  | \i[1542]  | \i[1540] );
  assign new_n4977_ = ~\i[943]  & ~\i[942]  & ~\i[940]  & ~\i[941] ;
  assign new_n4978_ = ~new_n4979_ & ((\i[2767]  & ~new_n4981_ & (\i[2766]  | \i[2765] )) | (~new_n4980_ & new_n4981_));
  assign new_n4979_ = ~\i[2547]  & ~\i[2546]  & ~\i[2544]  & ~\i[2545] ;
  assign new_n4980_ = ~\i[2543]  & (~\i[2542]  | (~\i[2541]  & ~\i[2540] ));
  assign new_n4981_ = \i[1871]  & (\i[1870]  | \i[1869] );
  assign new_n4982_ = new_n4979_ & (\i[2765]  | \i[2766]  | \i[2767] ) & (\i[2402]  | \i[2403] );
  assign new_n4983_ = \i[1031]  & \i[1030]  & \i[1028]  & \i[1029] ;
  assign new_n4984_ = new_n4972_ & (new_n4987_ ? ~new_n4699_ : (new_n4986_ ? \i[2411]  : ~new_n4985_));
  assign new_n4985_ = ~\i[2311]  & ~\i[2310]  & ~\i[2308]  & ~\i[2309] ;
  assign new_n4986_ = ~\i[2391]  & (~\i[2390]  | ~\i[2389] );
  assign new_n4987_ = \i[1530]  & \i[1531] ;
  assign new_n4988_ = (new_n4998_ & (\i[1379]  ? ~new_n4995_ : ~new_n4989_)) | (~new_n4992_ & ~new_n4997_ & ~new_n4998_);
  assign new_n4989_ = ~new_n4991_ & (\i[878]  | \i[879]  | (new_n4968_ ? ~new_n4990_ : ~new_n3320_));
  assign new_n4990_ = new_n3438_ & ~\i[2048]  & ~\i[2049] ;
  assign new_n4991_ = ~\i[639]  & (\i[878]  | \i[879] ) & (~\i[638]  | (~\i[636]  & ~\i[637] ));
  assign new_n4992_ = new_n4993_ & (~\i[2203]  | (~\i[2202]  & (~\i[2201]  | ~\i[2200] )));
  assign new_n4993_ = ~new_n4066_ & new_n4994_ & \i[943]  & (\i[942]  | (\i[940]  & \i[941] ));
  assign new_n4994_ = \i[2191]  & \i[2189]  & \i[2190] ;
  assign new_n4995_ = new_n4996_ & (~\i[1044]  | ~\i[1045]  | ~\i[1046] );
  assign new_n4996_ = ~\i[1047]  & ((\i[624]  & \i[625] ) | \i[627]  | \i[626] );
  assign new_n4997_ = ~new_n3321_ & new_n4066_ & ((~\i[1618]  & ~\i[1619] ) | new_n4817_ | ~new_n3395_);
  assign new_n4998_ = ~\i[1275]  & (~\i[1273]  | ~\i[1274]  | ~\i[1272] );
  assign new_n4999_ = ~new_n3479_ & ~new_n4850_ & ~new_n4847_ & new_n4848_ & (\i[2753]  | ~new_n3849_);
  assign new_n5000_ = new_n5001_ ? (new_n5057_ ^ new_n4999_) : (~new_n5057_ ^ new_n4999_);
  assign new_n5001_ = new_n5002_ ? (~new_n5026_ ^ new_n5043_) : (new_n5026_ ^ new_n5043_);
  assign new_n5002_ = new_n3520_ ? (new_n3670_ ? ~new_n5003_ : ~new_n5009_) : new_n5015_;
  assign new_n5003_ = (new_n5004_ | ~new_n5008_) & (~new_n4334_ | ~new_n5006_ | new_n5008_);
  assign new_n5004_ = (\i[1711]  & (\i[1708]  | \i[1709]  | \i[1710] )) ? ~new_n4087_ : ~new_n5005_;
  assign new_n5005_ = \i[1951]  & \i[1950]  & \i[1948]  & \i[1949] ;
  assign new_n5006_ = new_n5007_ & ~\i[1184]  & ~\i[1185] ;
  assign new_n5007_ = ~\i[1186]  & ~\i[1187] ;
  assign new_n5008_ = \i[1735]  & (\i[1734]  | (\i[1733]  & \i[1732] ));
  assign new_n5009_ = new_n3602_ ? ((new_n5013_ | ~new_n5014_) & (new_n4942_ | ~\i[1499]  | new_n5014_)) : ~new_n5010_;
  assign new_n5010_ = (new_n5011_ | new_n5012_) & (~\i[2038]  | ~\i[2039]  | ~new_n5012_);
  assign new_n5011_ = \i[2639]  & (\i[2638]  | \i[2637] );
  assign new_n5012_ = ~\i[494]  & ~\i[495]  & (~\i[493]  | ~\i[492] );
  assign new_n5013_ = \i[1183]  & (\i[1182]  | (\i[1181]  & \i[1180] ));
  assign new_n5014_ = ~\i[1295]  & ~\i[1293]  & ~\i[1294] ;
  assign new_n5015_ = ~new_n5020_ & (~new_n5016_ | (new_n5017_ & (new_n5024_ ? ~new_n4207_ : ~new_n5025_)));
  assign new_n5016_ = ~new_n5019_ & (new_n5017_ | (new_n3666_ & ~new_n5018_) | (\i[1762]  & \i[1763]  & new_n5018_));
  assign new_n5017_ = ~\i[1987]  & ~\i[1986]  & ~\i[1984]  & ~\i[1985] ;
  assign new_n5018_ = \i[2055]  & \i[2053]  & \i[2054] ;
  assign new_n5019_ = ~\i[2547]  & ~\i[2545]  & ~\i[2546] ;
  assign new_n5020_ = ~new_n5023_ & new_n5019_ & (new_n5021_ ? ~new_n4232_ : new_n5022_);
  assign new_n5021_ = ~\i[1771]  & (~\i[1770]  | ~\i[1769] );
  assign new_n5022_ = ~\i[1178]  & ~\i[1179]  & (~\i[1177]  | ~\i[1176] );
  assign new_n5023_ = ~\i[2215]  & ~\i[2213]  & ~\i[2214] ;
  assign new_n5024_ = ~\i[1150]  & ~\i[1151]  & (~\i[1149]  | ~\i[1148] );
  assign new_n5025_ = ~\i[2399]  & ~\i[2398]  & ~\i[2396]  & ~\i[2397] ;
  assign new_n5026_ = new_n3423_ ? ((~new_n5037_ & ~new_n5041_) | (~new_n5040_ & new_n5042_ & new_n5041_)) : new_n5027_;
  assign new_n5027_ = new_n3468_ ? ((new_n5033_ | new_n3367_) & (new_n5035_ | ~new_n5036_ | ~new_n3367_)) : new_n5028_;
  assign new_n5028_ = new_n5031_ ? (new_n4067_ ? ~new_n4851_ : new_n5032_) : new_n5029_;
  assign new_n5029_ = new_n4783_ ? new_n5030_ : ~new_n4769_;
  assign new_n5030_ = \i[2387]  & \i[2386]  & \i[2384]  & \i[2385] ;
  assign new_n5031_ = ~\i[1283]  & (~\i[1281]  | ~\i[1282]  | ~\i[1280] );
  assign new_n5032_ = ~\i[2431]  & ~\i[2430]  & ~\i[2428]  & ~\i[2429] ;
  assign new_n5033_ = ~\i[2546]  & ~\i[2547]  & new_n5034_ & (~\i[2545]  | ~\i[2544] );
  assign new_n5034_ = ~\i[2099]  & ~\i[2098]  & ~\i[2096]  & ~\i[2097] ;
  assign new_n5035_ = \i[2066]  & \i[2067]  & (\i[2065]  | \i[2064] );
  assign new_n5036_ = ~\i[1935]  & ~\i[1934]  & ~\i[1932]  & ~\i[1933] ;
  assign new_n5037_ = (~new_n3269_ | ~new_n5038_ | ~new_n4030_) & (new_n3526_ | \i[1714]  | \i[1715]  | new_n4030_);
  assign new_n5038_ = new_n5039_ & (~\i[1601]  | ~\i[1600] );
  assign new_n5039_ = ~\i[1602]  & ~\i[1603] ;
  assign new_n5040_ = new_n4667_ ? (~\i[1031]  & (~\i[1028]  | ~\i[1029]  | ~\i[1030] )) : new_n4723_;
  assign new_n5041_ = new_n4851_ & ~\i[1380]  & ~\i[1381] ;
  assign new_n5042_ = ~\i[1479]  & ~\i[1477]  & ~\i[1478] ;
  assign new_n5043_ = new_n4437_ ? new_n5046_ : (new_n5056_ ? ~new_n5055_ : ~new_n5044_);
  assign new_n5044_ = (~new_n5045_ | new_n3538_) & (~\i[2553]  | ~\i[2554]  | ~\i[2555] ) & (new_n4100_ | ~new_n3538_);
  assign new_n5045_ = ~\i[2343]  & ~\i[2342]  & ~\i[2340]  & ~\i[2341] ;
  assign new_n5046_ = new_n5052_ ? new_n5047_ : ((~new_n5050_ | ~new_n5053_) & (new_n3238_ | ~new_n5054_ | new_n5053_));
  assign new_n5047_ = (new_n5034_ | ~\i[2198]  | ~\i[2199]  | new_n4872_) & (~new_n4872_ | (~new_n5049_ & ~new_n5048_));
  assign new_n5048_ = ~\i[2747]  & ~\i[2746]  & ~\i[2744]  & ~\i[2745] ;
  assign new_n5049_ = ~\i[1831]  & (~\i[1830]  | (~\i[1829]  & ~\i[1828] ));
  assign new_n5050_ = new_n5051_ & (\i[1435]  | \i[1434] );
  assign new_n5051_ = ~\i[2218]  & ~\i[2219]  & (~\i[2217]  | ~\i[2216] );
  assign new_n5052_ = ~\i[1282]  & ~\i[1283] ;
  assign new_n5053_ = ~\i[1779]  & ~\i[1777]  & ~\i[1778] ;
  assign new_n5054_ = ~\i[1311]  & ~\i[1309]  & ~\i[1310] ;
  assign new_n5055_ = ~\i[1755]  & new_n4256_ & new_n4418_ & (~\i[1754]  | (~\i[1752]  & ~\i[1753] ));
  assign new_n5056_ = ~\i[1607]  & (~\i[1605]  | ~\i[1606]  | ~\i[1604] );
  assign new_n5057_ = new_n5058_ ? (~new_n5074_ ^ new_n5090_) : (new_n5074_ ^ new_n5090_);
  assign new_n5058_ = (new_n5059_ | ~new_n5067_) & (new_n5069_ | new_n5071_ | new_n5073_ | ~new_n3462_ | new_n5067_);
  assign new_n5059_ = new_n4278_ ? new_n5060_ : ((new_n5064_ | ~new_n4437_) & (new_n4077_ | ~new_n5066_ | new_n4437_));
  assign new_n5060_ = (~new_n3392_ | new_n5061_ | new_n3438_) & (~new_n3438_ | (new_n5032_ ? ~new_n5062_ : new_n5063_));
  assign new_n5061_ = ~\i[1483]  & (~\i[1482]  | (~\i[1481]  & ~\i[1480] ));
  assign new_n5062_ = ~\i[2211]  & ~\i[2210]  & ~\i[2208]  & ~\i[2209] ;
  assign new_n5063_ = ~\i[2094]  & ~\i[2095]  & (~\i[2093]  | ~\i[2092] );
  assign new_n5064_ = (~\i[2526]  & ~\i[2527]  & new_n5065_) | (~new_n5065_ & (\i[1601]  | ~new_n5039_));
  assign new_n5065_ = ~\i[1039]  & ~\i[1038]  & ~\i[1036]  & ~\i[1037] ;
  assign new_n5066_ = new_n4808_ & new_n5039_;
  assign new_n5067_ = new_n5068_ & ~\i[1392]  & ~\i[1393] ;
  assign new_n5068_ = ~\i[1394]  & ~\i[1395] ;
  assign new_n5069_ = ~new_n5070_ & (\i[2529]  | ~new_n3510_);
  assign new_n5070_ = ~\i[1982]  & ~\i[1983]  & (~\i[1981]  | ~\i[1980] );
  assign new_n5071_ = \i[1857]  & \i[1856]  & new_n5072_ & ~\i[2531]  & ~\i[2529]  & ~\i[2530] ;
  assign new_n5072_ = \i[1858]  & \i[1859] ;
  assign new_n5073_ = ~\i[2323]  & ~\i[2322]  & ~\i[2320]  & ~\i[2321] ;
  assign new_n5074_ = new_n5088_ ? ((new_n5081_ | new_n5087_) & (~new_n5085_ | ~new_n5089_ | ~new_n5087_)) : new_n5075_;
  assign new_n5075_ = new_n4678_ ? (~new_n5080_ | (~new_n4132_ & \i[1478]  & \i[1479] )) : new_n5076_;
  assign new_n5076_ = (~new_n5079_ | ~new_n3394_ | new_n5077_) & (~new_n5077_ | (new_n4075_ ? new_n3645_ : ~new_n4661_));
  assign new_n5077_ = new_n5078_ & ~\i[2076]  & ~\i[2077] ;
  assign new_n5078_ = ~\i[2078]  & ~\i[2079] ;
  assign new_n5079_ = ~\i[2387]  & ~\i[2386]  & ~\i[2384]  & ~\i[2385] ;
  assign new_n5080_ = ~\i[1771]  & ~\i[1770]  & ~\i[1768]  & ~\i[1769] ;
  assign new_n5081_ = (~new_n5083_ | new_n4879_ | ~new_n5082_) & (new_n5082_ | (new_n5084_ ? ~new_n3491_ : ~\i[2115] ));
  assign new_n5082_ = new_n4323_ & ~\i[1384]  & ~\i[1385] ;
  assign new_n5083_ = new_n4657_ & ~\i[1948]  & ~\i[1949] ;
  assign new_n5084_ = \i[2551]  & (\i[2550]  | \i[2549] );
  assign new_n5085_ = new_n5086_ & (\i[1895]  | (\i[1894]  & (\i[1893]  | \i[1892] )));
  assign new_n5086_ = ~\i[2259]  & ~\i[2258]  & ~\i[2256]  & ~\i[2257] ;
  assign new_n5087_ = ~\i[499]  & ~\i[498]  & ~\i[496]  & ~\i[497] ;
  assign new_n5088_ = ~\i[2335]  & ~\i[2334]  & ~\i[2332]  & ~\i[2333] ;
  assign new_n5089_ = ~\i[2114]  & ~\i[2115]  & (~\i[2113]  | ~\i[2112] );
  assign new_n5090_ = new_n4056_ ? new_n5096_ : ((new_n5091_ | ~new_n5100_) & (new_n5095_ | ~new_n5102_ | new_n5100_));
  assign new_n5091_ = (~\i[1922]  | ~\i[1923]  | ~new_n5093_) & (new_n5092_ | new_n5093_ | (~new_n5094_ & ~new_n3384_));
  assign new_n5092_ = new_n3384_ & ~\i[1767]  & ~\i[1765]  & ~\i[1766] ;
  assign new_n5093_ = ~\i[2227]  & ~\i[2225]  & ~\i[2226] ;
  assign new_n5094_ = ~\i[1883]  & ~\i[1882]  & ~\i[1880]  & ~\i[1881] ;
  assign new_n5095_ = (~\i[1710]  & ~\i[1711] ) ? ~new_n4469_ : ~new_n4087_;
  assign new_n5096_ = ~new_n5097_ & (~new_n3223_ | (new_n3778_ & new_n5099_) | (~new_n3396_ & ~new_n5098_ & ~new_n5099_));
  assign new_n5097_ = new_n3368_ & new_n5087_ & ~\i[1375]  & ~\i[1374]  & ~new_n3223_ & ~\i[1373] ;
  assign new_n5098_ = ~\i[1375]  & ~\i[1374]  & ~\i[1372]  & ~\i[1373] ;
  assign new_n5099_ = ~\i[2047]  & (~\i[2046]  | ~\i[2045] );
  assign new_n5100_ = new_n5101_ & ~\i[2044]  & ~\i[2045] ;
  assign new_n5101_ = ~\i[2046]  & ~\i[2047] ;
  assign new_n5102_ = ~\i[1171]  & ~\i[1170]  & ~\i[1168]  & ~\i[1169] ;
  assign new_n5103_ = (new_n5104_ | \i[1919] ) & (new_n4682_ | new_n5110_ | ~\i[1919] );
  assign new_n5104_ = ~new_n5105_ & (new_n5109_ | new_n4742_ | \i[1157]  | \i[1158]  | \i[1159] );
  assign new_n5105_ = new_n4742_ & (new_n5108_ ? (~new_n4764_ | ~new_n4657_) : ~new_n5106_);
  assign new_n5106_ = \i[951]  & new_n5107_ & ~\i[1374]  & ~\i[1375] ;
  assign new_n5107_ = \i[949]  & \i[950]  & (~\i[1373]  | ~\i[1372] );
  assign new_n5108_ = \i[2279]  & (\i[2277]  | \i[2278]  | \i[2276] );
  assign new_n5109_ = ~new_n4788_ & ~\i[1511]  & (~\i[1510]  | ~\i[1509]  | ~\i[1508] );
  assign new_n5110_ = ~\i[2095]  & (~\i[2094]  | (~\i[2093]  & ~\i[2092] ));
  assign new_n5111_ = new_n4007_ ? new_n5112_ : ((new_n5121_ | new_n5119_ | ~new_n5129_) & (new_n5123_ | new_n5129_));
  assign new_n5112_ = ~new_n5113_ & (~new_n3383_ | ((new_n5117_ | new_n5094_) & (~new_n3281_ | ~new_n3652_ | ~new_n5094_)));
  assign new_n5113_ = ~new_n3383_ & ~new_n5114_ & (\i[1665]  | \i[1666]  | \i[1667]  | ~new_n5116_);
  assign new_n5114_ = new_n5065_ & new_n5115_ & (\i[1555]  | \i[1554] );
  assign new_n5115_ = \i[1939]  & (\i[1938]  | (\i[1937]  & \i[1936] ));
  assign new_n5116_ = ~\i[1554]  & ~\i[1555]  & \i[1175]  & (\i[1174]  | \i[1173] );
  assign new_n5117_ = new_n4018_ ? new_n5118_ : (~\i[939]  | (~\i[937]  & ~\i[938] ));
  assign new_n5118_ = \i[2095]  & (\i[2094]  | \i[2093] );
  assign new_n5119_ = ~new_n4734_ & ((\i[2175]  & new_n5120_) | (~\i[2627]  & ~new_n5120_ & (~\i[2626]  | ~\i[2625] )));
  assign new_n5120_ = ~\i[2095]  & (~\i[2093]  | ~\i[2094]  | ~\i[2092] );
  assign new_n5121_ = ~new_n5122_ & new_n4734_ & (\i[1031]  | (\i[1029]  & \i[1030] ));
  assign new_n5122_ = ~\i[1827]  & (~\i[1826]  | (~\i[1825]  & ~\i[1824] ));
  assign new_n5123_ = new_n5128_ ? ((new_n5127_ & ~new_n5126_) | (new_n3614_ & \i[1843]  & new_n5126_)) : new_n5124_;
  assign new_n5124_ = (~new_n5125_ & (~\i[2617]  | ~\i[2618]  | ~\i[2619] )) | (~\i[2616]  & (~new_n5125_ | (~\i[2617]  & ~\i[2618]  & ~\i[2619] )));
  assign new_n5125_ = \i[1507]  & \i[1505]  & \i[1506] ;
  assign new_n5126_ = ~\i[1611]  & (~\i[1609]  | ~\i[1610]  | ~\i[1608] );
  assign new_n5127_ = ~\i[2150]  & ~\i[2151]  & (~\i[2149]  | ~\i[2148] );
  assign new_n5128_ = ~\i[1715]  & ~\i[1714]  & ~\i[1712]  & ~\i[1713] ;
  assign new_n5129_ = ~\i[1378]  & ~\i[1379]  & (~\i[1377]  | ~\i[1376] );
  assign new_n5130_ = (new_n5131_ & ~new_n4389_) | (~new_n5144_ & new_n4389_ & (~new_n5036_ | new_n5140_));
  assign new_n5131_ = new_n4235_ ? (new_n5139_ ? new_n5135_ : new_n5137_) : new_n5132_;
  assign new_n5132_ = (~new_n5053_ | ~new_n5133_ | ~new_n4731_) & (new_n5134_ | ~new_n3284_ | new_n4731_);
  assign new_n5133_ = ~\i[1399]  & ~\i[1397]  & ~\i[1398] ;
  assign new_n5134_ = ~\i[1875]  & ~\i[1874]  & ~\i[1872]  & ~\i[1873] ;
  assign new_n5135_ = new_n3299_ ? ~new_n5136_ : \i[1483] ;
  assign new_n5136_ = new_n4755_ & ~\i[2608]  & ~\i[2609] ;
  assign new_n5137_ = (~new_n4757_ | new_n5138_) & (\i[510]  | \i[511]  | ~new_n5138_ | (\i[509]  & \i[508] ));
  assign new_n5138_ = new_n3414_ & (~\i[1605]  | ~\i[1604] );
  assign new_n5139_ = ~\i[1383]  & (~\i[1381]  | ~\i[1382]  | ~\i[1380] );
  assign new_n5140_ = new_n4317_ ? (new_n5141_ | (~\i[586]  & ~\i[587]  & new_n4536_)) : new_n5142_;
  assign new_n5141_ = ~new_n4536_ & (\i[2533]  | ~new_n4735_);
  assign new_n5142_ = new_n5143_ & (~\i[1815]  | ~\i[1814] );
  assign new_n5143_ = ~\i[1670]  & ~\i[1671]  & (~\i[1669]  | ~\i[1668] );
  assign new_n5144_ = ~new_n4437_ & ~new_n5036_ & ~\i[499]  & (\i[2375]  | \i[2374]  | \i[2373] );
  assign new_n5145_ = new_n4659_ ? new_n5153_ : (~new_n5146_ & (~new_n5159_ | ~new_n5133_ | ~\i[2439] ));
  assign new_n5146_ = new_n5152_ & (new_n5147_ | (~new_n4080_ & ~new_n5150_ & ~new_n5151_));
  assign new_n5147_ = new_n4080_ & (new_n5148_ ? ~new_n5149_ : new_n3327_);
  assign new_n5148_ = new_n3339_ & ~\i[2052]  & ~\i[2053] ;
  assign new_n5149_ = \i[1934]  & \i[1935]  & (\i[1933]  | \i[1932] );
  assign new_n5150_ = ~\i[2331]  & ~\i[2330]  & ~\i[2328]  & ~\i[2329] ;
  assign new_n5151_ = ~\i[1162]  & ~\i[1163]  & (~\i[1161]  | ~\i[1160] );
  assign new_n5152_ = ~\i[2635]  & ~\i[2633]  & ~\i[2634] ;
  assign new_n5153_ = ~new_n5154_ & (~new_n5157_ | (\i[2631]  & (new_n5158_ | ~new_n4214_)));
  assign new_n5154_ = new_n3447_ & ((new_n3845_ & new_n3254_ & ~new_n5155_) | (~new_n4469_ & ~new_n5156_ & new_n5155_));
  assign new_n5155_ = new_n3659_ & ~\i[612]  & ~\i[613] ;
  assign new_n5156_ = ~\i[1046]  & ~\i[1047]  & (~\i[1045]  | ~\i[1044] );
  assign new_n5157_ = ~new_n3447_ & (\i[2631]  | (new_n3494_ & new_n4072_));
  assign new_n5158_ = \i[2059]  & (\i[2058]  | \i[2057] );
  assign new_n5159_ = ~\i[2119]  & ~\i[2118]  & ~new_n5152_ & ~\i[2117] ;
  assign \o[15]  = new_n5161_ ^ new_n5294_;
  assign new_n5161_ = new_n5162_ ? (~new_n5292_ ^ new_n5293_) : (new_n5292_ ^ new_n5293_);
  assign new_n5162_ = new_n5163_ ? (~new_n5277_ ^ new_n5278_) : (new_n5277_ ^ new_n5278_);
  assign new_n5163_ = new_n5164_ ? (~new_n5247_ ^ new_n5248_) : (new_n5247_ ^ new_n5248_);
  assign new_n5164_ = new_n5165_ ? (~new_n5216_ ^ new_n5246_) : (new_n5216_ ^ new_n5246_);
  assign new_n5165_ = new_n5166_ ? (~new_n5190_ ^ new_n5191_) : (new_n5190_ ^ new_n5191_);
  assign new_n5166_ = new_n5167_ ^ new_n5181_;
  assign new_n5167_ = new_n4056_ ? ((~new_n5178_ & ~new_n5180_ & new_n3223_) | (new_n5174_ & ~new_n3223_)) : new_n5168_;
  assign new_n5168_ = new_n5100_ ? (new_n5093_ ? new_n5172_ : ~new_n5092_) : new_n5169_;
  assign new_n5169_ = new_n5102_ ? new_n5170_ : (new_n4939_ ? new_n5171_ : ~new_n5080_);
  assign new_n5170_ = (~\i[1710]  & ~\i[1711] ) ? new_n4469_ : ~new_n4087_;
  assign new_n5171_ = ~\i[2007]  & ~\i[2006]  & ~\i[2004]  & ~\i[2005] ;
  assign new_n5172_ = (\i[1922]  & \i[1923] ) ? ~new_n5173_ : (~\i[1779]  | (~\i[1778]  & ~\i[1777] ));
  assign new_n5173_ = \i[1746]  & \i[1747]  & (\i[1745]  | \i[1744] );
  assign new_n5174_ = new_n3368_ ? new_n5175_ : (new_n5073_ ? new_n5177_ : new_n4206_);
  assign new_n5175_ = ~new_n5176_ & (\i[1373]  | \i[1374]  | \i[1375] );
  assign new_n5176_ = ~\i[1599]  & ~\i[1597]  & ~\i[1598] ;
  assign new_n5177_ = ~\i[1995]  & ~\i[1994]  & ~\i[1992]  & ~\i[1993] ;
  assign new_n5178_ = new_n5099_ & (~new_n5179_ | new_n3778_) & (\i[2005]  | \i[2006]  | \i[2007]  | ~new_n3778_);
  assign new_n5179_ = ~\i[2659]  & ~\i[2658]  & ~\i[2656]  & ~\i[2657] ;
  assign new_n5180_ = new_n5098_ & ~\i[1399]  & ~new_n5099_ & ~\i[1398] ;
  assign new_n5181_ = new_n5088_ ? new_n5187_ : new_n5182_;
  assign new_n5182_ = new_n4678_ ? new_n5185_ : ((~new_n5183_ & ~new_n5077_) | (~new_n3645_ & new_n4075_ & new_n5077_));
  assign new_n5183_ = new_n5079_ ? ~new_n3394_ : new_n5184_;
  assign new_n5184_ = \i[1770]  & \i[1771]  & (\i[1769]  | \i[1768] );
  assign new_n5185_ = (~\i[1478]  | ~\i[1479]  | ~new_n5080_) & (new_n5186_ | ~new_n4219_ | new_n5080_);
  assign new_n5186_ = \i[1954]  & \i[1955]  & (\i[1953]  | \i[1952] );
  assign new_n5187_ = ~new_n5188_ & (~new_n5087_ | (new_n5189_ & ~new_n5089_) | (~new_n5086_ & \i[1959]  & new_n5089_));
  assign new_n5188_ = ~new_n5087_ & (~new_n5129_ | new_n5083_ | ~new_n5082_) & (new_n5084_ | ~\i[2115]  | new_n5082_);
  assign new_n5189_ = ~\i[2839]  & ~\i[2838]  & ~\i[2837]  & ~\i[2836]  & ~\i[1486]  & ~\i[1487] ;
  assign new_n5190_ = (~new_n5074_ & ~new_n5090_) | (~new_n5058_ & (~new_n5074_ | ~new_n5090_));
  assign new_n5191_ = new_n5192_ ? (~new_n5201_ ^ new_n5207_) : (new_n5201_ ^ new_n5207_);
  assign new_n5192_ = (new_n5193_ & new_n4389_) | (~new_n5199_ & ~new_n4389_ & (new_n5139_ | ~new_n5198_));
  assign new_n5193_ = new_n5036_ ? ((~new_n5141_ | ~new_n4317_) & (new_n5143_ | ~new_n5197_ | new_n4317_)) : new_n5194_;
  assign new_n5194_ = (new_n5196_ | ~\i[499]  | new_n4437_) & (~new_n4437_ | (new_n3511_ ? ~new_n5195_ : new_n4677_));
  assign new_n5195_ = ~\i[1371]  & (~\i[1370]  | ~\i[1369] );
  assign new_n5196_ = ~\i[1979]  & (~\i[1978]  | (~\i[1977]  & ~\i[1976] ));
  assign new_n5197_ = ~\i[831]  & (~\i[830]  | ~\i[829] );
  assign new_n5198_ = new_n5138_ & new_n4235_ & ((\i[508]  & \i[509] ) | \i[511]  | \i[510] );
  assign new_n5199_ = ~new_n4235_ & ((~new_n5053_ & ~\i[1487]  & new_n4731_) | (new_n5134_ & new_n5200_ & ~new_n4731_));
  assign new_n5200_ = ~\i[1487]  & ~\i[1486]  & ~\i[1484]  & ~\i[1485] ;
  assign new_n5201_ = (~new_n5159_ & ~new_n5202_ & ~new_n4659_) | (~new_n5204_ & new_n4659_ & (new_n5206_ | ~new_n5157_));
  assign new_n5202_ = new_n5152_ & (new_n5147_ | (~new_n5203_ & ~new_n4080_));
  assign new_n5203_ = (new_n5151_ | new_n5150_) & (\i[1896]  | \i[1897]  | \i[1898]  | \i[1899]  | ~new_n5150_);
  assign new_n5204_ = new_n3447_ & (new_n5155_ ? ~new_n5205_ : (new_n3254_ ? ~new_n3845_ : ~new_n4851_));
  assign new_n5205_ = new_n4469_ ? (\i[2043]  & (\i[2040]  | \i[2041]  | \i[2042] )) : new_n5156_;
  assign new_n5206_ = \i[2631]  & new_n5158_ & ~\i[1975]  & ~\i[1974]  & ~\i[1972]  & ~\i[1973] ;
  assign new_n5207_ = (new_n5211_ | new_n5208_ | new_n5067_) & (~new_n5067_ | (new_n4278_ ? new_n5214_ : new_n5213_));
  assign new_n5208_ = new_n3462_ & (new_n5073_ ? (new_n5209_ ? ~new_n4823_ : ~new_n5210_) : ~new_n5071_);
  assign new_n5209_ = ~\i[1883]  & (~\i[1882]  | (~\i[1881]  & ~\i[1880] ));
  assign new_n5210_ = ~\i[2419]  & (~\i[2418]  | (~\i[2417]  & ~\i[2416] ));
  assign new_n5211_ = ~new_n3462_ & new_n5212_ & (~\i[2667]  | (~\i[2664]  & ~\i[2665]  & ~\i[2666] ));
  assign new_n5212_ = (~\i[1895]  & (~\i[1893]  | ~\i[1894] ) & (~\i[1822]  | ~\i[1823] )) | (~new_n3511_ & \i[1822]  & \i[1823] );
  assign new_n5213_ = (~new_n5066_ | ~new_n4077_ | new_n4437_) & (\i[2526]  | \i[2527]  | ~new_n5065_ | ~new_n4437_);
  assign new_n5214_ = (~new_n3438_ | (new_n5032_ ? new_n5062_ : ~new_n5063_)) & (~new_n5061_ | ~new_n5215_ | new_n3438_);
  assign new_n5215_ = ~\i[2738]  & ~\i[2739]  & (~\i[2737]  | ~\i[2736] );
  assign new_n5216_ = new_n5217_ ? (new_n5244_ ^ new_n5245_) : (~new_n5244_ ^ new_n5245_);
  assign new_n5217_ = new_n5218_ ? (new_n5225_ ^ new_n5234_) : (~new_n5225_ ^ new_n5234_);
  assign new_n5218_ = new_n3736_ ? ((new_n5222_ | new_n4784_ | ~new_n3697_) & (new_n5224_ | new_n3697_)) : new_n5219_;
  assign new_n5219_ = (new_n5221_ | new_n5220_ | new_n4788_) & (new_n3585_ | new_n4789_ | new_n4790_ | ~new_n4788_);
  assign new_n5220_ = new_n4190_ & (~new_n4794_ | ~\i[2197]  | ~\i[2198]  | ~\i[2199] );
  assign new_n5221_ = ~new_n4190_ & (~new_n4792_ | (new_n4705_ & \i[2409] ));
  assign new_n5222_ = (~new_n5223_ | new_n4785_) & (\i[1442]  | \i[1443]  | ~new_n4785_);
  assign new_n5223_ = ~\i[959]  & (~\i[958]  | (~\i[957]  & ~\i[956] ));
  assign new_n5224_ = (new_n4779_ | ~new_n4780_ | ~new_n3615_) & (~new_n3365_ | new_n3615_ | (~\i[835]  & ~\i[834] ));
  assign new_n5225_ = new_n3423_ ? new_n5226_ : ((~new_n5232_ & ~new_n3468_) | (~new_n3367_ & new_n5233_ & new_n3468_));
  assign new_n5226_ = ~new_n5227_ & (new_n5041_ | (~new_n5229_ & ~new_n4030_) | (~new_n5038_ & \i[2671]  & new_n4030_));
  assign new_n5227_ = new_n5041_ & (new_n5042_ ? ~new_n4667_ : (new_n5228_ | ~new_n4864_));
  assign new_n5228_ = \i[1375]  & (\i[1373]  | \i[1374]  | \i[1372] );
  assign new_n5229_ = (new_n5231_ & (new_n3526_ | \i[1714]  | \i[1715] )) | (~\i[1714]  & ~\i[1715]  & new_n5230_ & ~new_n3526_);
  assign new_n5230_ = ~\i[2166]  & ~\i[2167] ;
  assign new_n5231_ = ~\i[1619]  & (~\i[1618]  | (~\i[1617]  & ~\i[1616] ));
  assign new_n5232_ = (new_n4783_ | ~new_n4769_ | new_n5031_) & (~new_n5031_ | (new_n4067_ ? ~new_n4851_ : new_n5032_));
  assign new_n5233_ = (~new_n5034_ & ~\i[2546]  & ~\i[2547]  & (~\i[2544]  | ~\i[2545] )) | (new_n4739_ & (\i[2546]  | \i[2547]  | (\i[2544]  & \i[2545] )));
  assign new_n5234_ = new_n4437_ ? new_n5235_ : (new_n5056_ ? new_n5239_ : ~new_n5243_);
  assign new_n5235_ = (new_n5236_ | new_n5052_) & (new_n4872_ | ~new_n5034_ | ~new_n5238_ | ~new_n5052_);
  assign new_n5236_ = (new_n5051_ | new_n5237_ | ~new_n5053_) & (~new_n3238_ | ~new_n5054_ | new_n5053_);
  assign new_n5237_ = ~\i[610]  & ~\i[611]  & (~\i[609]  | ~\i[608] );
  assign new_n5238_ = ~\i[1482]  & ~\i[1483]  & (~\i[1481]  | ~\i[1480] );
  assign new_n5239_ = (new_n4418_ | ~new_n5242_ | ~new_n4256_) & (new_n4256_ | (new_n4847_ ? new_n5240_ : ~new_n5241_));
  assign new_n5240_ = ~\i[1175]  & (~\i[1174]  | ~\i[1173] );
  assign new_n5241_ = \i[1362]  & \i[1363]  & (\i[1361]  | \i[1360] );
  assign new_n5242_ = ~\i[1611]  & (~\i[1610]  | (~\i[1609]  & ~\i[1608] ));
  assign new_n5243_ = \i[2555]  & \i[2554]  & ~new_n3638_ & \i[2553] ;
  assign new_n5244_ = (~new_n4943_ & ~new_n4969_) | (~new_n4925_ & (~new_n4943_ | ~new_n4969_));
  assign new_n5245_ = (~new_n5043_ & new_n5026_) | (new_n5002_ & (~new_n5043_ | new_n5026_));
  assign new_n5246_ = (~new_n5057_ & new_n4999_) | (~new_n5001_ & (~new_n5057_ | new_n4999_));
  assign new_n5247_ = (~new_n5000_ & ~new_n5103_) | (~new_n4923_ & (~new_n5000_ | ~new_n5103_));
  assign new_n5248_ = new_n5249_ ? (new_n5250_ ^ new_n5276_) : (~new_n5250_ ^ new_n5276_);
  assign new_n5249_ = (~new_n4852_ & ~new_n4706_) | (~new_n4798_ & (~new_n4852_ | ~new_n4706_));
  assign new_n5250_ = new_n5251_ ? (new_n5252_ ^ new_n5271_) : (~new_n5252_ ^ new_n5271_);
  assign new_n5251_ = (~new_n4825_ & ~new_n4838_) | (~new_n4799_ & (~new_n4825_ | ~new_n4838_));
  assign new_n5252_ = new_n5253_ ? (~new_n5259_ ^ new_n5267_) : (new_n5259_ ^ new_n5267_);
  assign new_n5253_ = new_n3520_ ? new_n5254_ : new_n5257_;
  assign new_n5254_ = (new_n4334_ | new_n5008_ | new_n5256_ | ~new_n3670_) & (new_n5255_ | new_n3670_);
  assign new_n5255_ = (new_n5010_ | new_n3602_) & (~new_n5013_ | ~new_n5014_ | ~new_n3602_);
  assign new_n5256_ = ~\i[2191]  & ~\i[2190]  & ~\i[2188]  & ~\i[2189] ;
  assign new_n5257_ = (~new_n5024_ | ~new_n5017_ | ~new_n4207_ | new_n5019_) & (~new_n5023_ | new_n5258_ | ~new_n5019_);
  assign new_n5258_ = ~\i[2771]  & (~\i[2770]  | (~\i[2769]  & ~\i[2768] ));
  assign new_n5259_ = new_n4007_ ? (new_n3383_ ? new_n5265_ : ~new_n5114_) : new_n5260_;
  assign new_n5260_ = new_n5129_ ? (~new_n5264_ & (new_n4734_ | ~new_n5120_ | ~\i[2175] )) : new_n5261_;
  assign new_n5261_ = (~new_n5126_ | ~new_n3614_ | ~\i[1843]  | ~new_n5128_) & (~new_n5125_ | ~new_n5262_ | new_n5128_);
  assign new_n5262_ = new_n5263_ & ~\i[2616]  & ~\i[2617] ;
  assign new_n5263_ = ~\i[2618]  & ~\i[2619] ;
  assign new_n5264_ = new_n5122_ & new_n4734_ & (\i[2871]  | (\i[2869]  & \i[2870] ));
  assign new_n5265_ = (new_n5266_ | ~new_n5094_) & (~new_n4018_ | ~new_n5118_ | new_n5094_);
  assign new_n5266_ = (new_n3652_ | ~new_n3281_) & (~\i[1539]  | new_n3281_ | (~\i[1538]  & (~\i[1536]  | ~\i[1537] )));
  assign new_n5267_ = ~new_n5268_ & (new_n4774_ | (~new_n5270_ & ~new_n3275_) | (new_n4754_ & new_n4756_ & new_n3275_));
  assign new_n5268_ = ~new_n5269_ & new_n4774_ & (new_n4219_ | new_n4771_ | new_n5030_ | ~new_n4772_);
  assign new_n5269_ = ~\i[1635]  & new_n4219_ & new_n4767_ & new_n4769_ & (~\i[1634]  | ~\i[1633] );
  assign new_n5270_ = (~new_n4763_ | new_n4764_) & (new_n4676_ | new_n4760_ | ~new_n4764_);
  assign new_n5271_ = new_n5272_ ? (new_n5274_ ^ new_n5275_) : (~new_n5274_ ^ new_n5275_);
  assign new_n5272_ = (~new_n5273_ | ~new_n4820_) & (new_n4985_ | new_n4986_ | new_n4987_ | ~new_n4972_ | new_n4820_);
  assign new_n5273_ = ~\i[1627]  & new_n4983_ & new_n3905_ & (~\i[1626]  | ~\i[1625] );
  assign new_n5274_ = new_n4704_ & new_n4913_ & new_n4912_ & ~new_n3728_ & ~new_n4918_;
  assign new_n5275_ = new_n4957_ & new_n3275_ & ~new_n4968_ & ~new_n4956_ & ~new_n4958_;
  assign new_n5276_ = (~new_n4988_ & new_n4999_) | (~new_n4924_ & (~new_n4988_ | new_n4999_));
  assign new_n5277_ = (~new_n4922_ & ~new_n5111_) | (~new_n4796_ & (~new_n4922_ | ~new_n5111_));
  assign new_n5278_ = new_n5279_ ? (new_n5280_ ^ new_n5291_) : (~new_n5280_ ^ new_n5291_);
  assign new_n5279_ = (~new_n4728_ & ~new_n4743_) | (~new_n4645_ & (~new_n4728_ | ~new_n4743_));
  assign new_n5280_ = new_n5281_ ? (new_n5282_ ^ new_n5290_) : (~new_n5282_ ^ new_n5290_);
  assign new_n5281_ = (~new_n4706_ & ~new_n4712_) | (~new_n4646_ & (~new_n4706_ | ~new_n4712_));
  assign new_n5282_ = new_n5283_ ? (new_n5284_ ^ new_n5285_) : (~new_n5284_ ^ new_n5285_);
  assign new_n5283_ = (~new_n4669_ & ~new_n4686_) | (~new_n4647_ & (~new_n4669_ | ~new_n4686_));
  assign new_n5284_ = (~new_n4866_ & new_n4882_) | (~new_n4853_ & (~new_n4866_ | new_n4882_));
  assign new_n5285_ = ((\i[1487]  | \i[1519]  | ~new_n5288_ | ~new_n4837_) & (new_n5286_ ^ new_n5289_)) | (~\i[1487]  & ~\i[1519]  & new_n5288_ & new_n4837_ & (new_n5286_ ^ ~new_n5289_));
  assign new_n5286_ = ~new_n5287_ & (new_n4165_ | ~new_n3258_ | ~new_n3349_ | ~new_n4802_ | ~new_n4804_);
  assign new_n5287_ = new_n4814_ & new_n4821_ & ~new_n4813_ & ~new_n3258_ & ~new_n4078_;
  assign new_n5288_ = ~new_n3849_ & ~new_n4666_;
  assign new_n5289_ = ~new_n4682_ & ~\i[2095]  & \i[1919]  & (~\i[2094]  | (~\i[2092]  & ~\i[2093] ));
  assign new_n5290_ = ~new_n4726_ & ~new_n4719_ & ~\i[2087]  & new_n4718_ & (~\i[2086]  | ~\i[2085] );
  assign new_n5291_ = (~new_n4886_ & ~new_n4909_) | (~new_n4797_ & (~new_n4886_ | ~new_n4909_));
  assign new_n5292_ = (~new_n4795_ & ~new_n5130_) | (~new_n4643_ & (~new_n4795_ | ~new_n5130_));
  assign new_n5293_ = (~new_n4751_ & ~new_n4775_) | (~new_n4644_ & (~new_n4751_ | ~new_n4775_));
  assign new_n5294_ = ~new_n4642_ & ~new_n5145_;
  assign \o[16]  = ~new_n5296_ ^ new_n5297_;
  assign new_n5296_ = new_n5161_ & new_n5294_;
  assign new_n5297_ = new_n5298_ ^ new_n5299_;
  assign new_n5298_ = (new_n5292_ & new_n5293_) | (new_n5162_ & (new_n5292_ | new_n5293_));
  assign new_n5299_ = new_n5300_ ? (~new_n5301_ ^ new_n5335_) : (new_n5301_ ^ new_n5335_);
  assign new_n5300_ = (new_n5277_ & new_n5278_) | (new_n5163_ & (new_n5277_ | new_n5278_));
  assign new_n5301_ = new_n5302_ ? (new_n5303_ ^ new_n5327_) : (~new_n5303_ ^ new_n5327_);
  assign new_n5302_ = (new_n5247_ & new_n5248_) | (new_n5164_ & (new_n5247_ | new_n5248_));
  assign new_n5303_ = new_n5304_ ? (new_n5305_ ^ new_n5323_) : (~new_n5305_ ^ new_n5323_);
  assign new_n5304_ = (new_n5216_ & new_n5246_) | (new_n5165_ & (new_n5216_ | new_n5246_));
  assign new_n5305_ = new_n5306_ ? (new_n5307_ ^ new_n5320_) : (~new_n5307_ ^ new_n5320_);
  assign new_n5306_ = (new_n5190_ & new_n5191_) | (new_n5166_ & (new_n5190_ | new_n5191_));
  assign new_n5307_ = ~new_n5308_ ^ new_n5309_;
  assign new_n5308_ = ~new_n5181_ & new_n5167_;
  assign new_n5309_ = ~new_n5310_ ^ new_n5319_;
  assign new_n5310_ = new_n5088_ ? new_n5311_ : ((~new_n5315_ & new_n4678_) | (~new_n5079_ & new_n5318_ & ~new_n4678_));
  assign new_n5311_ = new_n5087_ ? new_n5312_ : ((~new_n5314_ & new_n5082_) | (new_n3491_ & new_n5084_ & ~new_n5082_));
  assign new_n5312_ = (new_n5189_ | new_n5313_ | new_n5089_) & (new_n5085_ | ~new_n5089_ | (\i[1959]  & ~new_n5086_));
  assign new_n5313_ = ~\i[1776]  & ~\i[1777]  & ~\i[1778]  & ~\i[1779]  & (\i[1487]  | \i[1486] );
  assign new_n5314_ = new_n5083_ ? ~new_n4879_ : ~new_n5129_;
  assign new_n5315_ = (new_n5317_ | ~new_n5080_ | (\i[1479]  & \i[1478] )) & (new_n4219_ | new_n5316_ | new_n5080_);
  assign new_n5316_ = new_n4277_ & ~\i[1728]  & ~\i[1729] ;
  assign new_n5317_ = \i[1387]  & (\i[1386]  | \i[1385] );
  assign new_n5318_ = ~new_n5077_ & ~new_n5184_;
  assign new_n5319_ = new_n4820_ & ~new_n3905_ & new_n4982_;
  assign new_n5320_ = ~new_n5321_ ^ new_n5322_;
  assign new_n5321_ = (~new_n5234_ & new_n5225_) | (~new_n5218_ & (~new_n5234_ | new_n5225_));
  assign new_n5322_ = (~new_n5207_ & new_n5201_) | (~new_n5192_ & (~new_n5207_ | new_n5201_));
  assign new_n5323_ = new_n5324_ ? (new_n5325_ ^ new_n5326_) : (~new_n5325_ ^ new_n5326_);
  assign new_n5324_ = (new_n5244_ & new_n5245_) | (~new_n5217_ & (new_n5244_ | new_n5245_));
  assign new_n5325_ = (new_n5252_ & new_n5271_) | (new_n5251_ & (new_n5252_ | new_n5271_));
  assign new_n5326_ = (~new_n5259_ & new_n5267_) | (~new_n5253_ & (~new_n5259_ | new_n5267_));
  assign new_n5327_ = new_n5328_ ? (~new_n5329_ ^ new_n5334_) : (new_n5329_ ^ new_n5334_);
  assign new_n5328_ = (new_n5282_ & new_n5290_) | (new_n5281_ & (new_n5282_ | new_n5290_));
  assign new_n5329_ = new_n5330_ ^ new_n5331_;
  assign new_n5330_ = (~new_n5285_ & new_n5284_) | (new_n5283_ & (~new_n5285_ | new_n5284_));
  assign new_n5331_ = new_n5332_ ^ new_n5333_;
  assign new_n5332_ = (new_n5286_ | (~new_n5289_ & (\i[1487]  | \i[1519]  | ~new_n5288_ | ~new_n4837_))) & (\i[1487]  | \i[1519]  | ~new_n5289_ | ~new_n5288_ | ~new_n4837_);
  assign new_n5333_ = (new_n5274_ & new_n5275_) | (~new_n5272_ & (new_n5274_ | new_n5275_));
  assign new_n5334_ = (~new_n5250_ & new_n5276_) | (new_n5249_ & (~new_n5250_ | new_n5276_));
  assign new_n5335_ = (~new_n5280_ & new_n5291_) | (new_n5279_ & (~new_n5280_ | new_n5291_));
  assign \o[17]  = ((new_n5337_ | new_n5338_) & (~new_n5339_ ^ ~new_n5340_)) | (~new_n5337_ & ~new_n5338_ & (~new_n5339_ ^ new_n5340_));
  assign new_n5337_ = ~new_n5297_ & new_n5296_;
  assign new_n5338_ = ~new_n5299_ & new_n5298_;
  assign new_n5339_ = (~new_n5301_ & new_n5335_) | (new_n5300_ & (~new_n5301_ | new_n5335_));
  assign new_n5340_ = new_n5341_ ? (~new_n5342_ ^ new_n5354_) : (new_n5342_ ^ new_n5354_);
  assign new_n5341_ = (~new_n5303_ & ~new_n5327_) | (new_n5302_ & (~new_n5303_ | ~new_n5327_));
  assign new_n5342_ = new_n5343_ ? (new_n5344_ ^ new_n5350_) : (~new_n5344_ ^ new_n5350_);
  assign new_n5343_ = (~new_n5305_ & ~new_n5323_) | (new_n5304_ & (~new_n5305_ | ~new_n5323_));
  assign new_n5344_ = new_n5345_ ? (~new_n5346_ ^ new_n5349_) : (new_n5346_ ^ new_n5349_);
  assign new_n5345_ = (~new_n5307_ & ~new_n5320_) | (new_n5306_ & (~new_n5307_ | ~new_n5320_));
  assign new_n5346_ = new_n5347_ ^ new_n5348_;
  assign new_n5347_ = ~new_n5308_ & ~new_n5309_;
  assign new_n5348_ = new_n5310_ & new_n5319_;
  assign new_n5349_ = new_n5321_ & new_n5322_;
  assign new_n5350_ = new_n5351_ ? (new_n5352_ ^ new_n5353_) : (~new_n5352_ ^ new_n5353_);
  assign new_n5351_ = (new_n5325_ & new_n5326_) | (new_n5324_ & (new_n5325_ | new_n5326_));
  assign new_n5352_ = ~new_n5331_ & new_n5330_;
  assign new_n5353_ = ~new_n5332_ & new_n5333_;
  assign new_n5354_ = (~new_n5329_ & new_n5334_) | (new_n5328_ & (~new_n5329_ | new_n5334_));
  assign \o[18]  = ~new_n5356_ ^ new_n5357_;
  assign new_n5356_ = (new_n5339_ | (~new_n5340_ & (new_n5338_ | new_n5337_))) & (new_n5338_ | new_n5337_ | ~new_n5340_);
  assign new_n5357_ = new_n5358_ ^ new_n5359_;
  assign new_n5358_ = (~new_n5342_ & new_n5354_) | (new_n5341_ & (~new_n5342_ | new_n5354_));
  assign new_n5359_ = new_n5360_ ? (~new_n5361_ ^ new_n5364_) : (new_n5361_ ^ new_n5364_);
  assign new_n5360_ = (~new_n5344_ & ~new_n5350_) | (new_n5343_ & (~new_n5344_ | ~new_n5350_));
  assign new_n5361_ = new_n5362_ ^ new_n5363_;
  assign new_n5362_ = (~new_n5346_ & new_n5349_) | (new_n5345_ & (~new_n5346_ | new_n5349_));
  assign new_n5363_ = ~new_n5347_ & ~new_n5348_;
  assign new_n5364_ = (new_n5352_ & new_n5353_) | (new_n5351_ & (new_n5352_ | new_n5353_));
  assign \o[19]  = ((new_n5366_ | new_n5367_) & (~new_n5368_ ^ new_n5369_)) | (~new_n5366_ & ~new_n5367_ & (~new_n5368_ ^ ~new_n5369_));
  assign new_n5366_ = ~new_n5357_ & new_n5356_;
  assign new_n5367_ = ~new_n5359_ & new_n5358_;
  assign new_n5368_ = (~new_n5361_ & new_n5364_) | (new_n5360_ & (~new_n5361_ | new_n5364_));
  assign new_n5369_ = ~new_n5363_ & new_n5362_;
  assign \o[20]  = (new_n5369_ | new_n5366_ | new_n5367_) & (new_n5368_ | (new_n5369_ & (new_n5366_ | new_n5367_)));
  assign \o[21]  = new_n5372_ ^ new_n5838_;
  assign new_n5372_ = new_n5373_ ? (new_n5811_ ^ new_n5830_) : (~new_n5811_ ^ new_n5830_);
  assign new_n5373_ = new_n5374_ ? (~new_n5782_ ^ new_n5798_) : (new_n5782_ ^ new_n5798_);
  assign new_n5374_ = new_n5375_ ? (new_n5500_ ^ new_n5766_) : (~new_n5500_ ^ new_n5766_);
  assign new_n5375_ = new_n5376_ ? (~new_n5473_ ^ new_n5487_) : (new_n5473_ ^ new_n5487_);
  assign new_n5376_ = new_n5377_ ? (~new_n5451_ ^ new_n5467_) : (new_n5451_ ^ new_n5467_);
  assign new_n5377_ = new_n5378_ ? (~new_n5432_ ^ new_n5447_) : (new_n5432_ ^ new_n5447_);
  assign new_n5378_ = new_n5379_ ? (~new_n5402_ ^ new_n5417_) : (new_n5402_ ^ new_n5417_);
  assign new_n5379_ = (\i[2310]  & \i[2311] ) ? (new_n5392_ | new_n5400_) : new_n5380_;
  assign new_n5380_ = (new_n5388_ & \i[2298]  & \i[2299]  & (\i[2296]  | \i[2297] )) | (new_n5381_ & (~\i[2298]  | ~\i[2299]  | (~\i[2296]  & ~\i[2297] )));
  assign new_n5381_ = new_n5385_ ? new_n5382_ : (new_n3789_ ? new_n5387_ : new_n5386_);
  assign new_n5382_ = (~new_n5384_ | ~new_n5383_) & (~\i[2753]  | ~\i[2754]  | ~\i[2755]  | new_n5383_);
  assign new_n5383_ = new_n4657_ & (~\i[1949]  | ~\i[1948] );
  assign new_n5384_ = \i[1402]  & \i[1403]  & (\i[1401]  | \i[1400] );
  assign new_n5385_ = ~\i[2539]  & (~\i[2537]  | ~\i[2538]  | ~\i[2536] );
  assign new_n5386_ = ~\i[2206]  & ~\i[2207]  & (~\i[2205]  | ~\i[2204] );
  assign new_n5387_ = \i[1751]  & \i[1749]  & \i[1750] ;
  assign new_n5388_ = new_n3462_ ? new_n5389_ : (new_n5391_ | (~new_n5078_ & ~\i[2730]  & ~\i[2731] ));
  assign new_n5389_ = (\i[1063]  & (\i[1062]  | (\i[1060]  & \i[1061] ))) ? new_n5390_ : ~new_n5034_;
  assign new_n5390_ = ~\i[1167]  & (~\i[1166]  | ~\i[1165] );
  assign new_n5391_ = new_n5078_ & \i[2407]  & (\i[2406]  | \i[2405] );
  assign new_n5392_ = ~new_n5399_ & (new_n4186_ ? (new_n5397_ ? ~new_n5398_ : new_n4225_) : new_n5393_);
  assign new_n5393_ = new_n5395_ ? (~\i[1879]  | (~new_n5396_ & ~\i[1878] )) : ~new_n5394_;
  assign new_n5394_ = ~\i[1079]  & (~\i[1078]  | ~\i[1077] );
  assign new_n5395_ = ~\i[959]  & (~\i[957]  | ~\i[958]  | ~\i[956] );
  assign new_n5396_ = \i[1876]  & \i[1877] ;
  assign new_n5397_ = \i[1283]  & (\i[1281]  | \i[1282]  | \i[1280] );
  assign new_n5398_ = \i[607]  & \i[605]  & \i[606] ;
  assign new_n5399_ = \i[2622]  & \i[2623]  & (\i[2621]  | \i[2620] );
  assign new_n5400_ = ~new_n5401_ & new_n5399_ & (\i[2619]  | (\i[2618]  & (\i[2617]  | \i[2616] )));
  assign new_n5401_ = new_n4210_ ? ~new_n3320_ : (~\i[647]  & (~\i[644]  | ~\i[645]  | ~\i[646] ));
  assign new_n5402_ = (new_n5409_ | new_n5415_ | ~new_n5416_) & (new_n5403_ | new_n5416_ | (new_n5414_ & ~new_n5412_));
  assign new_n5403_ = new_n5405_ & (~new_n5408_ | ~new_n5406_) & (\i[2431]  | ~new_n5407_ | ~new_n5404_ | new_n5406_);
  assign new_n5404_ = new_n4740_ & ~\i[2100]  & ~\i[2101] ;
  assign new_n5405_ = \i[2647]  & \i[2645]  & \i[2646] ;
  assign new_n5406_ = \i[2863]  & (\i[2862]  | (\i[2861]  & \i[2860] ));
  assign new_n5407_ = ~\i[2429]  & ~\i[2430] ;
  assign new_n5408_ = \i[1735]  & \i[1733]  & \i[1734] ;
  assign new_n5409_ = new_n5410_ & (~new_n4694_ | ~new_n4324_);
  assign new_n5410_ = ~\i[1159]  & ~new_n5411_ & (~\i[1263]  | (~\i[1261]  & ~\i[1262] ));
  assign new_n5411_ = \i[1157]  & \i[1158] ;
  assign new_n5412_ = ~new_n5413_ & ~new_n4939_ & ~\i[1771]  & (~\i[1770]  | ~\i[1769]  | ~\i[1768] );
  assign new_n5413_ = \i[2863]  & (\i[2862]  | \i[2861] );
  assign new_n5414_ = ~new_n5405_ & (\i[1035]  | ~new_n5413_ | (\i[1034]  & (\i[1032]  | \i[1033] )));
  assign new_n5415_ = ~new_n4673_ & (new_n4091_ | \i[1174]  | \i[1175] ) & (new_n5411_ | \i[1159] );
  assign new_n5416_ = \i[1499]  & (\i[1498]  | (\i[1497]  & \i[1496] ));
  assign new_n5417_ = (~new_n5427_ & ~new_n5418_ & ~new_n4019_) | (new_n4019_ & (new_n5431_ ? new_n5424_ : ~new_n5430_));
  assign new_n5418_ = ~new_n5422_ & ((new_n5419_ & new_n5423_) | (\i[519]  & ~new_n5423_ & (~\i[2619]  | ~\i[2618] )));
  assign new_n5419_ = (~new_n5421_ & ~new_n5420_) | (new_n4705_ & new_n5420_ & (\i[2409]  | \i[2408] ));
  assign new_n5420_ = ~\i[1611]  & ~\i[1609]  & ~\i[1610] ;
  assign new_n5421_ = \i[2174]  & \i[2175] ;
  assign new_n5422_ = \i[1279]  & \i[1278]  & \i[1276]  & \i[1277] ;
  assign new_n5423_ = \i[1379]  & (\i[1377]  | \i[1378]  | \i[1376] );
  assign new_n5424_ = ~new_n5425_ & (~new_n5426_ | (\i[409]  & \i[410]  & \i[411] ));
  assign new_n5425_ = ~\i[1083]  & new_n3550_ & new_n4166_ & (~\i[1082]  | (~\i[1080]  & ~\i[1081] ));
  assign new_n5426_ = ~new_n4166_ & ~\i[619]  & (~\i[618]  | ~\i[617] );
  assign new_n5427_ = new_n5422_ & (new_n5429_ ? (~new_n5428_ | ~new_n4100_) : ~new_n3417_);
  assign new_n5428_ = \i[611]  & (\i[610]  | \i[609] );
  assign new_n5429_ = ~\i[1491]  & ~\i[1489]  & ~\i[1490] ;
  assign new_n5430_ = ~new_n3498_ & ~\i[914]  & ~\i[915]  & (~\i[913]  | ~\i[912] );
  assign new_n5431_ = ~\i[942]  & ~\i[943]  & (~\i[941]  | ~\i[940] );
  assign new_n5432_ = (~\i[1711]  & (~\i[1710]  | (~\i[1708]  & ~\i[1709] ))) ? new_n5438_ : new_n5433_;
  assign new_n5433_ = new_n5437_ ? new_n5434_ : ((new_n4021_ & new_n5435_) | (~new_n5436_ & new_n4345_ & ~new_n5435_));
  assign new_n5434_ = (~\i[1174]  & ~\i[1175] ) ? new_n4440_ : ~new_n3538_;
  assign new_n5435_ = \i[2067]  & (\i[2065]  | \i[2066]  | \i[2064] );
  assign new_n5436_ = \i[1751]  & (\i[1750]  | \i[1749] );
  assign new_n5437_ = \i[635]  & (\i[633]  | \i[634]  | \i[632] );
  assign new_n5438_ = new_n3339_ ? new_n5444_ : (new_n3223_ ? new_n5439_ : new_n5441_);
  assign new_n5439_ = new_n5440_ ? (\i[1843]  & (\i[1841]  | \i[1842]  | \i[1840] )) : \i[2315] ;
  assign new_n5440_ = \i[2067]  & \i[2065]  & \i[2066] ;
  assign new_n5441_ = new_n5443_ ? new_n5442_ : \i[1303] ;
  assign new_n5442_ = \i[2754]  & \i[2755]  & (\i[2753]  | \i[2752] );
  assign new_n5443_ = \i[1839]  & (\i[1838]  | \i[1837] );
  assign new_n5444_ = new_n5445_ ? ((\i[1494]  & \i[1495] ) ? new_n4130_ : new_n5031_) : ~new_n5446_;
  assign new_n5445_ = \i[1731]  & \i[1730]  & \i[1728]  & \i[1729] ;
  assign new_n5446_ = \i[1961]  & \i[1962]  & \i[1963]  & (~\i[507]  | ~\i[506] );
  assign new_n5447_ = new_n4364_ & new_n5449_ & new_n5448_ & ~new_n5450_ & new_n5420_;
  assign new_n5448_ = ~\i[2715]  & ~\i[2713]  & ~\i[2714] ;
  assign new_n5449_ = \i[1379]  & \i[1378]  & \i[1376]  & \i[1377] ;
  assign new_n5450_ = \i[494]  & \i[495]  & (\i[493]  | \i[492] );
  assign new_n5451_ = (~new_n5457_ & ~new_n5463_ & ~new_n5462_) | (new_n5462_ & (new_n5466_ ? ~new_n5452_ : new_n5459_));
  assign new_n5452_ = ~new_n5453_ & (new_n5454_ | ~new_n4412_ | ~new_n5456_);
  assign new_n5453_ = new_n5454_ & ~new_n3867_ & ~new_n5455_;
  assign new_n5454_ = ~\i[2727]  & ~\i[2726]  & ~\i[2724]  & ~\i[2725] ;
  assign new_n5455_ = ~\i[2262]  & ~\i[2263]  & (~\i[2261]  | ~\i[2260] );
  assign new_n5456_ = ~\i[2282]  & ~\i[2283]  & (~\i[2281]  | ~\i[2280] );
  assign new_n5457_ = new_n4136_ & ((~\i[1421]  & ~\i[1422] ) | ~\i[1423]  | ~new_n5458_);
  assign new_n5458_ = new_n5048_ & (~\i[1312]  | ~\i[1313]  | ~\i[1314]  | ~\i[1315] );
  assign new_n5459_ = new_n5460_ & ~new_n5461_ & (~\i[940]  | ~\i[941]  | ~\i[942]  | ~\i[943] );
  assign new_n5460_ = \i[1179]  & (\i[1178]  | (\i[1177]  & \i[1176] ));
  assign new_n5461_ = \i[935]  & (\i[934]  | (\i[933]  & \i[932] ));
  assign new_n5462_ = new_n3409_ & (~\i[1545]  | ~\i[1544] );
  assign new_n5463_ = ~new_n4136_ & (new_n3647_ | new_n5464_ | ~new_n5465_);
  assign new_n5464_ = ~\i[1419]  & (~\i[1418]  | (~\i[1417]  & ~\i[1416] ));
  assign new_n5465_ = \i[2147]  & (\i[2146]  | \i[2145] );
  assign new_n5466_ = ~\i[495]  & (~\i[493]  | ~\i[494]  | ~\i[492] );
  assign new_n5467_ = ~new_n3348_ & ((~new_n5468_ & new_n5472_) | (~new_n5471_ & ~new_n5472_ & (new_n4651_ | new_n3627_)));
  assign new_n5468_ = (new_n5469_ | new_n5448_) & (~new_n5470_ | ~\i[1532]  | ~\i[1533]  | ~\i[1534]  | ~new_n5448_);
  assign new_n5469_ = (\i[1959]  | \i[1958]  | new_n5456_) & (\i[2378]  | \i[2379]  | ~new_n5456_);
  assign new_n5470_ = \i[1535]  & \i[1095]  & \i[1093]  & \i[1094] ;
  assign new_n5471_ = ~new_n4340_ & new_n3627_ & (~\i[1395]  | (~\i[1392]  & ~\i[1393]  & ~\i[1394] ));
  assign new_n5472_ = ~\i[491]  & (~\i[489]  | ~\i[490]  | ~\i[488] );
  assign new_n5473_ = new_n5484_ ? ((~new_n4241_ & new_n5486_) | (~new_n5482_ & ~new_n5485_ & ~new_n5486_)) : new_n5474_;
  assign new_n5474_ = new_n5481_ ? ((\i[2406]  & \i[2407] ) ? ~new_n5479_ : ~new_n5475_) : new_n5477_;
  assign new_n5475_ = new_n5476_ ? ~new_n3703_ : ~new_n4168_;
  assign new_n5476_ = new_n3539_ & (\i[1393]  | \i[1392] );
  assign new_n5477_ = (new_n5478_ | \i[1922]  | \i[1923] ) & (\i[2282]  | \i[2283]  | \i[2379]  | (~\i[1922]  & ~\i[1923] ));
  assign new_n5478_ = (~\i[2178]  | ~\i[2179] ) & (~\i[1715]  | (~\i[1714]  & ~new_n3526_));
  assign new_n5479_ = new_n5480_ & ~\i[2832]  & ~\i[2833] ;
  assign new_n5480_ = ~\i[2834]  & ~\i[2835] ;
  assign new_n5481_ = \i[2851]  & (\i[2849]  | \i[2850]  | \i[2848] );
  assign new_n5482_ = ~new_n5483_ & ~\i[2647]  & (~\i[2646]  | (~\i[2644]  & ~\i[2645] ));
  assign new_n5483_ = ~\i[1079]  & ~\i[1078]  & ~\i[1076]  & ~\i[1077] ;
  assign new_n5484_ = \i[699]  & (\i[697]  | \i[698]  | \i[696] );
  assign new_n5485_ = \i[1150]  & \i[1151] ;
  assign new_n5486_ = \i[1970]  & \i[1971]  & (\i[1969]  | \i[1968] );
  assign new_n5487_ = new_n5491_ ? ((new_n5496_ | ~new_n5498_) & (~new_n5493_ | new_n5492_)) : new_n5488_;
  assign new_n5488_ = (new_n5489_ | new_n5490_ | new_n4285_) & (~new_n4285_ | (new_n3284_ & (~\i[1403]  | ~\i[1402] )));
  assign new_n5489_ = ~\i[1431]  & new_n3350_ & (\i[2083]  | (\i[2082]  & (\i[2081]  | \i[2080] )));
  assign new_n5490_ = ~new_n3350_ & ~\i[1523]  & (~\i[1522]  | ~\i[1521] );
  assign new_n5491_ = new_n5480_ & (~\i[2833]  | ~\i[2832] );
  assign new_n5492_ = \i[1991]  & (~new_n4425_ | ~\i[1967] ) & (\i[534]  | \i[535]  | \i[533]  | \i[1967] );
  assign new_n5493_ = new_n5495_ & (new_n5494_ | \i[1991]  | (\i[1203]  & (\i[1201]  | \i[1202] )));
  assign new_n5494_ = ~\i[2178]  & ~\i[2179] ;
  assign new_n5495_ = ~\i[1431]  & (~\i[1430]  | (~\i[1429]  & ~\i[1428] ));
  assign new_n5496_ = new_n5497_ & new_n5176_ & ~\i[2255]  & ~\i[2254]  & ~\i[2252]  & ~\i[2253] ;
  assign new_n5497_ = ~\i[963]  & ~\i[961]  & ~\i[962] ;
  assign new_n5498_ = ~new_n5495_ & ((\i[1921]  & \i[1922]  & \i[1923] ) | new_n5499_ | new_n5176_);
  assign new_n5499_ = \i[759]  & (\i[758]  | (\i[757]  & \i[756] ));
  assign new_n5500_ = new_n5501_ ? (~new_n5658_ ^ new_n5451_) : (new_n5658_ ^ new_n5451_);
  assign new_n5501_ = new_n5502_ ? (new_n5595_ ^ new_n5656_) : (~new_n5595_ ^ new_n5656_);
  assign new_n5502_ = new_n5503_ ? (new_n5546_ ^ new_n5592_) : (~new_n5546_ ^ new_n5592_);
  assign new_n5503_ = new_n5504_ ? (~new_n5519_ ^ new_n5535_) : (new_n5519_ ^ new_n5535_);
  assign new_n5504_ = \i[1403]  ? ((~new_n5514_ & ~new_n3437_) | (~new_n5517_ & new_n5151_ & new_n3437_)) : new_n5505_;
  assign new_n5505_ = ~new_n5509_ & (~new_n5506_ | (~new_n4470_ & (new_n5512_ ? new_n5513_ : ~new_n3697_)));
  assign new_n5506_ = new_n3560_ & (new_n5507_ | \i[1954]  | \i[1955]  | ~new_n4470_);
  assign new_n5507_ = new_n5508_ & ~\i[2172]  & ~\i[2173] ;
  assign new_n5508_ = ~\i[2174]  & ~\i[2175] ;
  assign new_n5509_ = ~new_n5510_ & ~new_n3560_ & (new_n3451_ | (~\i[1287]  & ~new_n4334_) | (new_n5511_ & new_n4334_));
  assign new_n5510_ = ~\i[939]  & \i[611]  & new_n3451_ & (\i[610]  | (\i[608]  & \i[609] ));
  assign new_n5511_ = ~\i[2594]  & ~\i[2595]  & (~\i[2593]  | ~\i[2592] );
  assign new_n5512_ = ~\i[695]  & ~\i[693]  & ~\i[694] ;
  assign new_n5513_ = \i[1291]  & (\i[1290]  | \i[1289] );
  assign new_n5514_ = (~new_n5515_ | ~new_n4249_ | new_n3696_) & (~new_n3696_ | (~new_n4199_ & (~new_n5516_ | ~new_n5396_)));
  assign new_n5515_ = ~\i[2146]  & ~\i[2147]  & (~\i[2145]  | ~\i[2144] );
  assign new_n5516_ = \i[1878]  & \i[1879] ;
  assign new_n5517_ = new_n5518_ ? ~new_n4091_ : new_n3564_;
  assign new_n5518_ = ~\i[1946]  & ~\i[1947]  & (~\i[1945]  | ~\i[1944] );
  assign new_n5519_ = (new_n5524_ | new_n5528_ | ~new_n3301_) & (new_n5531_ | new_n3301_ | (~new_n5532_ & ~new_n5520_));
  assign new_n5520_ = new_n5522_ ? ((~new_n5523_ & ~new_n3669_) | (~new_n3658_ & new_n3659_ & new_n3669_)) : new_n5521_;
  assign new_n5521_ = (~new_n5316_ & ~new_n3670_) | (\i[1620]  & \i[1621]  & \i[1622]  & \i[1623]  & new_n3670_);
  assign new_n5522_ = ~\i[1303]  & (~\i[1302]  | ~\i[1301] );
  assign new_n5523_ = \i[1811]  & \i[1810]  & \i[1808]  & \i[1809] ;
  assign new_n5524_ = new_n3322_ & ((~new_n5525_ & new_n5526_) | (~new_n5527_ & new_n5383_ & ~new_n5526_));
  assign new_n5525_ = \i[1375]  & ~new_n5024_ & \i[1374] ;
  assign new_n5526_ = ~\i[2063]  & (~\i[2061]  | ~\i[2062]  | ~\i[2060] );
  assign new_n5527_ = \i[1754]  & \i[1755]  & (\i[1753]  | \i[1752] );
  assign new_n5528_ = ~new_n3322_ & new_n5529_ & new_n3394_ & (\i[2163]  | (\i[2161]  & \i[2162] ));
  assign new_n5529_ = \i[1625]  & new_n5530_ & \i[1624] ;
  assign new_n5530_ = \i[1626]  & \i[1627] ;
  assign new_n5531_ = new_n5532_ & new_n5384_ & ((~new_n5533_ & ~new_n5534_) | (\i[2214]  & \i[2215]  & new_n5534_));
  assign new_n5532_ = ~\i[2491]  & ~\i[2490]  & ~\i[2488]  & ~\i[2489] ;
  assign new_n5533_ = ~\i[731]  & ~\i[730]  & ~\i[728]  & ~\i[729] ;
  assign new_n5534_ = ~\i[855]  & (~\i[853]  | ~\i[854]  | ~\i[852] );
  assign new_n5535_ = ~new_n5538_ & (new_n3800_ | (~new_n5536_ & new_n4105_) | (new_n3548_ & new_n5545_ & ~new_n4105_));
  assign new_n5536_ = (~new_n5537_ | ~new_n5086_) & (new_n4323_ | ~new_n4021_ | new_n5086_);
  assign new_n5537_ = new_n3689_ & \i[1299] ;
  assign new_n5538_ = new_n5542_ & (~new_n5540_ | (new_n5390_ & (new_n5539_ ? ~new_n5544_ : new_n5543_)));
  assign new_n5539_ = new_n3225_ & ~\i[1042]  & ~\i[1043] ;
  assign new_n5540_ = ~new_n4158_ & (new_n5390_ | (~new_n4094_ & new_n5541_) | (\i[703]  & ~new_n5541_));
  assign new_n5541_ = ~\i[1599]  & ~\i[1598]  & ~\i[1596]  & ~\i[1597] ;
  assign new_n5542_ = new_n3800_ & (~new_n5390_ | ~new_n4158_ | (\i[1371]  ? new_n3575_ : new_n4012_));
  assign new_n5543_ = ~\i[1391]  & (~\i[1389]  | ~\i[1390]  | ~\i[1388] );
  assign new_n5544_ = \i[619]  & \i[617]  & \i[618] ;
  assign new_n5545_ = ~new_n4779_ & \i[2839]  & (\i[2838]  | (\i[2836]  & \i[2837] ));
  assign new_n5546_ = new_n5547_ ? (new_n5554_ ^ new_n5572_) : (~new_n5554_ ^ new_n5572_);
  assign new_n5547_ = new_n5462_ ? new_n5548_ : new_n5552_;
  assign new_n5548_ = (new_n5453_ | new_n5549_ | ~new_n5466_) & (new_n5459_ | new_n5466_ | (new_n5551_ & new_n5461_));
  assign new_n5549_ = ~new_n5454_ & (new_n5456_ ? new_n4412_ : ~new_n5550_);
  assign new_n5550_ = new_n5508_ & (~\i[2173]  | ~\i[2172] );
  assign new_n5551_ = (~\i[2110]  | ~\i[2111] ) & (~\i[2376]  | ~\i[2377]  | ~\i[2378]  | ~\i[2379] );
  assign new_n5552_ = ~new_n5553_ & (~new_n5457_ | (new_n5464_ & (~\i[1423]  | (~\i[1421]  & ~\i[1422] ))));
  assign new_n5553_ = ~new_n4136_ & (\i[914]  | \i[915]  | new_n5465_) & (new_n5464_ | new_n3647_ | ~new_n5465_);
  assign new_n5554_ = new_n5571_ ? new_n5555_ : (~new_n5564_ & (new_n5569_ | ~new_n3627_ | ~new_n5570_));
  assign new_n5555_ = new_n5561_ ? new_n5556_ : ((new_n5560_ | new_n3394_) & (new_n5562_ | ~new_n5563_ | ~new_n3394_));
  assign new_n5556_ = (new_n5557_ | ~new_n4293_) & (~new_n4328_ | ~new_n5559_ | new_n4293_);
  assign new_n5557_ = (\i[1283]  | ~new_n5558_) & (~\i[2099]  | new_n5558_ | (~\i[2098]  & (~\i[2096]  | ~\i[2097] )));
  assign new_n5558_ = ~\i[1387]  & (~\i[1386]  | (~\i[1385]  & ~\i[1384] ));
  assign new_n5559_ = ~\i[918]  & ~\i[919] ;
  assign new_n5560_ = (new_n4206_ | ~new_n4757_) & (~\i[1033]  | ~\i[1034]  | ~\i[1035]  | new_n4757_);
  assign new_n5561_ = \i[1623]  & \i[1621]  & \i[1622] ;
  assign new_n5562_ = ~\i[503]  & (~\i[501]  | ~\i[502]  | ~\i[500] );
  assign new_n5563_ = ~\i[939]  & ~\i[938]  & ~\i[936]  & ~\i[937] ;
  assign new_n5564_ = ~new_n5565_ & new_n5569_ & (new_n5566_ | (~new_n3796_ & new_n5568_) | (~new_n5567_ & ~new_n5568_));
  assign new_n5565_ = new_n5566_ & \i[738]  & \i[739]  & \i[1623]  & (\i[737]  | \i[736] );
  assign new_n5566_ = ~\i[1507]  & ~\i[1505]  & ~\i[1506] ;
  assign new_n5567_ = ~\i[1295]  & ~\i[1294]  & ~\i[1292]  & ~\i[1293] ;
  assign new_n5568_ = ~\i[983]  & ~\i[981]  & ~\i[982] ;
  assign new_n5569_ = ~\i[2399]  & (~\i[2398]  | (~\i[2397]  & ~\i[2396] ));
  assign new_n5570_ = ~new_n4660_ & new_n4656_;
  assign new_n5571_ = ~\i[2839]  & ~\i[2837]  & ~\i[2838] ;
  assign new_n5572_ = (~new_n5128_ & (new_n5591_ ? new_n5578_ : new_n5573_)) | (~new_n5582_ & ~new_n5587_ & new_n5128_);
  assign new_n5573_ = (new_n5575_ | new_n5574_ | ~new_n5576_) & (~new_n5577_ | new_n5576_ | (\i[1031]  & \i[1030] ));
  assign new_n5574_ = ~\i[2211]  & new_n3731_ & (~\i[2210]  | (~\i[2208]  & ~\i[2209] ));
  assign new_n5575_ = ~\i[2711]  & ~\i[2710]  & ~new_n3731_ & ~\i[2709] ;
  assign new_n5576_ = ~\i[915]  & ~\i[913]  & ~\i[914] ;
  assign new_n5577_ = ~\i[1259]  & ~\i[1257]  & ~\i[1258] ;
  assign new_n5578_ = (new_n5579_ | new_n5454_) & (~new_n5559_ | ~new_n5581_ | ~new_n5454_);
  assign new_n5579_ = (new_n4862_ | new_n5580_) & (~\i[2318]  | ~\i[2319]  | ~new_n5580_ | (~\i[2317]  & ~\i[2316] ));
  assign new_n5580_ = \i[2051]  & (\i[2050]  | \i[2049] );
  assign new_n5581_ = \i[1303]  & (\i[1301]  | \i[1302]  | \i[1300] );
  assign new_n5582_ = new_n5585_ & (new_n5532_ ? new_n5583_ : (new_n5148_ ? ~new_n5586_ : new_n3993_));
  assign new_n5583_ = new_n5584_ ? ~new_n4352_ : ~new_n4509_;
  assign new_n5584_ = ~\i[2179]  & ~\i[2177]  & ~\i[2178] ;
  assign new_n5585_ = ~\i[2095]  & ~\i[2093]  & ~\i[2094] ;
  assign new_n5586_ = \i[1734]  & \i[1735]  & (\i[1733]  | \i[1732] );
  assign new_n5587_ = ~new_n5585_ & ((~new_n5589_ & new_n5588_ & ~new_n4722_) | (new_n4722_ & (~new_n5590_ | ~new_n3229_)));
  assign new_n5588_ = ~\i[387]  & ~\i[386]  & ~\i[384]  & ~\i[385] ;
  assign new_n5589_ = \i[2071]  & \i[2069]  & \i[2070] ;
  assign new_n5590_ = ~\i[699]  & ~\i[697]  & ~\i[698] ;
  assign new_n5591_ = ~\i[1379]  & ~\i[1377]  & ~\i[1378] ;
  assign new_n5592_ = new_n5593_ & new_n5594_;
  assign new_n5593_ = ~\i[2087]  & ~new_n4239_ & ~\i[2663]  & \i[383]  & (~\i[2662]  | ~\i[2661] );
  assign new_n5594_ = \i[2511]  & (\i[2510]  | (\i[2509]  & \i[2508] ));
  assign new_n5595_ = new_n5596_ ? (~new_n5639_ ^ new_n5592_) : (new_n5639_ ^ new_n5592_);
  assign new_n5596_ = new_n5597_ ? (new_n5613_ ^ new_n5627_) : (~new_n5613_ ^ new_n5627_);
  assign new_n5597_ = new_n5612_ ? (new_n5607_ | (~new_n5610_ & ~new_n5609_ & new_n5611_)) : new_n5598_;
  assign new_n5598_ = new_n3633_ ? (new_n5606_ ? new_n5599_ : new_n5601_) : new_n5602_;
  assign new_n5599_ = (new_n5600_ | ~new_n5136_) & (\i[2154]  | \i[2155]  | new_n5136_ | (\i[2153]  & \i[2152] ));
  assign new_n5600_ = ~\i[1294]  & ~\i[1295]  & (~\i[1293]  | ~\i[1292] );
  assign new_n5601_ = new_n5529_ ? (~\i[1931]  & (~\i[1928]  | ~\i[1929]  | ~\i[1930] )) : ~\i[1603] ;
  assign new_n5602_ = (new_n5603_ | new_n5604_) & (~new_n3428_ | ~new_n5605_ | ~new_n5604_);
  assign new_n5603_ = (new_n4381_ | ~\i[1402]  | ~\i[1403] ) & (~\i[2714]  | ~\i[2715]  | (\i[1402]  & \i[1403] ));
  assign new_n5604_ = \i[1418]  & \i[1419]  & (\i[1417]  | \i[1416] );
  assign new_n5605_ = ~\i[1871]  & (~\i[1870]  | ~\i[1869] );
  assign new_n5606_ = ~\i[2162]  & ~\i[2163]  & (~\i[2161]  | ~\i[2160] );
  assign new_n5607_ = new_n5609_ & ((new_n5608_ & new_n4288_) | (~new_n3533_ & ~new_n4288_ & (~\i[2083]  | ~\i[2082] )));
  assign new_n5608_ = (\i[1279]  | new_n3400_) & (~\i[2629]  | ~\i[2630]  | ~\i[2631]  | ~new_n3400_);
  assign new_n5609_ = ~\i[2271]  & ~\i[2269]  & ~\i[2270] ;
  assign new_n5610_ = (~\i[2155]  & (~\i[2153]  | ~\i[2154] )) ? ~new_n4216_ : new_n4164_;
  assign new_n5611_ = ~\i[1415]  & ~\i[1414]  & ~\i[1412]  & ~\i[1413] ;
  assign new_n5612_ = ~\i[1943]  & ~\i[1941]  & ~\i[1942] ;
  assign new_n5613_ = ~new_n5618_ & (new_n3348_ | (new_n5622_ & ~new_n5626_) | (new_n5614_ & new_n5626_));
  assign new_n5614_ = (new_n5615_ | new_n4236_) & (\i[2387]  | \i[2386]  | ~new_n4236_ | (\i[2543]  & \i[2542] ));
  assign new_n5615_ = (~\i[2715]  & (~\i[2713]  | ~\i[2714] )) ? ~new_n5617_ : new_n5616_;
  assign new_n5616_ = new_n4806_ & ~\i[2272]  & ~\i[2273] ;
  assign new_n5617_ = ~\i[1151]  & ~\i[1149]  & ~\i[1150] ;
  assign new_n5618_ = new_n5619_ & new_n5620_ & (\i[2375]  | ~\i[2373]  | ~\i[2374]  | ~\i[2372] );
  assign new_n5619_ = ~\i[695]  & ~\i[2375]  & ~\i[694]  & new_n3348_ & (~\i[2871]  | ~\i[2870] );
  assign new_n5620_ = ~new_n5621_ & ((~\i[693]  & ~\i[692] ) | \i[695]  | \i[694] );
  assign new_n5621_ = ~\i[2870]  & \i[2871]  & (\i[2869]  | \i[2868] );
  assign new_n5622_ = (~new_n5072_ | ~new_n5625_ | ~new_n5624_) & (new_n5624_ | (new_n3797_ ? \i[1607]  : ~new_n5623_));
  assign new_n5623_ = ~\i[731]  & (~\i[729]  | ~\i[730]  | ~\i[728] );
  assign new_n5624_ = ~\i[2850]  & ~\i[2851] ;
  assign new_n5625_ = ~\i[1623]  & ~\i[1622]  & ~\i[1620]  & ~\i[1621] ;
  assign new_n5626_ = ~\i[2423]  & ~\i[2422]  & ~\i[2420]  & ~\i[2421] ;
  assign new_n5627_ = (new_n5637_ | ~new_n4035_ | new_n5480_) & (~new_n5480_ | (new_n5638_ ? ~new_n5633_ : ~new_n5628_));
  assign new_n5628_ = (~new_n5632_ | ~new_n3996_ | (~\i[1539]  & (~\i[1537]  | ~\i[1538] ))) & (new_n5629_ | new_n3996_);
  assign new_n5629_ = (~\i[979]  & (~\i[977]  | ~\i[978] )) ? new_n5631_ : new_n5630_;
  assign new_n5630_ = \i[2519]  & (\i[2518]  | (\i[2517]  & \i[2516] ));
  assign new_n5631_ = \i[967]  & (\i[965]  | \i[966]  | \i[964] );
  assign new_n5632_ = ~\i[1067]  & (~\i[1066]  | ~\i[1065] );
  assign new_n5633_ = ~new_n5634_ & (new_n5636_ | \i[2426]  | \i[2427]  | (\i[623]  & \i[622] ));
  assign new_n5634_ = \i[622]  & new_n5635_ & \i[623]  & ~\i[2498]  & ~\i[2499] ;
  assign new_n5635_ = ~\i[1079]  & (~\i[1078]  | (~\i[1077]  & ~\i[1076] ));
  assign new_n5636_ = new_n4372_ & (~\i[1749]  | ~\i[1748] );
  assign new_n5637_ = ~new_n5483_ & ~new_n3408_ & ~new_n4977_;
  assign new_n5638_ = \i[1187]  & (\i[1186]  | \i[1185] );
  assign new_n5639_ = new_n5655_ ? new_n5640_ : ((~new_n5647_ & new_n5101_) | (~new_n5650_ & ~new_n5653_ & ~new_n5101_));
  assign new_n5640_ = ~new_n5641_ & (~\i[2175]  | (new_n5645_ & ~new_n5646_) | (~new_n3778_ & new_n5646_));
  assign new_n5641_ = ~\i[2175]  & (new_n5643_ ? ~new_n5644_ : (new_n5642_ ? ~\i[1743]  : new_n4705_));
  assign new_n5642_ = \i[2295]  & (\i[2294]  | (\i[2293]  & \i[2292] ));
  assign new_n5643_ = \i[2063]  & (\i[2062]  | (\i[2061]  & \i[2060] ));
  assign new_n5644_ = ~\i[714]  & ~\i[715]  & ~\i[713]  & (\i[2171]  | (\i[2169]  & \i[2170] ));
  assign new_n5645_ = (~new_n3576_ & new_n4257_) | (\i[1953]  & \i[1954]  & \i[1955]  & ~new_n4257_);
  assign new_n5646_ = ~\i[1643]  & ~\i[1641]  & ~\i[1642] ;
  assign new_n5647_ = (new_n5648_ | ~new_n5649_ | new_n3557_) & (new_n3996_ | new_n4391_ | ~new_n3557_);
  assign new_n5648_ = ~\i[1655]  & (~\i[1654]  | (~\i[1653]  & ~\i[1652] ));
  assign new_n5649_ = ~\i[2098]  & ~\i[2099]  & (~\i[2097]  | ~\i[2096] );
  assign new_n5650_ = new_n5651_ & ~new_n4361_ & ~new_n5652_;
  assign new_n5651_ = ~\i[1943]  & (~\i[1942]  | (~\i[1941]  & ~\i[1940] ));
  assign new_n5652_ = \i[515]  & (\i[514]  | (\i[513]  & \i[512] ));
  assign new_n5653_ = new_n5652_ & (~new_n5654_ | (~\i[1834]  & ~\i[1835] ));
  assign new_n5654_ = ~\i[1651]  & (~\i[1650]  | ~\i[1649] );
  assign new_n5655_ = ~\i[2379]  & ~\i[2378]  & ~\i[2376]  & ~\i[2377] ;
  assign new_n5656_ = ~new_n5657_ & (new_n3633_ | new_n5612_ | new_n5605_ | ~new_n5604_ | ~new_n5581_);
  assign new_n5657_ = new_n5612_ & new_n4814_ & new_n4767_ & ~new_n5609_ & ~new_n5611_;
  assign new_n5658_ = new_n5659_ ? (new_n5755_ ^ new_n5656_) : (~new_n5755_ ^ new_n5656_);
  assign new_n5659_ = new_n5660_ ? (~new_n5707_ ^ new_n5447_) : (new_n5707_ ^ new_n5447_);
  assign new_n5660_ = new_n5661_ ? (~new_n5680_ ^ new_n5696_) : (new_n5680_ ^ new_n5696_);
  assign new_n5661_ = (~new_n5676_ & ~new_n5666_ & \i[843] ) | (~\i[843]  & (new_n5671_ | (new_n5673_ & ~new_n5662_)));
  assign new_n5662_ = (new_n5663_ | ~new_n4533_) & (new_n5665_ | ~new_n5664_ | new_n4533_);
  assign new_n5663_ = ~new_n4847_ & (~\i[2109]  | ~\i[2110]  | ~\i[2111] );
  assign new_n5664_ = \i[1255]  & \i[1254]  & \i[1252]  & \i[1253] ;
  assign new_n5665_ = \i[963]  & \i[962]  & \i[960]  & \i[961] ;
  assign new_n5666_ = ~new_n5670_ & ((\i[1383]  & (\i[1381]  | \i[1382] )) ? new_n5669_ : new_n5667_);
  assign new_n5667_ = new_n5668_ ? ~new_n3740_ : \i[1487] ;
  assign new_n5668_ = new_n4245_ & (\i[1061]  | \i[1060] );
  assign new_n5669_ = new_n3240_ ? ~new_n3399_ : ~new_n4087_;
  assign new_n5670_ = \i[1278]  & \i[1279]  & (\i[1277]  | \i[1276] );
  assign new_n5671_ = new_n5672_ & ((~\i[1054]  & ~\i[1055] ) ? ~new_n5674_ : new_n3659_);
  assign new_n5672_ = ~new_n5673_ & (~\i[2872]  | ~\i[2873]  | ~\i[2874]  | ~\i[2875] );
  assign new_n5673_ = \i[1155]  & (\i[1154]  | \i[1153] );
  assign new_n5674_ = new_n5675_ & (~\i[621]  | ~\i[620] );
  assign new_n5675_ = ~\i[622]  & ~\i[623] ;
  assign new_n5676_ = new_n5670_ & ((~new_n5677_ & ~new_n5460_) | (~new_n5679_ & new_n4190_ & new_n5460_));
  assign new_n5677_ = ~new_n5678_ & (\i[701]  | \i[702]  | \i[703] );
  assign new_n5678_ = ~\i[1871]  & ~\i[1870]  & ~\i[1868]  & ~\i[1869] ;
  assign new_n5679_ = \i[1750]  & \i[1751] ;
  assign new_n5680_ = (new_n5686_ | new_n5688_ | ~new_n3672_) & (new_n3672_ | (new_n5651_ ? new_n5694_ : new_n5681_));
  assign new_n5681_ = new_n3564_ ? ~new_n5685_ : new_n5682_;
  assign new_n5682_ = (new_n5683_ | new_n5684_) & (\i[2147]  | ~new_n5684_ | (\i[2146]  & (\i[2144]  | \i[2145] )));
  assign new_n5683_ = ~\i[739]  & ~\i[738]  & ~\i[736]  & ~\i[737] ;
  assign new_n5684_ = ~\i[927]  & ~\i[926]  & ~\i[924]  & ~\i[925] ;
  assign new_n5685_ = \i[1843]  & (\i[1842]  | (\i[1841]  & \i[1840] ));
  assign new_n5686_ = new_n4328_ & ((~new_n5687_ & ~new_n4078_) | (new_n4291_ & new_n5563_ & new_n4078_));
  assign new_n5687_ = new_n3533_ ? new_n4703_ : (\i[1747]  & (\i[1744]  | \i[1745]  | \i[1746] ));
  assign new_n5688_ = ~new_n5689_ & ~new_n4328_ & (new_n5693_ | ~new_n5692_ | new_n3754_);
  assign new_n5689_ = ~new_n5692_ & (new_n5691_ | ~new_n5690_) & (~\i[701]  | ~\i[702]  | ~\i[703]  | new_n5690_);
  assign new_n5690_ = \i[2323]  & (\i[2322]  | (\i[2321]  & \i[2320] ));
  assign new_n5691_ = ~\i[1511]  & (~\i[1510]  | (~\i[1509]  & ~\i[1508] ));
  assign new_n5692_ = \i[2299]  & (\i[2298]  | (\i[2297]  & \i[2296] ));
  assign new_n5693_ = \i[1411]  & (\i[1410]  | \i[1409] );
  assign new_n5694_ = new_n4930_ ? (new_n3230_ ? ~new_n3801_ : new_n5695_) : ~new_n5158_;
  assign new_n5695_ = \i[2407]  & \i[2406]  & \i[2404]  & \i[2405] ;
  assign new_n5696_ = ~new_n5705_ & ((~new_n5697_ & new_n5450_) | ~new_n5448_ | new_n5702_);
  assign new_n5697_ = (~new_n5698_ | new_n5700_ | ~new_n5699_) & (new_n5699_ | (new_n3750_ ? new_n5701_ : new_n5150_));
  assign new_n5698_ = new_n4057_ & (~\i[1389]  | ~\i[1388] );
  assign new_n5699_ = ~\i[627]  & (~\i[625]  | ~\i[626]  | ~\i[624] );
  assign new_n5700_ = ~\i[815]  & ~\i[814]  & ~\i[812]  & ~\i[813] ;
  assign new_n5701_ = \i[1298]  & \i[1299]  & (\i[1297]  | \i[1296] );
  assign new_n5702_ = ~new_n5450_ & ((~new_n5703_ & ~new_n5704_ & ~new_n4364_) | (new_n4364_ & (\i[1059]  | new_n5449_)));
  assign new_n5703_ = new_n4158_ & ~\i[1264]  & ~\i[1265] ;
  assign new_n5704_ = \i[947]  & \i[945]  & \i[946] ;
  assign new_n5705_ = new_n5706_ & (new_n3572_ | \i[1081]  | \i[1082]  | \i[1083] );
  assign new_n5706_ = ~new_n5448_ & ~\i[2171]  & (~\i[879]  | (~\i[876]  & ~\i[877]  & ~\i[878] ));
  assign new_n5707_ = new_n5708_ ? (~new_n5727_ ^ new_n5745_) : (new_n5727_ ^ new_n5745_);
  assign new_n5708_ = (new_n5715_ | ~new_n5726_) & (new_n5709_ | new_n5723_ | new_n5726_);
  assign new_n5709_ = new_n5472_ & (new_n5714_ ? (new_n5712_ ? ~\i[1159]  : ~new_n5713_) : ~new_n5710_);
  assign new_n5710_ = new_n3781_ ? ~new_n5711_ : ~\i[1771] ;
  assign new_n5711_ = ~\i[871]  & ~\i[870]  & ~\i[868]  & ~\i[869] ;
  assign new_n5712_ = \i[719]  & (\i[717]  | \i[718]  | \i[716] );
  assign new_n5713_ = ~\i[499]  & (~\i[498]  | ~\i[497] );
  assign new_n5714_ = ~\i[1422]  & ~\i[1423]  & (~\i[1421]  | ~\i[1420] );
  assign new_n5715_ = ~new_n5716_ & (~new_n4835_ | (~new_n5722_ & (new_n3399_ ? ~new_n5721_ : ~new_n5720_)));
  assign new_n5716_ = ~new_n4835_ & (new_n4900_ ? (new_n3240_ ? ~new_n5717_ : ~new_n5719_) : new_n5718_);
  assign new_n5717_ = new_n5230_ & ~\i[2164]  & ~\i[2165] ;
  assign new_n5718_ = (new_n3557_ & new_n4275_) | (~\i[2831]  & ~new_n4275_ & (~\i[2830]  | ~\i[2829] ));
  assign new_n5719_ = \i[843]  & (\i[842]  | \i[841] );
  assign new_n5720_ = \i[1851]  & (\i[1849]  | \i[1850]  | \i[1848] );
  assign new_n5721_ = \i[1862]  & \i[1863]  & (\i[1861]  | \i[1860] );
  assign new_n5722_ = \i[2854]  & \i[2855]  & (\i[2853]  | \i[2852] );
  assign new_n5723_ = ~new_n5472_ & ((~new_n5724_ & ~new_n5725_ & new_n3569_) | (~new_n3368_ & new_n3639_ & ~new_n3569_));
  assign new_n5724_ = ~\i[2215]  & (~\i[2214]  | (~\i[2213]  & ~\i[2212] ));
  assign new_n5725_ = ~\i[499]  & (~\i[497]  | ~\i[498]  | ~\i[496] );
  assign new_n5726_ = \i[1634]  & \i[1635]  & (\i[1633]  | \i[1632] );
  assign new_n5727_ = new_n5743_ ? new_n5728_ : ((~new_n5741_ | ~new_n5744_) & (new_n5739_ | new_n5736_ | new_n5744_));
  assign new_n5728_ = new_n5735_ ? (new_n5729_ | (new_n4094_ & new_n5472_ & new_n5730_)) : new_n5731_;
  assign new_n5729_ = ~\i[1515]  & ~new_n5730_ & ~\i[1514]  & \i[2399]  & (\i[2398]  | \i[2397] );
  assign new_n5730_ = \i[1643]  & (\i[1642]  | \i[1641] );
  assign new_n5731_ = new_n5494_ ? ((~new_n4424_ & ~new_n5733_) | (~new_n5732_ & \i[2075]  & new_n5733_)) : new_n5734_;
  assign new_n5732_ = ~\i[2074]  & (~\i[2073]  | ~\i[2072] );
  assign new_n5733_ = ~\i[1539]  & ~\i[1538]  & ~\i[1536]  & ~\i[1537] ;
  assign new_n5734_ = ~\i[2271]  & (~\i[711]  | ~\i[710] ) & (~\i[2269]  | ~\i[2270]  | ~\i[2268] );
  assign new_n5735_ = \i[1531]  & (\i[1530]  | (\i[1529]  & \i[1528] ));
  assign new_n5736_ = new_n5738_ & new_n5008_ & new_n5737_;
  assign new_n5737_ = ~\i[1087]  & (~\i[1085]  | ~\i[1086]  | ~\i[1084] );
  assign new_n5738_ = \i[1975]  & \i[1974]  & \i[1972]  & \i[1973] ;
  assign new_n5739_ = ~new_n5008_ & ((~new_n4226_ & ~new_n5740_) | (~\i[1387]  & new_n5740_ & (~\i[1386]  | ~\i[1385] )));
  assign new_n5740_ = \i[2218]  & \i[2219] ;
  assign new_n5741_ = new_n5742_ & ~\i[1710]  & ~\i[1711] ;
  assign new_n5742_ = \i[1171]  & \i[1170]  & \i[1168]  & \i[1169] ;
  assign new_n5743_ = ~\i[1719]  & (~\i[1718]  | (~\i[1717]  & ~\i[1716] ));
  assign new_n5744_ = \i[1271]  & (\i[1269]  | \i[1270]  | \i[1268] );
  assign new_n5745_ = new_n5754_ ? ((new_n5751_ | new_n5748_ | ~new_n4239_) & (~new_n5746_ | new_n4239_)) : new_n5752_;
  assign new_n5746_ = (new_n5384_ | new_n5747_ | \i[383] ) & (~\i[383]  | (new_n5594_ ? \i[2087]  : ~new_n5022_));
  assign new_n5747_ = ~\i[1299]  & (~\i[1297]  | ~\i[1298]  | ~\i[1296] );
  assign new_n5748_ = new_n5750_ & ((~new_n4389_ & ~new_n5749_) | (\i[1847]  & new_n5749_ & (\i[1846]  | \i[1845] )));
  assign new_n5749_ = ~\i[1191]  & (~\i[1190]  | (~\i[1189]  & ~\i[1188] ));
  assign new_n5750_ = ~\i[1743]  & (~\i[1741]  | ~\i[1742]  | ~\i[1740] );
  assign new_n5751_ = ~new_n5750_ & ~new_n4467_ & \i[2059]  & (\i[2058]  | \i[2057]  | \i[2056] );
  assign new_n5752_ = (~new_n3445_ | ~new_n5753_) & (~\i[2088]  | ~\i[2089]  | ~\i[2090]  | ~\i[2091]  | new_n5753_);
  assign new_n5753_ = \i[2443]  & \i[2442]  & \i[2440]  & \i[2441] ;
  assign new_n5754_ = ~\i[2663]  & (~\i[2662]  | ~\i[2661] );
  assign new_n5755_ = ~new_n5756_ & (~new_n5760_ | ((~new_n5763_ | ~new_n4470_) & (new_n5764_ | new_n5765_ | new_n4470_)));
  assign new_n5756_ = new_n5757_ & (new_n5759_ | ((~new_n5761_ | new_n4463_) & (new_n4057_ | new_n5762_ | ~new_n4463_)));
  assign new_n5757_ = ~new_n5760_ & (~new_n5758_ | (new_n3361_ & (new_n4217_ ? \i[2075]  : new_n3854_)));
  assign new_n5758_ = new_n5759_ & (new_n3361_ | \i[1047]  | ~new_n3717_ | (\i[1046]  & \i[1045] ));
  assign new_n5759_ = \i[1271]  & (\i[1270]  | (\i[1269]  & \i[1268] ));
  assign new_n5760_ = \i[1374]  & \i[1375]  & (\i[1373]  | \i[1372] );
  assign new_n5761_ = \i[1387]  & \i[1386]  & \i[1311]  & \i[1309]  & \i[1310] ;
  assign new_n5762_ = ~\i[947]  & ~\i[946]  & ~\i[944]  & ~\i[945] ;
  assign new_n5763_ = new_n4167_ & ~\i[1488]  & ~\i[1489] ;
  assign new_n5764_ = ~new_n4441_ & (~\i[2519]  | ~new_n3242_ | (~\i[2516]  & ~\i[2517]  & ~\i[2518] ));
  assign new_n5765_ = new_n4441_ & new_n3703_ & \i[2763]  & (\i[2762]  | (\i[2760]  & \i[2761] ));
  assign new_n5766_ = (~new_n5776_ & ~new_n5767_ & ~new_n5781_) | (new_n5781_ & (new_n5774_ | (~new_n5772_ & ~new_n4340_)));
  assign new_n5767_ = new_n3288_ & (new_n5771_ ? new_n5768_ : (new_n5770_ ? \i[2507]  : new_n5125_));
  assign new_n5768_ = new_n5646_ ? new_n5769_ : \i[2215] ;
  assign new_n5769_ = new_n4471_ & (~\i[1273]  | ~\i[1272] );
  assign new_n5770_ = \i[1619]  & (\i[1617]  | \i[1618]  | \i[1616] );
  assign new_n5771_ = ~\i[2503]  & ~\i[2502]  & ~\i[2500]  & ~\i[2501] ;
  assign new_n5772_ = (~new_n5416_ | new_n5041_ | ~new_n5052_) & (new_n5052_ | (new_n4417_ ? ~new_n5773_ : ~new_n4463_));
  assign new_n5773_ = \i[1163]  & (\i[1162]  | \i[1161] );
  assign new_n5774_ = new_n4340_ & (new_n3854_ ? new_n5775_ : (\i[2875]  | new_n5624_));
  assign new_n5775_ = ~new_n5617_ & (~\i[1059]  | ~\i[1058] );
  assign new_n5776_ = ~new_n3288_ & (new_n5779_ | ~new_n5777_ | ~new_n5778_) & (~new_n5780_ | new_n3703_ | new_n5778_);
  assign new_n5777_ = ~\i[523]  & (~\i[522]  | (~\i[521]  & ~\i[520] ));
  assign new_n5778_ = ~\i[1839]  & (~\i[1838]  | (~\i[1837]  & ~\i[1836] ));
  assign new_n5779_ = \i[1255]  & (\i[1254]  | \i[1253] );
  assign new_n5780_ = ~\i[2599]  & ~\i[2597]  & ~\i[2598] ;
  assign new_n5781_ = ~\i[1719]  & (~\i[1718]  | ~\i[1717] );
  assign new_n5782_ = (new_n5783_ & (\i[804]  | \i[805]  | \i[806]  | \i[807] )) | (new_n5789_ & ~\i[804]  & ~\i[805]  & ~\i[806]  & ~\i[807] );
  assign new_n5783_ = (new_n5784_ | new_n5032_) & (~new_n3625_ | ~new_n5032_ | (new_n5787_ ? new_n5788_ : ~new_n4028_));
  assign new_n5784_ = new_n5098_ ? ~new_n5785_ : ((~new_n4912_ | ~new_n5786_) & (~\i[1178]  | ~\i[1179]  | new_n5786_));
  assign new_n5785_ = ~new_n5404_ & (\i[2112]  | \i[2113]  | \i[2114]  | \i[2115] );
  assign new_n5786_ = ~\i[1147]  & (~\i[1145]  | ~\i[1146]  | ~\i[1144] );
  assign new_n5787_ = ~\i[2619]  & (~\i[2617]  | ~\i[2618]  | ~\i[2616] );
  assign new_n5788_ = ~\i[915]  & ~\i[914]  & ~\i[912]  & ~\i[913] ;
  assign new_n5789_ = new_n5139_ ? new_n5790_ : ((new_n5795_ | ~new_n5012_) & (new_n5797_ | ~new_n5796_ | new_n5012_));
  assign new_n5790_ = (~new_n4171_ | new_n5793_ | new_n5792_) & (new_n5791_ | ~new_n5792_ | (new_n5794_ & ~new_n3634_));
  assign new_n5791_ = new_n3634_ & (\i[2028]  | \i[2029]  | \i[2030]  | \i[2031] );
  assign new_n5792_ = ~\i[1171]  & (~\i[1169]  | ~\i[1170]  | ~\i[1168] );
  assign new_n5793_ = \i[495]  & (\i[494]  | (\i[493]  & \i[492] ));
  assign new_n5794_ = \i[1275]  & (\i[1274]  | (\i[1273]  & \i[1272] ));
  assign new_n5795_ = (~new_n3265_ & ~\i[1169]  & ~\i[1170]  & ~\i[1171] ) | (new_n4334_ & (\i[1169]  | \i[1170]  | \i[1171] ));
  assign new_n5796_ = ~\i[1159]  & (~\i[1158]  | (~\i[1157]  & ~\i[1156] ));
  assign new_n5797_ = ~\i[934]  & ~\i[935]  & (~\i[933]  | ~\i[932] );
  assign new_n5798_ = (new_n5799_ | \i[1595]  | (\i[1593]  & \i[1594] )) & (new_n5809_ | ~new_n5810_ | (~\i[1595]  & (~\i[1593]  | ~\i[1594] )));
  assign new_n5799_ = new_n5808_ ? new_n5800_ : (new_n5805_ | (~new_n5807_ & new_n5006_));
  assign new_n5800_ = (new_n5801_ | ~new_n5803_) & (~new_n4651_ | ~new_n5804_ | new_n5803_);
  assign new_n5801_ = (~\i[515]  & (~\i[513]  | ~\i[514] )) ? ~\i[2855]  : new_n5802_;
  assign new_n5802_ = ~\i[1183]  & ~\i[1182]  & ~\i[1180]  & ~\i[1181] ;
  assign new_n5803_ = ~\i[2214]  & ~\i[2215]  & (~\i[2213]  | ~\i[2212] );
  assign new_n5804_ = ~\i[947]  & (~\i[946]  | ~\i[945] );
  assign new_n5805_ = ~new_n5806_ & ~new_n5006_ & new_n4806_ & (~\i[2273]  | ~\i[2272] );
  assign new_n5806_ = ~\i[2723]  & (~\i[2722]  | (~\i[2721]  & ~\i[2720] ));
  assign new_n5807_ = (~new_n4369_ & (\i[1398]  | \i[1399] )) | (~\i[1398]  & ~\i[1399]  & (\i[1631]  | (\i[1629]  & \i[1630] )));
  assign new_n5808_ = ~\i[735]  & (~\i[733]  | ~\i[734]  | ~\i[732] );
  assign new_n5809_ = (new_n5068_ | ~new_n5200_ | new_n3625_) & (~new_n3521_ | ~new_n3625_ | (\i[2323]  & \i[2322] ));
  assign new_n5810_ = ~\i[1146]  & ~\i[1147] ;
  assign new_n5811_ = (new_n4167_ & (~\i[1488]  | ~\i[1489] )) ? new_n5823_ : new_n5812_;
  assign new_n5812_ = new_n5822_ ? new_n5817_ : (~new_n5813_ & (new_n5816_ | ~new_n4244_ | ~\i[1155] ));
  assign new_n5813_ = new_n5814_ & (~\i[1427]  | new_n5815_ | (~\i[1424]  & ~\i[1425]  & ~\i[1426] ));
  assign new_n5814_ = new_n5816_ & (~new_n5815_ | ~\i[938]  | ~\i[939]  | (~\i[937]  & ~\i[936] ));
  assign new_n5815_ = \i[915]  & (\i[914]  | (\i[913]  & \i[912] ));
  assign new_n5816_ = ~\i[611]  & (~\i[610]  | ~\i[609] );
  assign new_n5817_ = (new_n5818_ | ~new_n5821_) & (\i[1153]  | \i[1154]  | \i[1155]  | ~new_n3905_ | new_n5821_);
  assign new_n5818_ = (new_n5819_ | ~new_n5820_) & (~\i[1193]  | ~\i[1194]  | ~\i[1195]  | new_n5820_);
  assign new_n5819_ = ~\i[2155]  & ~\i[2153]  & ~\i[2154] ;
  assign new_n5820_ = \i[1311]  & \i[1310]  & \i[1308]  & \i[1309] ;
  assign new_n5821_ = \i[2603]  & (\i[2602]  | (\i[2601]  & \i[2600] ));
  assign new_n5822_ = ~\i[1287]  & (~\i[1285]  | ~\i[1286]  | ~\i[1284] );
  assign new_n5823_ = ~new_n5824_ & (~new_n5829_ | (~new_n5497_ & (new_n4716_ ? new_n4902_ : ~new_n5440_)));
  assign new_n5824_ = new_n5828_ & (new_n5827_ ? (~new_n5512_ | new_n5769_) : new_n5825_);
  assign new_n5825_ = new_n5826_ ? ~new_n4245_ : ~new_n3309_;
  assign new_n5826_ = \i[2214]  & \i[2215]  & (\i[2213]  | \i[2212] );
  assign new_n5827_ = ~\i[1171]  & (~\i[1170]  | (~\i[1169]  & ~\i[1168] ));
  assign new_n5828_ = ~\i[2095]  & ~\i[2094]  & ~\i[2092]  & ~\i[2093] ;
  assign new_n5829_ = ~new_n5828_ & (new_n5699_ | ~new_n5497_ | (\i[1195]  & (\i[1193]  | \i[1194] )));
  assign new_n5830_ = ~new_n5831_ & (new_n5836_ | ~new_n5835_ | ~new_n5837_);
  assign new_n5831_ = (~new_n5516_ | (~\i[1876]  & ~\i[1877] )) & (new_n5416_ ? new_n5832_ : new_n5834_);
  assign new_n5832_ = (~new_n5833_ | ~new_n5796_) & (new_n4851_ | new_n5796_ | (\i[1955]  & (\i[1953]  | \i[1954] )));
  assign new_n5833_ = (~\i[2622]  & ~\i[2623]  & ~\i[1055] ) | (\i[1055]  & (~\i[2211]  | ~\i[2210] ));
  assign new_n5834_ = ~new_n4760_ & (\i[1753]  | \i[1754]  | \i[1755]  | ~new_n3452_);
  assign new_n5835_ = ~new_n5404_ & new_n5516_ & (\i[1877]  | \i[1876] );
  assign new_n5836_ = \i[1943]  & \i[1941]  & \i[1942] ;
  assign new_n5837_ = ~\i[1595]  & ~\i[1594]  & ~\i[1592]  & ~\i[1593] ;
  assign new_n5838_ = (~\i[1378]  & ~\i[1379] ) ? new_n5839_ : (new_n5857_ ? new_n5848_ : new_n5853_);
  assign new_n5839_ = ~new_n5840_ & (~new_n4948_ | (~new_n3377_ & ~new_n5847_ & new_n5846_) | (~new_n5844_ & ~new_n5846_));
  assign new_n5840_ = ~new_n4948_ & ~new_n5841_ & (new_n5842_ | (new_n5843_ & new_n4303_) | (~new_n4279_ & ~new_n4303_));
  assign new_n5841_ = new_n5842_ & ((~\i[2607]  & (~\i[2605]  | ~\i[2606] )) ? ~new_n5700_ : new_n4337_);
  assign new_n5842_ = new_n3309_ & ~\i[1072]  & ~\i[1073] ;
  assign new_n5843_ = ~\i[2751]  & ~\i[2750]  & ~\i[2748]  & ~\i[2749] ;
  assign new_n5844_ = (~\i[1822]  & ~\i[1823] ) ? new_n5845_ : ~new_n5626_;
  assign new_n5845_ = ~\i[1402]  & ~\i[1403]  & (~\i[1401]  | ~\i[1400] );
  assign new_n5846_ = ~\i[2371]  & ~\i[2370]  & ~\i[2368]  & ~\i[2369] ;
  assign new_n5847_ = ~\i[1943]  & (~\i[1942]  | ~\i[1941] );
  assign new_n5848_ = (\i[1043]  | new_n5852_) & (new_n5851_ | new_n5849_ | ~new_n5852_);
  assign new_n5849_ = ~new_n5850_ & (~\i[607]  | (~\i[606]  & (~\i[605]  | ~\i[604] )));
  assign new_n5850_ = \i[1511]  & (\i[1510]  | (\i[1509]  & \i[1508] ));
  assign new_n5851_ = ~\i[1971]  & new_n5850_ & (~\i[1970]  | ~\i[1969]  | ~\i[1968] );
  assign new_n5852_ = ~\i[503]  & (~\i[502]  | ~\i[501] );
  assign new_n5853_ = (~new_n5855_ | ~new_n5856_ | \i[1043] ) & (new_n5854_ | ~\i[1043]  | (\i[1403]  & new_n3618_));
  assign new_n5854_ = ~\i[1403]  & ~\i[2603]  & (~\i[2602]  | (~\i[2600]  & ~\i[2601] ));
  assign new_n5855_ = ~\i[590]  & ~\i[591]  & (~\i[589]  | ~\i[588] );
  assign new_n5856_ = \i[1294]  & \i[1295]  & (\i[1293]  | \i[1292] );
  assign new_n5857_ = \i[1179]  & (\i[1178]  | \i[1177] );
  assign \o[22]  = new_n5859_ ? (new_n5860_ ^ new_n5861_) : (~new_n5860_ ^ new_n5861_);
  assign new_n5859_ = ~new_n5372_ & ~new_n5838_;
  assign new_n5860_ = (~new_n5811_ & ~new_n5830_) | (new_n5373_ & (~new_n5811_ | ~new_n5830_));
  assign new_n5861_ = new_n5862_ ? (~new_n5863_ ^ new_n5967_) : (new_n5863_ ^ new_n5967_);
  assign new_n5862_ = (~new_n5782_ & ~new_n5798_) | (new_n5374_ & (~new_n5782_ | ~new_n5798_));
  assign new_n5863_ = new_n5864_ ? (~new_n5865_ ^ new_n5966_) : (new_n5865_ ^ new_n5966_);
  assign new_n5864_ = (~new_n5766_ & new_n5500_) | (new_n5375_ & (~new_n5766_ | new_n5500_));
  assign new_n5865_ = new_n5866_ ? (new_n5881_ ^ new_n5965_) : (~new_n5881_ ^ new_n5965_);
  assign new_n5866_ = new_n5867_ ? (~new_n5868_ ^ new_n5880_) : (new_n5868_ ^ new_n5880_);
  assign new_n5867_ = (new_n5451_ & new_n5467_) | (~new_n5377_ & (new_n5451_ | new_n5467_));
  assign new_n5868_ = new_n5869_ ? (new_n5870_ ^ new_n5878_) : (~new_n5870_ ^ new_n5878_);
  assign new_n5869_ = (new_n5432_ & new_n5447_) | (~new_n5378_ & (new_n5432_ | new_n5447_));
  assign new_n5870_ = new_n5871_ ? (~new_n5872_ ^ new_n5873_) : (new_n5872_ ^ new_n5873_);
  assign new_n5871_ = (new_n5402_ & new_n5417_) | (~new_n5379_ & (new_n5402_ | new_n5417_));
  assign new_n5872_ = (~new_n5727_ & ~new_n5745_) | (new_n5708_ & (~new_n5727_ | ~new_n5745_));
  assign new_n5873_ = new_n5874_ ? (~new_n5876_ ^ new_n5877_) : (new_n5876_ ^ new_n5877_);
  assign new_n5874_ = (new_n5472_ | ~new_n5875_ | ~new_n3569_ | new_n5726_) & (~new_n5722_ | ~new_n4835_ | ~new_n5726_);
  assign new_n5875_ = ~new_n5725_ & new_n5724_;
  assign new_n5876_ = ~new_n5484_ & ~new_n5476_ & ~new_n4168_ & new_n5481_ & (~\i[2407]  | ~\i[2406] );
  assign new_n5877_ = new_n5743_ & new_n3672_ & new_n4328_ & ~new_n5563_ & new_n4078_;
  assign new_n5878_ = (~new_n4217_ | ~new_n5879_ | ~new_n5759_ | new_n5760_) & (~new_n5765_ | new_n4470_ | ~new_n5760_);
  assign new_n5879_ = ~\i[2075]  & new_n3361_;
  assign new_n5880_ = (~new_n5755_ & ~new_n5656_) | (~new_n5659_ & (~new_n5755_ | ~new_n5656_));
  assign new_n5881_ = new_n5882_ ? (new_n5943_ ^ new_n5964_) : (~new_n5943_ ^ new_n5964_);
  assign new_n5882_ = new_n5883_ ? (new_n5919_ ^ new_n5942_) : (~new_n5919_ ^ new_n5942_);
  assign new_n5883_ = new_n5884_ ? (new_n5904_ ^ new_n5905_) : (~new_n5904_ ^ new_n5905_);
  assign new_n5884_ = new_n5885_ ? (new_n5890_ ^ new_n5899_) : (~new_n5890_ ^ new_n5899_);
  assign new_n5885_ = ~new_n5886_ & ((~\i[1378]  & ~\i[1379] ) | (~new_n5888_ & (new_n5857_ | new_n5889_)));
  assign new_n5886_ = new_n5887_ & (new_n4948_ | (~new_n5841_ & (new_n5842_ | (new_n4303_ & new_n5843_))));
  assign new_n5887_ = ~\i[1378]  & ~\i[1379]  & (new_n5846_ | \i[1822]  | \i[1823]  | ~new_n4948_);
  assign new_n5888_ = new_n5857_ & (new_n5852_ ? ~new_n5851_ : (\i[1043]  | ~new_n3396_));
  assign new_n5889_ = ~\i[1043]  & ~\i[1035]  & ~\i[1034]  & ~\i[1033]  & ~new_n5855_ & ~\i[1032] ;
  assign new_n5890_ = new_n3301_ ? ((new_n5898_ | new_n5526_ | ~new_n3322_) & (new_n5891_ | new_n3322_)) : new_n5894_;
  assign new_n5891_ = ~new_n5893_ & (~new_n5892_ | (~\i[695]  & (~\i[694]  | (~\i[692]  & ~\i[693] ))));
  assign new_n5892_ = ~new_n5529_ & (~\i[1195]  | (~\i[1192]  & ~\i[1193]  & ~\i[1194] ));
  assign new_n5893_ = ~new_n3715_ & ~\i[2163]  & new_n5529_ & (~\i[2162]  | ~\i[2161] );
  assign new_n5894_ = ~new_n5895_ & (new_n5532_ | ~new_n3670_ | ~new_n5897_);
  assign new_n5895_ = ~new_n5384_ & new_n5532_ & (new_n4955_ ? ~new_n5896_ : ~new_n5780_);
  assign new_n5896_ = ~\i[2855]  & ~\i[2854]  & ~\i[2852]  & ~\i[2853] ;
  assign new_n5897_ = \i[1623]  & \i[1622]  & \i[1621]  & ~new_n5522_ & \i[1620] ;
  assign new_n5898_ = new_n5383_ ? ~new_n5527_ : (~\i[695]  & (~\i[692]  | ~\i[693]  | ~\i[694] ));
  assign new_n5899_ = (new_n4167_ & (~\i[1488]  | ~\i[1489] )) ? new_n5902_ : new_n5900_;
  assign new_n5900_ = (~new_n5819_ | ~new_n5820_ | ~new_n5821_ | ~new_n5822_) & (new_n5901_ | new_n5814_ | new_n5822_);
  assign new_n5901_ = ~new_n5816_ & (\i[1155]  | (\i[1161]  & \i[1162]  & \i[1163] ));
  assign new_n5902_ = (new_n5440_ | new_n5497_ | new_n4716_ | new_n5828_) & (~new_n5903_ | new_n5827_ | ~new_n5828_);
  assign new_n5903_ = new_n4245_ & new_n5826_;
  assign new_n5904_ = (~new_n5535_ & new_n5519_) | (new_n5504_ & (~new_n5535_ | new_n5519_));
  assign new_n5905_ = new_n5906_ ^ new_n5915_;
  assign new_n5906_ = new_n3800_ ? new_n5907_ : ((~new_n5914_ & new_n4105_) | (~new_n5912_ & ~new_n5911_ & ~new_n4105_));
  assign new_n5907_ = new_n4158_ ? (~new_n5909_ & (new_n4012_ | \i[1371]  | ~new_n5390_)) : new_n5908_;
  assign new_n5908_ = (~new_n5544_ | ~new_n5539_ | ~new_n5390_) & (new_n5390_ | (new_n5541_ ? new_n4094_ : ~\i[703] ));
  assign new_n5909_ = new_n5910_ & (new_n3697_ | ~\i[1051]  | (~\i[1050]  & (~\i[1048]  | ~\i[1049] )));
  assign new_n5910_ = ~new_n5390_ & (\i[2141]  | \i[2142]  | \i[2143]  | ~new_n3697_);
  assign new_n5911_ = new_n3548_ & (new_n5545_ | (~new_n4756_ & new_n4779_));
  assign new_n5912_ = ~new_n3548_ & (new_n4471_ | new_n5913_) & (\i[2857]  | \i[2858]  | \i[2859]  | ~new_n5913_);
  assign new_n5913_ = ~\i[2627]  & ~\i[2625]  & ~\i[2626] ;
  assign new_n5914_ = (new_n5537_ | ~new_n5086_) & (new_n4021_ | ~new_n3285_ | new_n5086_);
  assign new_n5915_ = (new_n5916_ | \i[1403] ) & (~new_n3437_ | ~new_n5151_ | ~new_n5518_ | ~\i[1403] );
  assign new_n5916_ = (new_n5917_ | new_n3560_) & (new_n4470_ | new_n5512_ | ~new_n3697_ | ~new_n3560_);
  assign new_n5917_ = (new_n4413_ | new_n5918_ | ~new_n3451_) & (new_n4334_ | ~\i[1287]  | new_n3451_);
  assign new_n5918_ = \i[611]  & (\i[610]  | (\i[609]  & \i[608] ));
  assign new_n5919_ = new_n5920_ ? (~new_n5921_ ^ new_n5941_) : (new_n5921_ ^ new_n5941_);
  assign new_n5920_ = (~new_n5627_ & new_n5613_) | (~new_n5597_ & (~new_n5627_ | new_n5613_));
  assign new_n5921_ = new_n5922_ ? (~new_n5927_ ^ new_n5936_) : (new_n5927_ ^ new_n5936_);
  assign new_n5922_ = new_n5571_ ? new_n5923_ : ((new_n5926_ | ~new_n5569_) & (new_n3627_ | ~new_n5570_ | new_n5569_));
  assign new_n5923_ = (~new_n5562_ | ~new_n5924_ | new_n5561_) & (new_n5559_ | new_n4293_ | ~new_n5925_ | ~new_n5561_);
  assign new_n5924_ = \i[403]  & \i[402]  & \i[401]  & new_n3394_ & \i[400] ;
  assign new_n5925_ = ~\i[1091]  & ~\i[1089]  & ~\i[1090] ;
  assign new_n5926_ = ~new_n5565_ & (new_n5566_ | ~new_n3796_ | ~new_n5568_);
  assign new_n5927_ = (new_n5928_ & (\i[804]  | \i[805]  | \i[806]  | \i[807] )) | (new_n5933_ & ~\i[804]  & ~\i[805]  & ~\i[806]  & ~\i[807] );
  assign new_n5928_ = new_n5032_ ? new_n5929_ : (~new_n5932_ & (new_n5931_ | new_n5785_ | ~new_n5098_));
  assign new_n5929_ = (~new_n3351_ | ~new_n5930_ | new_n3625_) & (new_n4028_ | new_n5787_ | ~new_n3625_);
  assign new_n5930_ = \i[1203]  & (\i[1201]  | \i[1202]  | \i[1200] );
  assign new_n5931_ = new_n5404_ & \i[2307]  & (\i[2306]  | \i[2305]  | \i[2304] );
  assign new_n5932_ = new_n5786_ & ~new_n4912_ & ~new_n5098_;
  assign new_n5933_ = new_n5139_ ? (new_n5792_ ? ~new_n5791_ : ~new_n5935_) : ~new_n5934_;
  assign new_n5934_ = new_n5797_ & ~new_n5012_ & new_n4919_;
  assign new_n5935_ = new_n5793_ & (~\i[1727]  | ~\i[1726] );
  assign new_n5936_ = new_n5128_ ? ((new_n5937_ | ~new_n5585_) & (new_n5845_ | ~new_n5940_ | new_n5585_)) : new_n5938_;
  assign new_n5937_ = (~new_n5586_ | ~new_n5148_ | new_n5532_) & (~new_n5532_ | (new_n5584_ ? ~new_n4352_ : new_n4509_));
  assign new_n5938_ = (new_n5939_ | ~new_n5591_) & (~\i[1030]  | ~\i[1031]  | new_n5591_ | new_n5576_ | ~new_n5577_);
  assign new_n5939_ = (new_n5580_ | ~new_n4862_ | new_n5454_) & (new_n3221_ | new_n5559_ | ~new_n5454_);
  assign new_n5940_ = ~new_n4722_ & ~new_n5588_;
  assign new_n5941_ = (~new_n5554_ & ~new_n5572_) | (~new_n5547_ & (~new_n5554_ | ~new_n5572_));
  assign new_n5942_ = (new_n5546_ & new_n5592_) | (~new_n5503_ & (new_n5546_ | new_n5592_));
  assign new_n5943_ = new_n5944_ ? (~new_n5945_ ^ new_n5963_) : (new_n5945_ ^ new_n5963_);
  assign new_n5944_ = (new_n5707_ & new_n5447_) | (~new_n5660_ & (new_n5707_ | new_n5447_));
  assign new_n5945_ = new_n5946_ ? (new_n5947_ ^ new_n5954_) : (~new_n5947_ ^ new_n5954_);
  assign new_n5946_ = (~new_n5696_ & new_n5680_) | (new_n5661_ & (~new_n5696_ | new_n5680_));
  assign new_n5947_ = new_n5948_ ? (new_n5951_ ^ new_n5953_) : (~new_n5951_ ^ new_n5953_);
  assign new_n5948_ = (new_n5949_ | \i[1595]  | (\i[1593]  & \i[1594] )) & (~new_n5950_ | ~new_n5810_ | (~\i[1595]  & (~\i[1593]  | ~\i[1594] )));
  assign new_n5949_ = (~new_n5805_ | new_n5808_) & (new_n5803_ | new_n5804_ | ~new_n3468_ | ~new_n5808_);
  assign new_n5950_ = \i[2323]  & \i[2322]  & ~new_n3303_ & new_n3625_;
  assign new_n5951_ = (~new_n5952_ | ~new_n5770_) & (new_n3854_ | ~new_n5781_ | ~new_n4340_ | ~\i[2875] );
  assign new_n5952_ = new_n3288_ & ~\i[2507]  & ~new_n5781_ & ~new_n5771_;
  assign new_n5953_ = new_n3797_ & ~\i[1607]  & ~new_n5624_ & ~new_n3348_ & ~new_n5626_;
  assign new_n5954_ = new_n5955_ ? (~new_n5960_ ^ new_n5961_) : (new_n5960_ ^ new_n5961_);
  assign new_n5955_ = (~new_n5956_ & ~new_n5959_ & \i[843] ) | (~\i[843]  & (new_n5958_ | new_n5672_));
  assign new_n5956_ = new_n5957_ & new_n5670_ & ~\i[703]  & ~\i[702]  & ~new_n5460_ & ~\i[701] ;
  assign new_n5957_ = new_n5052_ & ~\i[1280]  & ~\i[1281] ;
  assign new_n5958_ = new_n5673_ & (new_n4533_ | new_n5747_ | ~new_n5665_);
  assign new_n5959_ = ~new_n5670_ & new_n3240_ & new_n3399_ & \i[1383]  & (\i[1382]  | \i[1381] );
  assign new_n5960_ = new_n5637_ & ~new_n5480_ & new_n4035_;
  assign new_n5961_ = new_n3350_ & ~new_n5962_ & ~new_n4285_ & ~new_n5491_;
  assign new_n5962_ = ~\i[1431]  & ~\i[2083]  & (~\i[2082]  | (~\i[2080]  & ~\i[2081] ));
  assign new_n5963_ = (~new_n5639_ & new_n5592_) | (~new_n5596_ & (~new_n5639_ | new_n5592_));
  assign new_n5964_ = (~new_n5656_ & new_n5595_) | (new_n5502_ & (~new_n5656_ | new_n5595_));
  assign new_n5965_ = (new_n5658_ & new_n5451_) | (new_n5501_ & (new_n5658_ | new_n5451_));
  assign new_n5966_ = (~new_n5487_ & new_n5473_) | (~new_n5376_ & (~new_n5487_ | new_n5473_));
  assign new_n5967_ = \i[2647]  & \i[2646]  & \i[2645]  & new_n5406_ & ~new_n5416_ & new_n5408_;
  assign \o[23]  = ~new_n5969_ ^ new_n5970_;
  assign new_n5969_ = (~new_n5861_ & new_n5860_) | (new_n5859_ & (~new_n5861_ | new_n5860_));
  assign new_n5970_ = new_n5971_ ^ new_n5972_;
  assign new_n5971_ = (~new_n5863_ & new_n5967_) | (new_n5862_ & (~new_n5863_ | new_n5967_));
  assign new_n5972_ = ~new_n5973_ ^ new_n5974_;
  assign new_n5973_ = (~new_n5865_ & new_n5966_) | (new_n5864_ & (~new_n5865_ | new_n5966_));
  assign new_n5974_ = new_n5975_ ? (new_n5976_ ^ new_n6010_) : (~new_n5976_ ^ new_n6010_);
  assign new_n5975_ = (~new_n5881_ & new_n5965_) | (~new_n5866_ & (~new_n5881_ | new_n5965_));
  assign new_n5976_ = new_n5977_ ? (new_n5985_ ^ new_n5986_) : (~new_n5985_ ^ new_n5986_);
  assign new_n5977_ = new_n5978_ ? (~new_n5979_ ^ new_n5984_) : (new_n5979_ ^ new_n5984_);
  assign new_n5978_ = (~new_n5870_ & ~new_n5878_) | (new_n5869_ & (~new_n5870_ | ~new_n5878_));
  assign new_n5979_ = ~new_n5980_ ^ new_n5981_;
  assign new_n5980_ = (~new_n5873_ & new_n5872_) | (new_n5871_ & (~new_n5873_ | new_n5872_));
  assign new_n5981_ = new_n5982_ ^ new_n5983_;
  assign new_n5982_ = (new_n5960_ & new_n5961_) | (~new_n5955_ & (new_n5960_ | new_n5961_));
  assign new_n5983_ = (new_n5876_ & new_n5877_) | (~new_n5874_ & (new_n5876_ | new_n5877_));
  assign new_n5984_ = (~new_n5945_ & new_n5963_) | (new_n5944_ & (~new_n5945_ | new_n5963_));
  assign new_n5985_ = (~new_n5943_ & new_n5964_) | (~new_n5882_ & (~new_n5943_ | new_n5964_));
  assign new_n5986_ = new_n5987_ ? (new_n5988_ ^ new_n6006_) : (~new_n5988_ ^ new_n6006_);
  assign new_n5987_ = (~new_n5919_ & new_n5942_) | (~new_n5883_ & (~new_n5919_ | new_n5942_));
  assign new_n5988_ = new_n5989_ ? (new_n5992_ ^ new_n5993_) : (~new_n5992_ ^ new_n5993_);
  assign new_n5989_ = ~new_n5990_ ^ new_n5991_;
  assign new_n5990_ = (~new_n5890_ & ~new_n5899_) | (new_n5885_ & (~new_n5890_ | ~new_n5899_));
  assign new_n5991_ = (~new_n5927_ & ~new_n5936_) | (~new_n5922_ & (~new_n5927_ | ~new_n5936_));
  assign new_n5992_ = (~new_n5905_ & new_n5904_) | (~new_n5884_ & (~new_n5905_ | new_n5904_));
  assign new_n5993_ = new_n5994_ ^ new_n5995_;
  assign new_n5994_ = new_n5906_ & new_n5915_;
  assign new_n5995_ = new_n5996_ ? (new_n6003_ ^ new_n6004_) : (~new_n6003_ ^ new_n6004_);
  assign new_n5996_ = \i[1403]  ? new_n5997_ : (new_n3560_ ? new_n6002_ : ~new_n5510_);
  assign new_n5997_ = new_n3437_ ? new_n5998_ : ((~new_n6000_ | ~new_n3696_) & (new_n5515_ | ~new_n6001_ | new_n3696_));
  assign new_n5998_ = new_n5151_ ? new_n5999_ : (new_n5769_ ? ~new_n5591_ : ~\i[595] );
  assign new_n5999_ = new_n5518_ ? new_n4091_ : ~new_n3564_;
  assign new_n6000_ = ~new_n3523_ & new_n4199_;
  assign new_n6001_ = ~\i[1719]  & ~\i[1717]  & ~\i[1718] ;
  assign new_n6002_ = (new_n3697_ | new_n5512_ | new_n4470_) & (~new_n5507_ | ~new_n5098_ | ~new_n4470_);
  assign new_n6003_ = new_n5845_ & new_n5940_ & ~new_n5585_ & new_n5128_;
  assign new_n6004_ = new_n5566_ & new_n6005_ & new_n5569_ & ~new_n5571_ & ~\i[1623] ;
  assign new_n6005_ = ~\i[871]  & (~\i[870]  | (~\i[869]  & ~\i[868] ));
  assign new_n6006_ = new_n6007_ ? (new_n6008_ ^ new_n6009_) : (~new_n6008_ ^ new_n6009_);
  assign new_n6007_ = (~new_n5947_ & ~new_n5954_) | (new_n5946_ & (~new_n5947_ | ~new_n5954_));
  assign new_n6008_ = (~new_n5921_ & new_n5941_) | (new_n5920_ & (~new_n5921_ | new_n5941_));
  assign new_n6009_ = (~new_n5951_ & new_n5953_) | (~new_n5948_ & (~new_n5951_ | new_n5953_));
  assign new_n6010_ = (~new_n5868_ & new_n5880_) | (new_n5867_ & (~new_n5868_ | new_n5880_));
  assign \o[24]  = ((new_n6012_ | new_n6013_) & (~new_n6014_ ^ ~new_n6015_)) | (~new_n6012_ & ~new_n6013_ & (~new_n6014_ ^ new_n6015_));
  assign new_n6012_ = ~new_n5970_ & new_n5969_;
  assign new_n6013_ = ~new_n5972_ & new_n5971_;
  assign new_n6014_ = new_n5973_ & new_n5974_;
  assign new_n6015_ = ~new_n6016_ ^ new_n6017_;
  assign new_n6016_ = (~new_n5976_ & new_n6010_) | (new_n5975_ & (~new_n5976_ | new_n6010_));
  assign new_n6017_ = new_n6018_ ? (new_n6019_ ^ new_n6031_) : (~new_n6019_ ^ new_n6031_);
  assign new_n6018_ = (~new_n5986_ & new_n5985_) | (~new_n5977_ & (~new_n5986_ | new_n5985_));
  assign new_n6019_ = new_n6020_ ? (new_n6024_ ^ new_n6025_) : (~new_n6024_ ^ new_n6025_);
  assign new_n6020_ = new_n6021_ ? (new_n6022_ ^ new_n6023_) : (~new_n6022_ ^ new_n6023_);
  assign new_n6021_ = new_n5980_ & new_n5981_;
  assign new_n6022_ = (new_n6008_ & new_n6009_) | (new_n6007_ & (new_n6008_ | new_n6009_));
  assign new_n6023_ = new_n5982_ & new_n5983_;
  assign new_n6024_ = (~new_n5988_ & ~new_n6006_) | (new_n5987_ & (~new_n5988_ | ~new_n6006_));
  assign new_n6025_ = new_n6026_ ? (~new_n6027_ ^ new_n6030_) : (new_n6027_ ^ new_n6030_);
  assign new_n6026_ = (~new_n5993_ & new_n5992_) | (~new_n5989_ & (~new_n5993_ | new_n5992_));
  assign new_n6027_ = new_n6028_ ^ new_n6029_;
  assign new_n6028_ = ~new_n5994_ & new_n5995_;
  assign new_n6029_ = (new_n6003_ & new_n6004_) | (~new_n5996_ & (new_n6003_ | new_n6004_));
  assign new_n6030_ = new_n5990_ & new_n5991_;
  assign new_n6031_ = (~new_n5979_ & new_n5984_) | (new_n5978_ & (~new_n5979_ | new_n5984_));
  assign \o[25]  = ~new_n6033_ ^ new_n6034_;
  assign new_n6033_ = (new_n6014_ | (~new_n6015_ & (new_n6013_ | new_n6012_))) & (new_n6013_ | new_n6012_ | ~new_n6015_);
  assign new_n6034_ = new_n6035_ ^ new_n6036_;
  assign new_n6035_ = new_n6016_ & new_n6017_;
  assign new_n6036_ = ~new_n6037_ ^ new_n6038_;
  assign new_n6037_ = (~new_n6019_ & new_n6031_) | (new_n6018_ & (~new_n6019_ | new_n6031_));
  assign new_n6038_ = new_n6039_ ? (new_n6040_ ^ new_n6043_) : (~new_n6040_ ^ new_n6043_);
  assign new_n6039_ = (~new_n6025_ & new_n6024_) | (~new_n6020_ & (~new_n6025_ | new_n6024_));
  assign new_n6040_ = new_n6041_ ^ new_n6042_;
  assign new_n6041_ = (~new_n6027_ & new_n6030_) | (new_n6026_ & (~new_n6027_ | new_n6030_));
  assign new_n6042_ = ~new_n6028_ & ~new_n6029_;
  assign new_n6043_ = (new_n6022_ & new_n6023_) | (new_n6021_ & (new_n6022_ | new_n6023_));
  assign \o[26]  = ((~new_n6048_ ^ ~new_n6049_) & ((new_n6047_ & (new_n6045_ | new_n6046_)) | (~new_n6045_ & ~new_n6046_ & ~new_n6047_))) | ((~new_n6048_ ^ new_n6049_) & ((~new_n6045_ & ~new_n6046_ & new_n6047_) | (~new_n6047_ & (new_n6045_ | new_n6046_))));
  assign new_n6045_ = ~new_n6034_ & new_n6033_;
  assign new_n6046_ = ~new_n6036_ & new_n6035_;
  assign new_n6047_ = new_n6037_ & new_n6038_;
  assign new_n6048_ = (~new_n6040_ & new_n6043_) | (new_n6039_ & (~new_n6040_ | new_n6043_));
  assign new_n6049_ = ~new_n6042_ & new_n6041_;
  assign \o[27]  = (~new_n6047_ | ~new_n6048_ | ~new_n6049_ | (~new_n6045_ & ~new_n6046_)) & (new_n6047_ | new_n6048_ | new_n6049_) & (new_n6045_ | new_n6046_ | ((new_n6048_ | new_n6049_) & (new_n6047_ | (new_n6048_ & new_n6049_))));
  assign \o[28]  = new_n6052_ ^ new_n6462_;
  assign new_n6052_ = new_n6053_ ? (~new_n6367_ ^ new_n6448_) : (new_n6367_ ^ new_n6448_);
  assign new_n6053_ = new_n6054_ ? (~new_n6183_ ^ new_n6349_) : (new_n6183_ ^ new_n6349_);
  assign new_n6054_ = new_n6055_ ? (new_n6156_ ^ new_n6173_) : (~new_n6156_ ^ new_n6173_);
  assign new_n6055_ = new_n6056_ ? (new_n6105_ ^ new_n6148_) : (~new_n6105_ ^ new_n6148_);
  assign new_n6056_ = new_n6057_ ? (new_n6075_ ^ new_n6088_) : (~new_n6075_ ^ new_n6088_);
  assign new_n6057_ = (new_n6070_ | new_n6058_ | ~new_n4150_) & (new_n4150_ | (new_n6065_ ? ~new_n6066_ : ~new_n6063_));
  assign new_n6058_ = new_n6061_ & (new_n6059_ | (~new_n6062_ & new_n5134_ & new_n4392_));
  assign new_n6059_ = new_n6060_ & (~\i[639]  | (~\i[638]  & (~\i[637]  | ~\i[636] )));
  assign new_n6060_ = ~new_n4392_ & ~\i[2099]  & (~\i[2098]  | (~\i[2096]  & ~\i[2097] ));
  assign new_n6061_ = \i[855]  & (\i[853]  | \i[854]  | \i[852] );
  assign new_n6062_ = ~\i[1971]  & ~\i[1969]  & ~\i[1970] ;
  assign new_n6063_ = ~new_n6064_ & (new_n3741_ | new_n5558_ | ~\i[1273]  | ~\i[1274]  | ~\i[1275] );
  assign new_n6064_ = new_n5558_ & (new_n5035_ ? ~new_n3459_ : (\i[723]  | (\i[721]  & \i[722] )));
  assign new_n6065_ = \i[733]  & new_n4414_ & \i[732] ;
  assign new_n6066_ = (~new_n3788_ | new_n4061_ | ~new_n3750_) & (new_n3750_ | (new_n6068_ ? new_n6069_ : new_n6067_));
  assign new_n6067_ = ~\i[2855]  & (~\i[2854]  | (~\i[2853]  & ~\i[2852] ));
  assign new_n6068_ = \i[854]  & \i[855] ;
  assign new_n6069_ = \i[1867]  & \i[1866]  & \i[1864]  & \i[1865] ;
  assign new_n6070_ = ~new_n6061_ & ((~new_n6074_ & new_n6073_ & ~new_n3592_) | (~new_n6071_ & new_n6072_ & new_n3592_));
  assign new_n6071_ = \i[751]  & (\i[750]  | (\i[749]  & \i[748] ));
  assign new_n6072_ = ~\i[1534]  & ~\i[1535]  & (~\i[1533]  | ~\i[1532] );
  assign new_n6073_ = ~\i[2070]  & ~\i[2071]  & (~\i[2069]  | ~\i[2068] );
  assign new_n6074_ = ~\i[835]  & ~\i[833]  & ~\i[834] ;
  assign new_n6075_ = (~new_n6086_ | ~new_n6087_ | ~new_n4070_) & (new_n6076_ | new_n6082_ | new_n4070_);
  assign new_n6076_ = new_n4266_ & ~new_n6077_ & ~new_n6079_;
  assign new_n6077_ = ~new_n6078_ & (~\i[2859]  | (~\i[2858]  & (~\i[2857]  | ~\i[2856] )));
  assign new_n6078_ = (~\i[963]  & ~\i[962]  & ~new_n4684_) | (\i[1763]  & new_n4684_ & (\i[1762]  | \i[1761] ));
  assign new_n6079_ = new_n6080_ & \i[2859]  & (\i[2858]  | (\i[2856]  & \i[2857] ));
  assign new_n6080_ = ~\i[946]  & ~\i[947]  & new_n6081_ & (~\i[945]  | ~\i[944] );
  assign new_n6081_ = \i[1391]  & \i[1390]  & \i[1388]  & \i[1389] ;
  assign new_n6082_ = ~new_n6083_ & ~new_n4266_ & (new_n5476_ | \i[845]  | ~new_n6085_ | ~new_n6084_);
  assign new_n6083_ = new_n3781_ & ~new_n6084_ & new_n3302_;
  assign new_n6084_ = \i[1067]  & (\i[1066]  | (\i[1065]  & \i[1064] ));
  assign new_n6085_ = ~\i[846]  & ~\i[847] ;
  assign new_n6086_ = new_n5836_ & ((~\i[2429]  & ~\i[2428] ) | ~\i[2431]  | ~\i[2430] );
  assign new_n6087_ = \i[2762]  & \i[2763] ;
  assign new_n6088_ = (\i[1391]  & (\i[1390]  | (\i[1388]  & \i[1389] ))) ? new_n6089_ : new_n6095_;
  assign new_n6089_ = new_n6094_ ? (new_n6093_ ? new_n6091_ : ~new_n6092_) : ~new_n6090_;
  assign new_n6090_ = \i[1943]  & \i[1942]  & \i[1941]  & new_n4244_ & \i[1940] ;
  assign new_n6091_ = new_n3683_ & (\i[979]  | \i[978] );
  assign new_n6092_ = \i[2655]  & (\i[2654]  | (\i[2653]  & \i[2652] ));
  assign new_n6093_ = ~\i[922]  & ~\i[923]  & (~\i[921]  | ~\i[920] );
  assign new_n6094_ = ~\i[519]  & (~\i[518]  | (~\i[517]  & ~\i[516] ));
  assign new_n6095_ = (new_n6103_ | new_n6099_ | ~\i[1271]  | (~\i[1269]  & ~\i[1270] )) & (new_n6096_ | (\i[1271]  & (\i[1269]  | \i[1270] )));
  assign new_n6096_ = new_n5052_ ? new_n6097_ : (new_n4214_ ? new_n3446_ : \i[2407] );
  assign new_n6097_ = (~\i[943]  | ~new_n4361_ | (~\i[942]  & (~\i[940]  | ~\i[941] ))) & (new_n6098_ | new_n4361_);
  assign new_n6098_ = ~\i[986]  & ~\i[987]  & (~\i[985]  | ~\i[984] );
  assign new_n6099_ = new_n3550_ & ((~\i[724]  & new_n6100_ & (\i[371]  | new_n6102_)) | (~\i[1055]  & (\i[724]  | ~new_n6100_)));
  assign new_n6100_ = ~\i[725]  & new_n6101_;
  assign new_n6101_ = ~\i[726]  & ~\i[727] ;
  assign new_n6102_ = \i[370]  & (\i[369]  | \i[368] );
  assign new_n6103_ = ~\i[1663]  & ~\i[1662]  & ~\i[1661]  & ~new_n3550_ & ~new_n6104_;
  assign new_n6104_ = \i[1590]  & \i[1591]  & (\i[1589]  | \i[1588] );
  assign new_n6105_ = new_n6106_ ? (~new_n6123_ ^ new_n6133_) : (new_n6123_ ^ new_n6133_);
  assign new_n6106_ = (~\i[1495]  & (~\i[1494]  | (~\i[1492]  & ~\i[1493] ))) ? new_n6107_ : new_n6112_;
  assign new_n6107_ = ~new_n6108_ & (~new_n6111_ | (~new_n5527_ & new_n3299_ & new_n3350_));
  assign new_n6108_ = ~\i[1601]  & new_n5039_ & (new_n4674_ ? (~\i[2283]  | new_n6110_) : new_n6109_);
  assign new_n6109_ = new_n4214_ ? new_n5584_ : new_n3312_;
  assign new_n6110_ = \i[947]  & \i[946]  & \i[944]  & \i[945] ;
  assign new_n6111_ = (\i[1601]  | ~new_n5039_) & (new_n3350_ | \i[2082]  | \i[2083]  | ~new_n4334_);
  assign new_n6112_ = new_n3893_ ? new_n6113_ : (new_n6121_ | (~new_n6118_ & new_n4378_));
  assign new_n6113_ = ~new_n6114_ & (~new_n4330_ | (~new_n6117_ & new_n6115_) | (~new_n6116_ & \i[863]  & ~new_n6115_));
  assign new_n6114_ = ~new_n4330_ & \i[1595]  & (\i[1594]  | (\i[1592]  & \i[1593] ));
  assign new_n6115_ = \i[1191]  & (\i[1189]  | \i[1190]  | \i[1188] );
  assign new_n6116_ = ~\i[862]  & (~\i[861]  | ~\i[860] );
  assign new_n6117_ = ~\i[1059]  & (~\i[1058]  | (~\i[1057]  & ~\i[1056] ));
  assign new_n6118_ = \i[1411]  ? new_n6120_ : new_n6119_;
  assign new_n6119_ = new_n4932_ & ~\i[1166]  & ~\i[1167] ;
  assign new_n6120_ = ~\i[2287]  & (~\i[2285]  | ~\i[2286]  | ~\i[2284] );
  assign new_n6121_ = ~new_n6122_ & ~new_n4378_ & \i[739]  & (\i[738]  | \i[737]  | \i[736] );
  assign new_n6122_ = ~\i[947]  & (~\i[946]  | (~\i[945]  & ~\i[944] ));
  assign new_n6123_ = new_n6131_ ? new_n6124_ : (~new_n6132_ | (~new_n3556_ & ~new_n4273_));
  assign new_n6124_ = new_n6128_ ? new_n6125_ : ((new_n6129_ | new_n6130_ | ~new_n4467_) & (~new_n4870_ | new_n4467_));
  assign new_n6125_ = (new_n6126_ | \i[2848]  | \i[2849]  | ~new_n5624_) & (~new_n4235_ | ~new_n6127_ | (~\i[2848]  & ~\i[2849]  & new_n5624_));
  assign new_n6126_ = (new_n4000_ | ~new_n6067_) & (\i[839]  | new_n6067_ | (\i[838]  & (\i[836]  | \i[837] )));
  assign new_n6127_ = ~\i[955]  & ~\i[954]  & ~\i[952]  & ~\i[953] ;
  assign new_n6128_ = ~\i[2283]  & (~\i[2281]  | ~\i[2282]  | ~\i[2280] );
  assign new_n6129_ = ~\i[859]  & (~\i[857]  | ~\i[858]  | ~\i[856] );
  assign new_n6130_ = \i[851]  & (\i[849]  | \i[850]  | \i[848] );
  assign new_n6131_ = new_n4031_ & ~\i[764]  & ~\i[765] ;
  assign new_n6132_ = new_n4947_ & (~\i[857]  | ~\i[856] );
  assign new_n6133_ = (new_n6144_ | new_n6141_ | new_n6147_) & (~new_n6147_ | (~new_n6137_ & (~new_n4412_ | new_n6134_)));
  assign new_n6134_ = new_n6135_ ? (new_n6136_ ? new_n5703_ : new_n4017_) : ~new_n4028_;
  assign new_n6135_ = ~\i[875]  & ~\i[873]  & ~\i[874] ;
  assign new_n6136_ = ~\i[1423]  & (~\i[1421]  | ~\i[1422]  | ~\i[1420] );
  assign new_n6137_ = ~new_n4412_ & (new_n5822_ ? ~new_n6140_ : (new_n6138_ ? new_n6139_ : ~new_n3582_));
  assign new_n6138_ = \i[1971]  & (\i[1969]  | \i[1970]  | \i[1968] );
  assign new_n6139_ = ~\i[983]  & (~\i[982]  | (~\i[981]  & ~\i[980] ));
  assign new_n6140_ = \i[851]  & (\i[849]  | \i[850] ) & (\i[867]  | (\i[865]  & \i[866] ));
  assign new_n6141_ = ~new_n3278_ & (new_n6142_ | (~new_n3584_ & ~new_n5533_ & new_n3476_));
  assign new_n6142_ = ~new_n3476_ & (new_n6143_ ? (~\i[1875]  | ~\i[1874] ) : ~new_n4920_);
  assign new_n6143_ = \i[855]  & (\i[854]  | \i[853] );
  assign new_n6144_ = new_n3278_ & (new_n6146_ ? new_n6145_ : (new_n3499_ ? ~new_n5431_ : ~new_n5836_));
  assign new_n6145_ = new_n4681_ & (\i[2187]  | (\i[2185]  & \i[2186] ));
  assign new_n6146_ = ~\i[2091]  & (~\i[2089]  | ~\i[2090]  | ~\i[2088] );
  assign new_n6147_ = \i[1599]  & (\i[1597]  | \i[1598]  | \i[1596] );
  assign new_n6148_ = ~\i[2967]  & (~\i[2965]  | ~\i[2966]  | ~\i[2964] ) & (new_n6152_ | new_n6149_);
  assign new_n6149_ = \i[747]  & (new_n4695_ ? (new_n3988_ ? ~new_n4895_ : ~new_n5678_) : ~new_n6150_);
  assign new_n6150_ = (new_n5684_ | new_n6151_) & (\i[971]  | ~new_n6151_ | (\i[970]  & (\i[968]  | \i[969] )));
  assign new_n6151_ = \i[1075]  & (\i[1073]  | \i[1074]  | \i[1072] );
  assign new_n6152_ = ~\i[747]  & (new_n6155_ ? (new_n5802_ ? ~new_n3495_ : ~new_n4895_) : ~new_n6153_);
  assign new_n6153_ = ~new_n6154_ & \i[839]  & (\i[838]  | \i[837]  | \i[836] );
  assign new_n6154_ = ~\i[962]  & ~\i[963]  & (~\i[961]  | ~\i[960] );
  assign new_n6155_ = new_n6085_ & ~\i[844]  & ~\i[845] ;
  assign new_n6156_ = new_n6171_ ? (new_n6172_ ? ~new_n6165_ : new_n6169_) : new_n6157_;
  assign new_n6157_ = new_n6164_ ? (new_n6162_ | (~new_n6158_ & new_n3750_)) : ~new_n6161_;
  assign new_n6158_ = ~new_n6159_ & (~new_n6160_ | new_n4379_);
  assign new_n6159_ = ~new_n6160_ & (~\i[729]  | ~\i[730]  | ~\i[731] );
  assign new_n6160_ = ~\i[1987]  & (~\i[1986]  | ~\i[1985] );
  assign new_n6161_ = (\i[954]  | \i[955]  | ~new_n5665_) & (new_n4029_ | ~new_n4342_ | new_n5665_);
  assign new_n6162_ = ~new_n3750_ & ((~new_n3687_ & new_n6163_) | (~\i[2417]  & ~\i[2418]  & ~\i[2419]  & ~new_n6163_));
  assign new_n6163_ = \i[859]  & (\i[858]  | (\i[857]  & \i[856] ));
  assign new_n6164_ = \i[739]  & (\i[738]  | (\i[737]  & \i[736] ));
  assign new_n6165_ = (~new_n6167_ | ~new_n6168_ | ~new_n5577_) & (new_n3427_ | new_n6166_ | new_n5577_);
  assign new_n6166_ = ~\i[1163]  & (~\i[1161]  | ~\i[1162]  | ~\i[1160] );
  assign new_n6167_ = ~\i[1535]  & (~\i[1534]  | (~\i[1533]  & ~\i[1532] ));
  assign new_n6168_ = \i[2055]  & \i[2054]  & \i[2052]  & \i[2053] ;
  assign new_n6169_ = new_n6170_ & ((~\i[2185]  & ~\i[2184] ) | ~\i[2187]  | ~\i[2186] );
  assign new_n6170_ = ~\i[767]  & (~\i[2862]  | ~\i[2863] ) & (~\i[766]  | (~\i[765]  & ~\i[764] ));
  assign new_n6171_ = new_n5078_ & (~\i[2077]  | ~\i[2076] );
  assign new_n6172_ = ~\i[2523]  & (~\i[2521]  | ~\i[2522]  | ~\i[2520] );
  assign new_n6173_ = new_n3761_ ? new_n6174_ : new_n6179_;
  assign new_n6174_ = new_n3221_ ? (new_n4861_ | (~new_n6178_ & new_n5533_)) : new_n6175_;
  assign new_n6175_ = ~new_n6176_ & (\i[837]  | \i[838]  | \i[839]  | ~new_n4245_);
  assign new_n6176_ = new_n6177_ & ((~\i[1170]  & ~\i[1171] ) ? ~new_n4061_ : new_n6101_);
  assign new_n6177_ = \i[839]  & (\i[838]  | \i[837] );
  assign new_n6178_ = \i[1927]  & (\i[1926]  | (\i[1925]  & \i[1924] ));
  assign new_n6179_ = (new_n3799_ | ~\i[1553]  | ~\i[1554]  | ~\i[1555] ) & (new_n6182_ | ~new_n6180_ | (\i[1553]  & \i[1554]  & \i[1555] ));
  assign new_n6180_ = \i[2267]  & new_n4031_ & ~\i[2207]  & new_n6181_;
  assign new_n6181_ = (\i[2265]  | \i[2266] ) & (~\i[2205]  | ~\i[2206] );
  assign new_n6182_ = \i[765]  & new_n4031_ & \i[764] ;
  assign new_n6183_ = new_n6184_ ? (~new_n6269_ ^ new_n6333_) : (new_n6269_ ^ new_n6333_);
  assign new_n6184_ = new_n6185_ ? (new_n6226_ ^ new_n6268_) : (~new_n6226_ ^ new_n6268_);
  assign new_n6185_ = new_n6186_ ? (~new_n6199_ ^ new_n6216_) : (new_n6199_ ^ new_n6216_);
  assign new_n6186_ = ~new_n6187_ & (~new_n6193_ | (new_n4285_ & (new_n5005_ ? ~new_n6197_ : new_n6198_)));
  assign new_n6187_ = ~new_n4682_ & (new_n6188_ | (\i[1395]  & (new_n3450_ ? new_n6190_ : new_n6192_)));
  assign new_n6188_ = ~\i[1395]  & new_n4470_ & (new_n5703_ ? ~new_n6189_ : ~new_n4061_);
  assign new_n6189_ = \i[1870]  & \i[1871]  & (\i[1869]  | \i[1868] );
  assign new_n6190_ = (new_n6191_ | (~\i[1834]  & ~\i[1835] )) & (~\i[753]  | ~\i[754]  | ~\i[755]  | \i[1834]  | \i[1835] );
  assign new_n6191_ = ~\i[1867]  & (~\i[1865]  | ~\i[1866]  | ~\i[1864] );
  assign new_n6192_ = \i[395]  & (~\i[1288]  | ~\i[1289]  | ~\i[1290]  | ~\i[1291] );
  assign new_n6193_ = new_n4682_ & (new_n4285_ | ((new_n6195_ | new_n6196_) & (~new_n6194_ | ~new_n4659_ | ~new_n6196_)));
  assign new_n6194_ = new_n4521_ & (~\i[1721]  | ~\i[1720] );
  assign new_n6195_ = (~\i[2746]  | ~\i[2747] ) & (~\i[1926]  | ~\i[1927]  | ~\i[1924]  | ~\i[1925] );
  assign new_n6196_ = \i[1599]  & (\i[1598]  | (\i[1597]  & \i[1596] ));
  assign new_n6197_ = new_n3576_ ? (~\i[927]  | (~\i[925]  & ~\i[926] )) : ~new_n4357_;
  assign new_n6198_ = ~\i[759]  & ~\i[758]  & ~\i[756]  & ~\i[757] ;
  assign new_n6199_ = ~new_n6207_ & (~new_n6212_ | ((~new_n6200_ | ~new_n3683_) & (new_n6205_ | new_n6213_ | new_n3683_)));
  assign new_n6200_ = (new_n6201_ | new_n6204_) & (new_n4167_ | new_n4684_ | ~new_n6204_);
  assign new_n6201_ = new_n6203_ ? (~\i[1887]  | (~\i[1885]  & ~\i[1886] )) : ~new_n6202_;
  assign new_n6202_ = ~\i[723]  & ~\i[721]  & ~\i[722] ;
  assign new_n6203_ = \i[1067]  & (\i[1066]  | \i[1065] );
  assign new_n6204_ = \i[1822]  & \i[1823]  & (\i[1821]  | \i[1820] );
  assign new_n6205_ = ~new_n6206_ & (new_n4336_ | ~new_n4019_) & (\i[1553]  | \i[1554]  | \i[1555]  | new_n4019_);
  assign new_n6206_ = ~\i[2323]  & ~\i[2321]  & ~\i[2322] ;
  assign new_n6207_ = ~new_n6212_ & (new_n3800_ ? new_n6210_ : (new_n4056_ ? new_n6208_ : new_n6209_));
  assign new_n6208_ = (new_n5449_ | ~new_n6069_) & (~\i[1382]  | ~\i[1383]  | new_n6069_ | (~\i[1381]  & ~\i[1380] ));
  assign new_n6209_ = \i[2627]  ? (~new_n4225_ & (\i[2626]  | \i[2624]  | \i[2625] )) : (new_n4225_ & (~\i[2626]  | (~\i[2624]  & ~\i[2625] )));
  assign new_n6210_ = (~new_n4428_ | (new_n5802_ ? new_n6001_ : ~new_n4002_)) & (~new_n4994_ | ~new_n6211_ | new_n4428_);
  assign new_n6211_ = \i[1598]  & \i[1599]  & (\i[1597]  | \i[1596] );
  assign new_n6212_ = \i[1747]  & \i[1746]  & \i[1744]  & \i[1745] ;
  assign new_n6213_ = new_n6206_ & (\i[859]  ? new_n6214_ : (~\i[635]  | new_n6215_));
  assign new_n6214_ = \i[1191]  & (\i[1190]  | (\i[1189]  & \i[1188] ));
  assign new_n6215_ = ~\i[634]  & (~\i[633]  | ~\i[632] );
  assign new_n6216_ = new_n6225_ ? (new_n6224_ | (new_n6223_ & new_n4820_ & new_n5588_)) : new_n6217_;
  assign new_n6217_ = (new_n6218_ | ~new_n6221_) & (new_n6220_ | ~new_n6222_ | new_n6221_);
  assign new_n6218_ = (~new_n6219_ | ~new_n4446_ | ~new_n3309_) & (new_n3309_ | (new_n3220_ & (~\i[998]  | ~\i[999] )));
  assign new_n6219_ = ~\i[1959]  & (~\i[1957]  | ~\i[1958]  | ~\i[1956] );
  assign new_n6220_ = (~new_n3313_ | ~new_n3988_) & (~\i[1316]  | ~\i[1317]  | ~\i[1318]  | ~\i[1319]  | new_n3988_);
  assign new_n6221_ = ~\i[747]  & ~\i[746]  & ~\i[744]  & ~\i[745] ;
  assign new_n6222_ = ~\i[1671]  & ~\i[1669]  & ~\i[1670] ;
  assign new_n6223_ = (~new_n4977_ | new_n5810_) & (\i[2962]  | \i[2963]  | ~new_n5810_ | (\i[2961]  & \i[2960] ));
  assign new_n6224_ = ~new_n5588_ & (~new_n3990_ | ~new_n3244_) & (~\i[277]  | ~\i[278]  | ~\i[279] );
  assign new_n6225_ = ~\i[2499]  & ~\i[2498]  & ~\i[2496]  & ~\i[2497] ;
  assign new_n6226_ = new_n6227_ ? (~new_n6244_ ^ new_n6255_) : (new_n6244_ ^ new_n6255_);
  assign new_n6227_ = (new_n6228_ | ~new_n6155_) & (new_n6239_ | new_n6242_ | new_n6155_);
  assign new_n6228_ = (new_n6229_ | ~new_n5066_) & (new_n3399_ | new_n6236_ | new_n5066_ | (~new_n6238_ & new_n6237_));
  assign new_n6229_ = new_n4837_ ? (new_n6233_ ? new_n6235_ : ~new_n6234_) : new_n6230_;
  assign new_n6230_ = new_n6231_ ? new_n5022_ : ~new_n6232_;
  assign new_n6231_ = ~\i[2207]  & ~\i[2206]  & ~\i[2204]  & ~\i[2205] ;
  assign new_n6232_ = \i[1974]  & \i[1975]  & (\i[1973]  | \i[1972] );
  assign new_n6233_ = \i[1706]  & \i[1707]  & (\i[1705]  | \i[1704] );
  assign new_n6234_ = \i[1503]  & (\i[1501]  | \i[1502]  | \i[1500] );
  assign new_n6235_ = ~\i[1834]  & ~\i[1835]  & (~\i[1833]  | ~\i[1832] );
  assign new_n6236_ = ~new_n6237_ & ~\i[2271]  & (~\i[2270]  | (~\i[2268]  & ~\i[2269] ));
  assign new_n6237_ = ~\i[651]  & ~\i[650]  & ~\i[648]  & ~\i[649] ;
  assign new_n6238_ = ~\i[2415]  & ~\i[2414]  & ~\i[2412]  & ~\i[2413] ;
  assign new_n6239_ = new_n5743_ & (new_n3775_ | (new_n6241_ & ~new_n6240_) | (new_n3269_ & new_n6240_));
  assign new_n6240_ = new_n3540_ & ~\i[848]  & ~\i[849] ;
  assign new_n6241_ = ~\i[2818]  & ~\i[2819]  & (~\i[2817]  | ~\i[2816] );
  assign new_n6242_ = ~new_n5743_ & ((~new_n5616_ & ~new_n6243_ & new_n4019_) | (~new_n4019_ & (~new_n4069_ | ~new_n6240_)));
  assign new_n6243_ = ~\i[2403]  & ~\i[2402]  & ~\i[2400]  & ~\i[2401] ;
  assign new_n6244_ = (new_n6248_ | ~new_n6254_) & (new_n6245_ | new_n6253_ | new_n6254_);
  assign new_n6245_ = (new_n6246_ | new_n5025_) & (~new_n4734_ | ~new_n4143_ | ~new_n5025_);
  assign new_n6246_ = (~new_n6247_ | ~new_n3613_) & (~\i[879]  | new_n3613_ | (~\i[878]  & (~\i[876]  | ~\i[877] )));
  assign new_n6247_ = ~\i[2731]  & new_n4407_;
  assign new_n6248_ = new_n5636_ ? new_n6249_ : ((new_n3628_ | new_n6127_) & (~new_n5808_ | ~\i[731]  | ~new_n6127_));
  assign new_n6249_ = (new_n6250_ | ~\i[1635]  | (~\i[1633]  & ~\i[1634] )) & (new_n6251_ | ~new_n6252_ | (\i[1635]  & (\i[1633]  | \i[1634] )));
  assign new_n6250_ = ~\i[1499]  & \i[1867]  & (~\i[1498]  | (~\i[1497]  & ~\i[1496] ));
  assign new_n6251_ = \i[1871]  & (\i[1869]  | \i[1870]  | \i[1868] );
  assign new_n6252_ = \i[1631]  & \i[1629]  & \i[1630] ;
  assign new_n6253_ = ~\i[1059]  & (~\i[1057]  | ~\i[1058]  | ~\i[1056] );
  assign new_n6254_ = ~\i[615]  & ~\i[613]  & ~\i[614] ;
  assign new_n6255_ = new_n6267_ ? new_n6258_ : ((new_n6256_ & new_n5079_) | (~new_n6262_ & ~new_n6265_ & ~new_n5079_));
  assign new_n6256_ = new_n3413_ ? (new_n4818_ ? ~new_n6257_ : ~new_n4002_) : \i[1391] ;
  assign new_n6257_ = ~\i[738]  & ~\i[739]  & (~\i[737]  | ~\i[736] );
  assign new_n6258_ = (new_n5843_ | new_n6260_ | new_n6238_) & (new_n6259_ | new_n6261_ | ~new_n6238_);
  assign new_n6259_ = (new_n3525_ | ~new_n4246_) & (\i[741]  | \i[742]  | \i[743]  | new_n4246_);
  assign new_n6260_ = new_n3285_ ? \i[1067]  : \i[2639] ;
  assign new_n6261_ = ~\i[1747]  & (~\i[1746]  | (~\i[1745]  & ~\i[1744] ));
  assign new_n6262_ = ~\i[769]  & ~\i[770]  & ~\i[771]  & (new_n6263_ ? new_n4172_ : ~new_n6264_);
  assign new_n6263_ = \i[1607]  & \i[1606]  & \i[1604]  & \i[1605] ;
  assign new_n6264_ = ~\i[1778]  & ~\i[1779]  & (~\i[1777]  | ~\i[1776] );
  assign new_n6265_ = (~new_n4810_ | new_n5035_) & (new_n6266_ | ~new_n5035_) & (\i[769]  | \i[770]  | \i[771] );
  assign new_n6266_ = ~\i[859]  & ~\i[857]  & ~\i[858] ;
  assign new_n6267_ = ~\i[1859]  & (~\i[1858]  | ~\i[1857] );
  assign new_n6268_ = new_n3221_ & new_n3761_ & ((new_n6178_ & ~new_n4861_) | (new_n5035_ & new_n3227_ & new_n4861_));
  assign new_n6269_ = new_n6270_ ? (new_n6321_ ^ new_n6268_) : (~new_n6321_ ^ new_n6268_);
  assign new_n6270_ = new_n6271_ ? (~new_n6293_ ^ new_n6309_) : (new_n6293_ ^ new_n6309_);
  assign new_n6271_ = new_n5675_ ? (new_n6203_ ? new_n6283_ : new_n6290_) : new_n6272_;
  assign new_n6272_ = new_n4946_ ? ((new_n6277_ | ~new_n3377_) & (new_n6279_ | new_n6282_ | new_n3377_)) : new_n6273_;
  assign new_n6273_ = new_n6276_ ? (new_n4831_ ? ~new_n4338_ : ~new_n6275_) : new_n6274_;
  assign new_n6274_ = ~new_n6214_ & \i[747]  & (\i[746]  | (\i[744]  & \i[745] ));
  assign new_n6275_ = ~\i[731]  & (~\i[729]  | ~\i[730]  | ~\i[728] );
  assign new_n6276_ = ~\i[1874]  & ~\i[1875]  & (~\i[1873]  | ~\i[1872] );
  assign new_n6277_ = (\i[519]  & (\i[517]  | \i[518] )) ? ~new_n6278_ : new_n4310_;
  assign new_n6278_ = ~\i[2291]  & ~\i[2290]  & ~\i[2288]  & ~\i[2289] ;
  assign new_n6279_ = ~new_n6281_ & new_n6280_;
  assign new_n6280_ = ~\i[2059]  & (~\i[2058]  | ~\i[2057] );
  assign new_n6281_ = \i[1718]  & \i[1719]  & (\i[1717]  | \i[1716] );
  assign new_n6282_ = ~new_n6280_ & (~\i[1639]  | (~\i[1637]  & ~\i[1638] ));
  assign new_n6283_ = new_n6287_ ? new_n6284_ : (new_n6289_ ? new_n6288_ : new_n4837_);
  assign new_n6284_ = (~new_n6286_ & ~new_n6285_) | (new_n4342_ & new_n6285_ & (\i[841]  | \i[840] ));
  assign new_n6285_ = ~\i[1079]  & (~\i[1077]  | ~\i[1078]  | ~\i[1076] );
  assign new_n6286_ = ~\i[1059]  & ~\i[1057]  & ~\i[1058] ;
  assign new_n6287_ = \i[1507]  & (\i[1505]  | \i[1506]  | \i[1504] );
  assign new_n6288_ = ~\i[1543]  & ~\i[1542]  & ~\i[1540]  & ~\i[1541] ;
  assign new_n6289_ = ~\i[1711]  & (~\i[1710]  | ~\i[1709] );
  assign new_n6290_ = ~new_n6291_ & (~new_n4471_ | (~new_n6292_ & ~new_n4246_) | (new_n5742_ & new_n4246_));
  assign new_n6291_ = ~new_n4471_ & ((\i[1178]  & \i[1179]  & (\i[607]  | \i[606] )) | (~new_n4379_ & (~\i[1178]  | ~\i[1179] )));
  assign new_n6292_ = \i[1727]  & \i[1726]  & \i[1724]  & \i[1725] ;
  assign new_n6293_ = new_n4190_ ? (new_n6308_ ? ~new_n6294_ : ~new_n6298_) : new_n6303_;
  assign new_n6294_ = new_n6297_ ? new_n6295_ : ~new_n6221_;
  assign new_n6295_ = new_n6296_ ? ~new_n3229_ : (\i[1423]  | (\i[1421]  & \i[1422] ));
  assign new_n6296_ = ~\i[1638]  & ~\i[1639]  & (~\i[1637]  | ~\i[1636] );
  assign new_n6297_ = ~\i[1079]  & ~\i[1077]  & ~\i[1078] ;
  assign new_n6298_ = (~new_n5039_ | ~\i[1511]  | new_n6302_) & (new_n6299_ | new_n6301_ | ~new_n6302_);
  assign new_n6299_ = ~\i[1755]  & new_n6300_ & \i[1541]  & (~\i[1754]  | ~\i[1753]  | ~\i[1752] );
  assign new_n6300_ = \i[1542]  & \i[1543] ;
  assign new_n6301_ = new_n3378_ & (~\i[1541]  | ~new_n6300_);
  assign new_n6302_ = ~\i[1519]  & (~\i[1518]  | ~\i[1517] );
  assign new_n6303_ = new_n5544_ ? ((~new_n6304_ & new_n4667_) | (~new_n6243_ & new_n4068_ & ~new_n4667_)) : new_n6305_;
  assign new_n6304_ = (new_n3726_ & ~new_n5683_) | (~\i[2176]  & ~\i[2177]  & new_n5494_ & new_n5683_);
  assign new_n6305_ = (~new_n6307_ & ~\i[2980]  & ~\i[2981]  & ~\i[2982]  & ~\i[2983] ) | (~new_n6306_ & (\i[2980]  | \i[2981]  | \i[2982]  | \i[2983] ));
  assign new_n6306_ = ~\i[2647]  & ~\i[2645]  & ~\i[2646] ;
  assign new_n6307_ = ~\i[391]  & ~\i[390]  & ~\i[388]  & ~\i[389] ;
  assign new_n6308_ = \i[1646]  & \i[1647]  & (\i[1645]  | \i[1644] );
  assign new_n6309_ = (new_n6315_ | ~new_n6132_ | new_n6131_) & (~new_n6131_ | (~new_n6312_ & (~new_n6319_ | new_n6310_)));
  assign new_n6310_ = ~new_n4017_ & (new_n6311_ ? \i[523]  : ~new_n4048_);
  assign new_n6311_ = ~\i[743]  & (~\i[742]  | (~\i[741]  & ~\i[740] ));
  assign new_n6312_ = ~new_n3666_ & (~new_n6313_ | new_n5674_ | ~new_n5421_) & (new_n5440_ | ~new_n6314_ | new_n5421_);
  assign new_n6313_ = ~\i[1323]  & ~\i[1322]  & ~\i[1320]  & ~\i[1321] ;
  assign new_n6314_ = ~\i[995]  & (~\i[993]  | ~\i[994]  | ~\i[992] );
  assign new_n6315_ = (~new_n6316_ | new_n6317_) & (new_n6318_ | ~new_n6317_ | (new_n4080_ & (\i[1190]  | \i[1191] )));
  assign new_n6316_ = ~\i[879]  & ~\i[877]  & ~\i[878] ;
  assign new_n6317_ = ~\i[643]  & ~\i[641]  & ~\i[642] ;
  assign new_n6318_ = ~\i[1190]  & ~\i[1191]  & ((~\i[620]  & ~\i[621] ) | ~\i[623]  | ~\i[622] );
  assign new_n6319_ = new_n3666_ & (new_n4723_ | ~new_n4017_ | ~new_n6320_);
  assign new_n6320_ = \i[975]  & (\i[974]  | (\i[973]  & \i[972] ));
  assign new_n6321_ = ~new_n6322_ & (\i[1646]  | \i[1647]  | (new_n4190_ ? new_n6329_ : new_n6326_));
  assign new_n6322_ = (new_n6323_ | ~new_n3710_) & (\i[1647]  | \i[1646] ) & (new_n4863_ | new_n4331_ | new_n3710_);
  assign new_n6323_ = (~new_n6324_ | new_n6325_ | ~new_n4470_) & (new_n4470_ | (new_n3518_ ? new_n4740_ : new_n4673_));
  assign new_n6324_ = ~\i[1819]  & (~\i[1818]  | (~\i[1817]  & ~\i[1816] ));
  assign new_n6325_ = \i[2434]  & \i[2435]  & (\i[2433]  | \i[2432] );
  assign new_n6326_ = ~new_n6327_ & (~new_n4725_ | ~new_n4903_ | ~new_n6328_);
  assign new_n6327_ = (\i[1967]  | \i[1966]  | (~\i[1978]  & ~\i[1979] )) & ~new_n6328_ & (new_n4134_ | \i[1978]  | \i[1979] );
  assign new_n6328_ = \i[2751]  & (\i[2750]  | \i[2749] );
  assign new_n6329_ = (~\i[1162]  & ~\i[1163]  & new_n6330_ & ~\i[1161] ) | (~new_n6332_ & (\i[1161]  | \i[1162]  | \i[1163] ));
  assign new_n6330_ = new_n6331_ ? (\i[839]  | (\i[837]  & \i[838] )) : new_n4673_;
  assign new_n6331_ = \i[1967]  & (\i[1966]  | (\i[1965]  & \i[1964] ));
  assign new_n6332_ = \i[1491]  & (\i[1489]  | \i[1490]  | \i[1488] );
  assign new_n6333_ = new_n6348_ ? new_n6334_ : (new_n5802_ ? new_n6345_ : new_n6342_);
  assign new_n6334_ = (new_n6337_ | new_n6339_ | new_n5125_) & (~new_n5125_ | (new_n6341_ ? new_n6335_ : new_n6340_));
  assign new_n6335_ = (new_n4074_ & (~\i[1525]  | ~\i[1526]  | ~\i[1527] )) | (new_n6336_ & \i[1525]  & \i[1526]  & \i[1527] );
  assign new_n6336_ = ~\i[727]  & (~\i[725]  | ~\i[726]  | ~\i[724] );
  assign new_n6337_ = new_n6338_ & (~new_n4215_ | (\i[840]  & \i[841] ));
  assign new_n6338_ = new_n4020_ & (~\i[1647]  | (~\i[1645]  & ~\i[1646] ));
  assign new_n6339_ = ~new_n4020_ & new_n5643_ & \i[1643]  & (\i[1642]  | \i[1641]  | \i[1640] );
  assign new_n6340_ = (\i[850]  & \i[851]  & (~\i[2651]  | (~\i[2649]  & ~\i[2650] ))) | (\i[627]  & (~\i[850]  | ~\i[851] ));
  assign new_n6341_ = ~\i[971]  & ~\i[969]  & ~\i[970] ;
  assign new_n6342_ = new_n4340_ ? new_n6343_ : (new_n4757_ ? new_n6344_ : ~new_n4288_);
  assign new_n6343_ = (\i[2539]  & (\i[2538]  | (\i[2536]  & \i[2537] ))) ? ~new_n4977_ : ~new_n6292_;
  assign new_n6344_ = \i[1171]  & \i[1169]  & \i[1170] ;
  assign new_n6345_ = (new_n6346_ & (~\i[2062]  | ~\i[2063] )) | (\i[2062]  & \i[2063]  & (new_n6347_ ? new_n3396_ : ~new_n4299_));
  assign new_n6346_ = (new_n3450_ & ~\i[735] ) | (~\i[1283]  & \i[735]  & (~\i[1282]  | ~\i[1281] ));
  assign new_n6347_ = \i[2399]  & (\i[2397]  | \i[2398]  | \i[2396] );
  assign new_n6348_ = \i[1855]  & (\i[1853]  | \i[1854]  | \i[1852] );
  assign new_n6349_ = new_n5674_ ? new_n6355_ : ((new_n6364_ | new_n6366_ | ~new_n4091_) & (new_n6350_ | new_n4091_));
  assign new_n6350_ = (new_n6352_ | new_n5155_) & (new_n3242_ | ~new_n6351_);
  assign new_n6351_ = new_n5155_ & new_n6101_ & (~\i[725]  | ~\i[724] );
  assign new_n6352_ = (\i[1098]  & \i[1099] ) ? ~new_n6354_ : ~new_n6353_;
  assign new_n6353_ = \i[1814]  & \i[1815]  & (\i[1813]  | \i[1812] );
  assign new_n6354_ = ~\i[631]  & ~\i[630]  & ~\i[628]  & ~\i[629] ;
  assign new_n6355_ = new_n6363_ ? new_n6359_ : (new_n5857_ ? new_n6358_ : new_n6356_);
  assign new_n6356_ = (~new_n4393_ | ~new_n6357_) & (\i[1995]  | new_n6357_ | (\i[1994]  & (\i[1992]  | \i[1993] )));
  assign new_n6357_ = new_n4289_ & (\i[845]  | \i[844] );
  assign new_n6358_ = (new_n4946_ | (~\i[849]  & new_n3540_)) & (~\i[1953]  | ~\i[1954]  | ~\i[1955]  | \i[849]  | ~new_n3540_);
  assign new_n6359_ = (new_n6360_ | new_n3415_) & (new_n6362_ | ~new_n3415_ | (~new_n5762_ & (\i[938]  | \i[939] )));
  assign new_n6360_ = new_n6147_ ? (\i[1315]  | (\i[1313]  & \i[1314] )) : ~new_n6361_;
  assign new_n6361_ = ~\i[955]  & ~\i[953]  & ~\i[954] ;
  assign new_n6362_ = \i[1859]  & \i[1858]  & \i[1857]  & ~\i[938]  & ~\i[939] ;
  assign new_n6363_ = \i[959]  & (\i[958]  | (\i[957]  & \i[956] ));
  assign new_n6364_ = ~new_n3446_ & (new_n3585_ ? new_n6191_ : new_n6365_);
  assign new_n6365_ = ~\i[2103]  & (~\i[2101]  | ~\i[2102]  | ~\i[2100] );
  assign new_n6366_ = new_n3512_ & new_n3446_ & (\i[2399]  | (\i[2397]  & \i[2398] ));
  assign new_n6367_ = new_n6368_ ? (~new_n6419_ ^ new_n6432_) : (new_n6419_ ^ new_n6432_);
  assign new_n6368_ = new_n6369_ ? (~new_n6394_ ^ new_n6409_) : (new_n6394_ ^ new_n6409_);
  assign new_n6369_ = new_n6370_ ? (new_n6378_ ^ new_n6388_) : (~new_n6378_ ^ new_n6388_);
  assign new_n6370_ = (~new_n6211_ & \i[2860]  & \i[2861]  & \i[2862]  & \i[2863] ) | (new_n6371_ & (~\i[2860]  | ~\i[2861]  | ~\i[2862]  | ~\i[2863] ));
  assign new_n6371_ = ~new_n6374_ & (~new_n4193_ | (~new_n6372_ & (new_n6377_ | ~new_n3219_)));
  assign new_n6372_ = new_n6373_ & (~\i[971]  | (~\i[968]  & ~\i[969]  & ~\i[970] ));
  assign new_n6373_ = ~new_n3219_ & ~\i[2527]  & (~\i[2526]  | ~\i[2525]  | ~\i[2524] );
  assign new_n6374_ = ~new_n4193_ & (new_n6376_ | new_n6375_) & (new_n6132_ | \i[1190]  | \i[1191]  | ~new_n6375_);
  assign new_n6375_ = \i[1391]  & (\i[1389]  | \i[1390]  | \i[1388] );
  assign new_n6376_ = \i[1591]  & \i[1590]  & \i[1588]  & \i[1589] ;
  assign new_n6377_ = ~\i[1539]  & ~\i[1537]  & ~\i[1538] ;
  assign new_n6378_ = (\i[2751]  & (\i[2748]  | \i[2749]  | \i[2750] )) ? new_n6379_ : new_n6383_;
  assign new_n6379_ = ~new_n6380_ & (\i[1735]  | ((new_n6382_ | ~new_n5115_) & (~new_n3731_ | ~new_n4061_ | new_n5115_)));
  assign new_n6380_ = new_n6381_ & (~new_n3714_ | ~\i[1519]  | (~\i[1518]  & (~\i[1516]  | ~\i[1517] )));
  assign new_n6381_ = \i[1735]  & (new_n3714_ | (~\i[2859]  & (\i[2189]  | \i[2190]  | \i[2191] )));
  assign new_n6382_ = \i[1603]  & ~new_n4808_ & \i[1602] ;
  assign new_n6383_ = new_n6387_ ? ((new_n6384_ | ~new_n4674_) & (new_n3761_ | ~new_n5025_ | new_n4674_)) : new_n4710_;
  assign new_n6384_ = (~new_n6385_ | new_n6386_) & (\i[719]  | ~new_n6386_ | (\i[718]  & (\i[716]  | \i[717] )));
  assign new_n6385_ = ~\i[967]  & (~\i[966]  | ~\i[965] );
  assign new_n6386_ = ~\i[2835]  & (~\i[2834]  | (~\i[2833]  & ~\i[2832] ));
  assign new_n6387_ = ~\i[2862]  & ~\i[2863]  & (~\i[2861]  | ~\i[2860] );
  assign new_n6388_ = ~\i[2955]  & ~\i[2954]  & ~\i[2953]  & ~new_n6389_ & ~\i[2952] ;
  assign new_n6389_ = ~new_n6390_ & (new_n4188_ | (~new_n6392_ & new_n5483_) | (~new_n6155_ & new_n6393_ & ~new_n5483_));
  assign new_n6390_ = new_n4188_ & (new_n6391_ | new_n5711_) & (\i[1826]  | \i[1827]  | ~new_n5231_ | ~new_n5711_);
  assign new_n6391_ = ~\i[2271]  & ~\i[2270]  & ~\i[2269]  & ~new_n4391_ & ~\i[2268] ;
  assign new_n6392_ = \i[1423]  & \i[1422]  & ~new_n3569_ & \i[1421] ;
  assign new_n6393_ = ~\i[1879]  & ~\i[1877]  & ~\i[1878] ;
  assign new_n6394_ = new_n3450_ ? new_n6395_ : ((new_n6404_ | new_n6405_ | ~new_n6408_) & (~new_n6402_ | new_n6408_));
  assign new_n6395_ = (new_n6396_ | new_n6397_ | (~\i[1949]  & new_n4657_)) & (new_n6398_ | new_n6401_ | \i[1949]  | ~new_n4657_);
  assign new_n6396_ = ~new_n5196_ & \i[1159]  & new_n5411_ & (\i[1719]  | (\i[1718]  & new_n4817_));
  assign new_n6397_ = new_n5196_ & ((~\i[1747]  & (~\i[1745]  | ~\i[1746] )) ? ~new_n6252_ : ~new_n4277_);
  assign new_n6398_ = (~new_n6399_ | new_n4656_) & (~\i[1826]  | ~\i[1827] ) & (~new_n6400_ | ~new_n4656_);
  assign new_n6399_ = \i[1147]  & \i[1146]  & \i[1144]  & \i[1145] ;
  assign new_n6400_ = ~\i[1207]  & ~\i[1206]  & ~\i[1204]  & ~\i[1205] ;
  assign new_n6401_ = \i[1827]  & \i[1826]  & ~new_n6069_ & new_n6281_;
  assign new_n6402_ = (~\i[1323]  | new_n3538_ | ~new_n3467_) & (new_n3467_ | (new_n5679_ ? new_n6403_ : ~new_n5913_));
  assign new_n6403_ = \i[1831]  & \i[1830]  & \i[1828]  & \i[1829] ;
  assign new_n6404_ = new_n4804_ & new_n3455_ & (~\i[723]  | (~\i[720]  & ~\i[721]  & ~\i[722] ));
  assign new_n6405_ = ~new_n3455_ & (new_n6127_ ? new_n6407_ : ~new_n6406_);
  assign new_n6406_ = ~\i[1051]  & ~\i[1049]  & ~\i[1050] ;
  assign new_n6407_ = \i[735]  & (\i[733]  | \i[734]  | \i[732] );
  assign new_n6408_ = ~\i[1538]  & ~\i[1539]  & (~\i[1537]  | ~\i[1536] );
  assign new_n6409_ = (new_n6410_ | ~new_n6131_) & (~new_n6418_ | new_n6131_ | (\i[967]  & (\i[965]  | \i[966] )));
  assign new_n6410_ = new_n6416_ ? ((~new_n6414_ & ~new_n4326_) | (new_n5913_ & new_n6417_ & new_n4326_)) : new_n6411_;
  assign new_n6411_ = (new_n6412_ | new_n3349_ | ~new_n6087_) & (new_n6087_ | (new_n6413_ ? ~new_n4189_ : ~new_n3628_));
  assign new_n6412_ = ~\i[2311]  & (~\i[2309]  | ~\i[2310]  | ~\i[2308] );
  assign new_n6413_ = ~\i[731]  & (~\i[730]  | (~\i[729]  & ~\i[728] ));
  assign new_n6414_ = new_n6415_ ? (\i[2615]  | (\i[2612]  & \i[2613]  & \i[2614] )) : ~new_n5005_;
  assign new_n6415_ = ~\i[1207]  & (~\i[1205]  | ~\i[1206]  | ~\i[1204] );
  assign new_n6416_ = \i[1954]  & \i[1955] ;
  assign new_n6417_ = ~\i[1983]  & ~\i[1982]  & ~\i[1980]  & ~\i[1981] ;
  assign new_n6418_ = ~\i[2266]  & ~\i[2267]  & (~\i[2265]  | ~\i[2264] );
  assign new_n6419_ = (~\i[1709]  & ~\i[1710]  & ~\i[1711] ) ? (new_n6428_ | new_n6430_) : new_n6420_;
  assign new_n6420_ = new_n4323_ ? new_n6421_ : ((~new_n6426_ | new_n6427_) & (new_n3869_ | ~new_n4062_ | ~new_n6427_));
  assign new_n6421_ = (~new_n4288_ | ~new_n6425_ | new_n6424_) & (new_n6422_ | ~new_n6424_ | (~new_n6423_ & new_n3229_));
  assign new_n6422_ = ~\i[619]  & new_n6423_ & (~\i[618]  | (~\i[616]  & ~\i[617] ));
  assign new_n6423_ = ~\i[1775]  & (~\i[1773]  | ~\i[1774]  | ~\i[1772] );
  assign new_n6424_ = ~\i[951]  & ~\i[949]  & ~\i[950] ;
  assign new_n6425_ = ~\i[1694]  & ~\i[1695]  & (~\i[1693]  | ~\i[1692] );
  assign new_n6426_ = (new_n6400_ | (~\i[966]  & ~\i[967] )) & (\i[629]  | \i[630]  | \i[631]  | \i[966]  | \i[967] );
  assign new_n6427_ = ~\i[1427]  & ~\i[1426]  & ~\i[1424]  & ~\i[1425] ;
  assign new_n6428_ = ~new_n3756_ & (~new_n4949_ | \i[2313] ) & (new_n4285_ ? ~\i[1975]  : ~new_n6429_);
  assign new_n6429_ = ~\i[1502]  & ~\i[1503]  & (~\i[1501]  | ~\i[1500] );
  assign new_n6430_ = ~new_n6104_ & new_n3756_ & (new_n6431_ | ~new_n6101_);
  assign new_n6431_ = ~\i[1495]  & (~\i[1493]  | ~\i[1494]  | ~\i[1492] );
  assign new_n6432_ = new_n6447_ ? (new_n6439_ | (~new_n6444_ & ~new_n6128_ & ~new_n6443_)) : new_n6433_;
  assign new_n6433_ = (new_n5006_ | new_n6436_ | new_n6438_) & (new_n6434_ | ~new_n6437_ | ~new_n6438_);
  assign new_n6434_ = (new_n6435_ & new_n6385_) | (~\i[1663]  & ~new_n6385_ & (~\i[1662]  | ~\i[1661] ));
  assign new_n6435_ = \i[1187]  & (\i[1186]  | (\i[1185]  & \i[1184] ));
  assign new_n6436_ = (new_n3253_ | \i[1719] ) & (\i[2514]  | \i[2515]  | ~\i[1719] );
  assign new_n6437_ = ~\i[515]  & ~\i[514]  & ~\i[512]  & ~\i[513] ;
  assign new_n6438_ = ~\i[747]  & (~\i[746]  | (~\i[745]  & ~\i[744] ));
  assign new_n6439_ = new_n6443_ & (new_n5533_ ? (new_n3540_ ? ~new_n6440_ : new_n6435_) : new_n6441_);
  assign new_n6440_ = new_n4000_ & ~\i[752]  & ~\i[753] ;
  assign new_n6441_ = (~\i[979]  & ~\i[978]  & ~\i[2051]  & (~new_n6442_ | ~\i[2048] )) | (~new_n5062_ & (\i[2051]  | (new_n6442_ & \i[2048] )));
  assign new_n6442_ = \i[2049]  & \i[2050] ;
  assign new_n6443_ = \i[718]  & \i[719]  & (\i[717]  | \i[716] );
  assign new_n6444_ = (~new_n6446_ & ~new_n6445_) | (\i[1597]  & \i[1598]  & \i[1599]  & new_n6445_);
  assign new_n6445_ = ~\i[2219]  & ~\i[2217]  & ~\i[2218] ;
  assign new_n6446_ = ~\i[1754]  & ~\i[1755]  & (~\i[1753]  | ~\i[1752] );
  assign new_n6447_ = ~\i[2502]  & ~\i[2503]  & (~\i[2501]  | ~\i[2500] );
  assign new_n6448_ = new_n6459_ ? new_n6449_ : ((new_n6455_ | ~new_n5435_) & (new_n6460_ | ~new_n4380_ | new_n5435_));
  assign new_n6449_ = (new_n6450_ | ~new_n6454_) & (new_n4659_ | new_n6454_ | (new_n6407_ ? ~new_n3446_ : new_n4494_));
  assign new_n6450_ = new_n6453_ ? (~new_n4362_ | (\i[1818]  & \i[1819] )) : new_n6451_;
  assign new_n6451_ = new_n6452_ & ((\i[733]  & \i[732] ) | \i[735]  | \i[734] );
  assign new_n6452_ = ~\i[2286]  & ~\i[2287]  & (~\i[2285]  | ~\i[2284] );
  assign new_n6453_ = ~\i[1746]  & ~\i[1747]  & (~\i[1745]  | ~\i[1744] );
  assign new_n6454_ = ~\i[834]  & ~\i[835]  & (~\i[833]  | ~\i[832] );
  assign new_n6455_ = (~new_n6458_ | (~\i[743]  & (~\i[741]  | ~\i[742] ))) & (new_n6457_ | new_n6456_ | \i[743]  | (\i[741]  & \i[742] ));
  assign new_n6456_ = new_n5420_ & ~new_n4817_ & new_n3395_;
  assign new_n6457_ = ~new_n5420_ & (\i[2613]  | \i[2614]  | \i[2615] );
  assign new_n6458_ = \i[1703]  & \i[1702]  & \i[1701]  & ~new_n4823_ & \i[1700] ;
  assign new_n6459_ = new_n3264_ & ~\i[2388]  & ~\i[2389] ;
  assign new_n6460_ = new_n6461_ & (~\i[2771]  | (~\i[2768]  & ~\i[2769]  & ~\i[2770] ));
  assign new_n6461_ = ~\i[1783]  & ~\i[1782]  & ~\i[1780]  & ~\i[1781] ;
  assign new_n6462_ = new_n4142_ ? new_n6463_ : ((new_n6467_ | ~new_n4080_) & (new_n6471_ | new_n6474_ | new_n4080_));
  assign new_n6463_ = new_n3775_ ? (~new_n6466_ & (new_n4002_ | new_n4299_ | ~\i[1639] )) : new_n6464_;
  assign new_n6464_ = (~new_n3594_ | ~new_n4285_ | ~new_n6465_) & (~new_n6266_ | new_n6465_ | (~\i[1281]  & new_n5052_));
  assign new_n6465_ = ~\i[771]  & (~\i[769]  | ~\i[770]  | ~\i[768] );
  assign new_n6466_ = ~\i[1639]  & \i[1095]  & new_n4362_ & (\i[1094]  | \i[1093]  | \i[1092] );
  assign new_n6467_ = (new_n6468_ | ~new_n5200_) & (~new_n6470_ | ~new_n4050_ | new_n5200_);
  assign new_n6468_ = new_n6469_ ? (~\i[1503]  | (~\i[1501]  & ~\i[1502] )) : new_n5563_;
  assign new_n6469_ = ~\i[1483]  & ~\i[1482]  & ~\i[1480]  & ~\i[1481] ;
  assign new_n6470_ = new_n4109_ & (~\i[1841]  | ~\i[1840] );
  assign new_n6471_ = new_n5062_ & ((~new_n6472_ & new_n6473_) | (\i[1597]  & \i[1598]  & \i[1599]  & ~new_n6473_));
  assign new_n6472_ = ~\i[1826]  & ~\i[1827]  & (~\i[1825]  | ~\i[1824] );
  assign new_n6473_ = ~\i[2279]  & (~\i[2278]  | (~\i[2277]  & ~\i[2276] ));
  assign new_n6474_ = ~new_n5062_ & (new_n6475_ ? new_n5108_ : ~new_n3239_);
  assign new_n6475_ = \i[1711]  & \i[1709]  & \i[1710] ;
  assign \o[29]  = new_n6477_ ^ new_n6478_;
  assign new_n6477_ = ~new_n6052_ & ~new_n6462_;
  assign new_n6478_ = new_n6479_ ? (~new_n6480_ ^ new_n6573_) : (new_n6480_ ^ new_n6573_);
  assign new_n6479_ = (~new_n6367_ & ~new_n6448_) | (~new_n6053_ & (~new_n6367_ | ~new_n6448_));
  assign new_n6480_ = new_n6481_ ? (~new_n6482_ ^ new_n6560_) : (new_n6482_ ^ new_n6560_);
  assign new_n6481_ = (~new_n6183_ & ~new_n6349_) | (~new_n6054_ & (~new_n6183_ | ~new_n6349_));
  assign new_n6482_ = new_n6483_ ? (~new_n6506_ ^ new_n6507_) : (new_n6506_ ^ new_n6507_);
  assign new_n6483_ = new_n6484_ ? (new_n6485_ ^ new_n6505_) : (~new_n6485_ ^ new_n6505_);
  assign new_n6484_ = (~new_n6105_ & new_n6148_) | (~new_n6056_ & (~new_n6105_ | new_n6148_));
  assign new_n6485_ = new_n6486_ ? (new_n6487_ ^ new_n6497_) : (~new_n6487_ ^ new_n6497_);
  assign new_n6486_ = (~new_n6088_ & new_n6075_) | (~new_n6057_ & (~new_n6088_ | new_n6075_));
  assign new_n6487_ = new_n6488_ ? (new_n6492_ ^ new_n6495_) : (~new_n6492_ ^ new_n6495_);
  assign new_n6488_ = new_n5674_ ? ((~new_n6491_ | new_n6363_) & (~new_n3415_ | ~new_n6362_ | ~new_n6363_)) : new_n6489_;
  assign new_n6489_ = (~new_n3446_ | ~new_n6490_ | ~new_n4091_) & (~new_n6351_ | ~new_n3242_ | new_n4091_);
  assign new_n6490_ = ~\i[2399]  & \i[1987]  & \i[1986]  & (~\i[2398]  | ~\i[2397] );
  assign new_n6491_ = new_n5857_ & new_n4946_ & (\i[851]  | \i[850]  | \i[849] );
  assign new_n6492_ = new_n4682_ & (new_n6494_ | (new_n6493_ & new_n6196_));
  assign new_n6493_ = ~new_n4285_ & ~new_n6194_ & ((~\i[968]  & ~\i[969] ) | ~\i[971]  | ~\i[970] );
  assign new_n6494_ = new_n3672_ & new_n4285_ & ~new_n5005_ & ~new_n6198_;
  assign new_n6495_ = new_n6447_ & (new_n6496_ | (~new_n6128_ & ~new_n6443_ & ~new_n6445_ & new_n6446_));
  assign new_n6496_ = new_n5533_ & new_n6443_ & (new_n3540_ ? ~new_n6440_ : new_n6435_);
  assign new_n6497_ = new_n6498_ ? (new_n6502_ ^ new_n6504_) : (~new_n6502_ ^ new_n6504_);
  assign new_n6498_ = (~new_n4946_ | new_n6499_ | new_n5675_) & (~new_n5675_ | (~new_n6500_ & (new_n6501_ | new_n6203_)));
  assign new_n6499_ = (~new_n6282_ | new_n3377_) & (~new_n4310_ | ~new_n3377_ | (\i[519]  & (\i[517]  | \i[518] )));
  assign new_n6500_ = new_n6285_ & new_n6287_ & new_n4342_ & new_n6203_ & (\i[841]  | \i[840] );
  assign new_n6501_ = (~new_n5742_ | ~new_n4246_ | ~new_n4471_) & (~new_n4379_ | new_n4471_ | (\i[1179]  & \i[1178] ));
  assign new_n6502_ = ~new_n6171_ & (new_n6164_ ? (new_n6162_ | (new_n6159_ & new_n3750_)) : ~new_n6503_);
  assign new_n6503_ = (\i[954]  | \i[955]  | ~new_n6413_ | ~new_n5665_) & (~new_n4342_ | new_n4029_ | new_n5665_);
  assign new_n6504_ = new_n6318_ & new_n6317_ & ~new_n6131_ & new_n6132_;
  assign new_n6505_ = (~new_n6321_ & new_n6268_) | (~new_n6270_ & (~new_n6321_ | new_n6268_));
  assign new_n6506_ = (~new_n6269_ & ~new_n6333_) | (~new_n6184_ & (~new_n6269_ | ~new_n6333_));
  assign new_n6507_ = new_n6508_ ? (~new_n6509_ ^ new_n6526_) : (new_n6509_ ^ new_n6526_);
  assign new_n6508_ = (~new_n6226_ & new_n6268_) | (~new_n6185_ & (~new_n6226_ | new_n6268_));
  assign new_n6509_ = new_n6510_ ? (new_n6511_ ^ new_n6512_) : (~new_n6511_ ^ new_n6512_);
  assign new_n6510_ = (~new_n6216_ & new_n6199_) | (new_n6186_ & (~new_n6216_ | new_n6199_));
  assign new_n6511_ = (~new_n6293_ & ~new_n6309_) | (~new_n6271_ & (~new_n6293_ | ~new_n6309_));
  assign new_n6512_ = new_n6513_ ? (new_n6521_ ^ new_n6524_) : (~new_n6521_ ^ new_n6524_);
  assign new_n6513_ = (~\i[1709]  & ~\i[1710]  & ~\i[1711] ) ? (new_n6518_ | ~new_n3756_) : new_n6514_;
  assign new_n6514_ = new_n4323_ ? new_n6515_ : (new_n6427_ ? new_n6516_ : ~new_n6517_);
  assign new_n6515_ = new_n6424_ ? ~new_n6422_ : new_n6425_;
  assign new_n6516_ = new_n4062_ ? ~new_n3869_ : (\i[2971]  & (\i[2968]  | \i[2969]  | \i[2970] ));
  assign new_n6517_ = ~\i[967]  & ~\i[966]  & ~\i[631]  & ~\i[629]  & ~\i[630] ;
  assign new_n6518_ = (~new_n6431_ | ~new_n6520_ | new_n6104_) & (new_n6198_ | new_n6519_ | ~new_n6104_);
  assign new_n6519_ = ~\i[1947]  & ~\i[1946]  & ~\i[1944]  & ~\i[1945] ;
  assign new_n6520_ = \i[2843]  & \i[2841]  & \i[2842] ;
  assign new_n6521_ = ~new_n6522_ & (~new_n6523_ | ~new_n3683_ | ~new_n4684_);
  assign new_n6522_ = new_n4056_ & new_n6069_ & new_n5449_ & ~new_n3800_ & ~new_n6212_;
  assign new_n6523_ = new_n6212_ & new_n6204_ & ~\i[2271]  & ~\i[2270]  & ~\i[2268]  & ~\i[2269] ;
  assign new_n6524_ = ~new_n6225_ & ((~new_n6222_ & ~new_n6221_) | (~new_n6219_ & ~new_n6525_ & new_n3309_ & new_n6221_));
  assign new_n6525_ = \i[1042]  & \i[1043] ;
  assign new_n6526_ = new_n6527_ ? (~new_n6528_ ^ new_n6550_) : (new_n6528_ ^ new_n6550_);
  assign new_n6527_ = (~new_n6244_ & ~new_n6255_) | (~new_n6227_ & (~new_n6244_ | ~new_n6255_));
  assign new_n6528_ = new_n6529_ ? (new_n6536_ ^ new_n6546_) : (~new_n6536_ ^ new_n6546_);
  assign new_n6529_ = new_n6459_ ? new_n6532_ : new_n6530_;
  assign new_n6530_ = (new_n6531_ | ~new_n5435_) & (new_n4380_ | \i[2158]  | \i[2159]  | ~new_n5483_ | new_n5435_);
  assign new_n6531_ = (~new_n4216_ | ~new_n4823_ | (~\i[743]  & (~\i[741]  | ~\i[742] ))) & (~new_n6457_ | \i[743]  | (\i[741]  & \i[742] ));
  assign new_n6532_ = (new_n6533_ | ~new_n6454_) & (new_n6534_ | ~new_n4946_ | ~new_n4659_ | new_n6454_);
  assign new_n6533_ = (~new_n6451_ | new_n6453_) & (~new_n4362_ | ~\i[1818]  | ~\i[1819]  | ~new_n6453_);
  assign new_n6534_ = new_n6535_ & ~\i[872]  & ~\i[873] ;
  assign new_n6535_ = ~\i[874]  & ~\i[875] ;
  assign new_n6536_ = new_n6254_ ? (new_n5636_ ? new_n6542_ : new_n6544_) : new_n6537_;
  assign new_n6537_ = new_n6253_ ? new_n6538_ : ((~new_n6541_ | ~new_n5025_) & (new_n6247_ | ~new_n3613_ | new_n5025_));
  assign new_n6538_ = (~new_n6540_ | ~new_n6539_) & (~new_n5668_ | ~new_n4285_ | new_n6539_);
  assign new_n6539_ = \i[1593]  & new_n3348_ & \i[1592] ;
  assign new_n6540_ = \i[1159]  & ((~\i[2209]  & ~\i[2208] ) | ~\i[2211]  | ~\i[2210] );
  assign new_n6541_ = ~new_n4143_ & (~\i[2291]  | (~\i[2288]  & ~\i[2289]  & ~\i[2290] ));
  assign new_n6542_ = (~new_n6250_ | ~\i[1635]  | (~\i[1633]  & ~\i[1634] )) & (~new_n6251_ | ~new_n6543_ | (\i[1635]  & (\i[1633]  | \i[1634] )));
  assign new_n6543_ = \i[1959]  & (\i[1958]  | \i[1957] );
  assign new_n6544_ = (~new_n6545_ | ~new_n6127_) & (\i[746]  | \i[747]  | ~new_n3628_ | new_n6127_);
  assign new_n6545_ = ~\i[731]  & ~\i[375]  & ~\i[374]  & ~\i[372]  & ~\i[373] ;
  assign new_n6546_ = (new_n6548_ | new_n6547_ | ~new_n4142_) & (new_n4142_ | (new_n4080_ ? new_n6549_ : ~new_n6471_));
  assign new_n6547_ = ~new_n3775_ & (new_n6465_ | \i[1281]  | \i[1282]  | \i[1283]  | ~new_n6266_);
  assign new_n6548_ = new_n3775_ & (~new_n4002_ | ~new_n6101_ | ~\i[1639]  | (\i[725]  & \i[724] ));
  assign new_n6549_ = (new_n6469_ | ~new_n5563_ | ~new_n5200_) & (new_n5200_ | (new_n4050_ ? new_n6470_ : new_n6135_));
  assign new_n6550_ = new_n6551_ ^ new_n6557_;
  assign new_n6551_ = ~new_n6552_ & (~new_n6267_ | (~new_n6554_ & (~new_n6238_ | new_n6556_)));
  assign new_n6552_ = ~new_n6267_ & (new_n6553_ | (~new_n3413_ & new_n5079_ & \i[1391] ));
  assign new_n6553_ = ~new_n5079_ & new_n5035_ & new_n6266_ & (\i[771]  | \i[770]  | \i[769] );
  assign new_n6554_ = new_n5843_ & new_n6555_ & new_n5230_ & (~\i[2165]  | ~\i[2164] );
  assign new_n6555_ = ~new_n6238_ & ((\i[253]  & \i[252] ) | \i[255]  | \i[254] );
  assign new_n6556_ = (new_n3800_ | ~new_n5730_ | ~new_n6261_) & (~new_n3525_ | ~new_n4246_ | new_n6261_);
  assign new_n6557_ = (new_n6558_ | new_n6155_) & (new_n5066_ | ~new_n6155_ | (new_n3399_ ? ~new_n6559_ : ~new_n6236_));
  assign new_n6558_ = (new_n4019_ | new_n5743_ | ~new_n4069_ | ~new_n6240_) & (~new_n4019_ | ~new_n5743_ | new_n4080_ | ~new_n3775_);
  assign new_n6559_ = new_n4785_ & new_n5675_;
  assign new_n6560_ = new_n6561_ ? (new_n6562_ ^ new_n6572_) : (~new_n6562_ ^ new_n6572_);
  assign new_n6561_ = (~new_n6156_ & new_n6173_) | (~new_n6055_ & (~new_n6156_ | new_n6173_));
  assign new_n6562_ = new_n6563_ ? (~new_n6564_ ^ new_n6565_) : (new_n6564_ ^ new_n6565_);
  assign new_n6563_ = (~new_n6123_ & ~new_n6133_) | (~new_n6106_ & (~new_n6123_ | ~new_n6133_));
  assign new_n6564_ = (~new_n6378_ & new_n6388_) | (~new_n6370_ & (~new_n6378_ | new_n6388_));
  assign new_n6565_ = (new_n4190_ & new_n6571_ & new_n6308_ & new_n6297_ & (new_n6566_ ^ ~new_n6567_)) | ((~new_n4190_ | ~new_n6571_ | ~new_n6308_ | ~new_n6297_) & (new_n6566_ ^ new_n6567_));
  assign new_n6566_ = ~new_n4070_ & (new_n4266_ ? new_n6079_ : new_n6083_);
  assign new_n6567_ = (~new_n6568_ & ~new_n6569_ & ~new_n6348_) | (new_n6348_ & (~new_n6336_ | ~new_n6570_));
  assign new_n6568_ = \i[2063]  & \i[2062]  & new_n5802_ & ~new_n4299_ & ~new_n6347_;
  assign new_n6569_ = new_n6344_ & new_n4757_ & ~new_n4340_ & ~new_n5802_;
  assign new_n6570_ = \i[1527]  & \i[1526]  & \i[1525]  & new_n5125_ & new_n6341_;
  assign new_n6571_ = new_n3229_ & new_n6296_;
  assign new_n6572_ = (~new_n6394_ & ~new_n6409_) | (~new_n6369_ & (~new_n6394_ | ~new_n6409_));
  assign new_n6573_ = (~new_n6419_ & ~new_n6432_) | (~new_n6368_ & (~new_n6419_ | ~new_n6432_));
  assign \o[30]  = ~new_n6575_ ^ new_n6576_;
  assign new_n6575_ = new_n6477_ & new_n6478_;
  assign new_n6576_ = new_n6577_ ^ new_n6578_;
  assign new_n6577_ = (new_n6480_ & new_n6573_) | (new_n6479_ & (new_n6480_ | new_n6573_));
  assign new_n6578_ = new_n6579_ ? (~new_n6580_ ^ new_n6608_) : (new_n6580_ ^ new_n6608_);
  assign new_n6579_ = (new_n6482_ & new_n6560_) | (new_n6481_ & (new_n6482_ | new_n6560_));
  assign new_n6580_ = new_n6581_ ? (new_n6587_ ^ new_n6588_) : (~new_n6587_ ^ new_n6588_);
  assign new_n6581_ = new_n6582_ ? (~new_n6583_ ^ new_n6584_) : (new_n6583_ ^ new_n6584_);
  assign new_n6582_ = (~new_n6485_ & new_n6505_) | (new_n6484_ & (~new_n6485_ | new_n6505_));
  assign new_n6583_ = (~new_n6565_ & new_n6564_) | (new_n6563_ & (~new_n6565_ | new_n6564_));
  assign new_n6584_ = new_n6585_ ^ new_n6586_;
  assign new_n6585_ = (~new_n6566_ | (new_n6567_ & (~new_n6308_ | ~new_n6297_ | ~new_n4190_ | ~new_n6571_))) & (new_n6567_ | ~new_n4190_ | ~new_n6571_ | ~new_n6308_ | ~new_n6297_);
  assign new_n6586_ = (new_n6502_ & new_n6504_) | (~new_n6498_ & (new_n6502_ | new_n6504_));
  assign new_n6587_ = (new_n6506_ & new_n6507_) | (new_n6483_ & (new_n6506_ | new_n6507_));
  assign new_n6588_ = new_n6589_ ? (new_n6593_ ^ new_n6594_) : (~new_n6593_ ^ new_n6594_);
  assign new_n6589_ = new_n6590_ ? (new_n6591_ ^ new_n6592_) : (~new_n6591_ ^ new_n6592_);
  assign new_n6590_ = (new_n6487_ & new_n6497_) | (new_n6486_ & (new_n6487_ | new_n6497_));
  assign new_n6591_ = (~new_n6512_ & new_n6511_) | (new_n6510_ & (~new_n6512_ | new_n6511_));
  assign new_n6592_ = (new_n6492_ & new_n6495_) | (~new_n6488_ & (new_n6492_ | new_n6495_));
  assign new_n6593_ = (new_n6509_ & new_n6526_) | (new_n6508_ & (new_n6509_ | new_n6526_));
  assign new_n6594_ = new_n6595_ ? (new_n6598_ ^ new_n6599_) : (~new_n6598_ ^ new_n6599_);
  assign new_n6595_ = ~new_n6596_ ^ new_n6597_;
  assign new_n6596_ = (~new_n6536_ & ~new_n6546_) | (~new_n6529_ & (~new_n6536_ | ~new_n6546_));
  assign new_n6597_ = (~new_n6521_ & new_n6524_) | (~new_n6513_ & (~new_n6521_ | new_n6524_));
  assign new_n6598_ = (new_n6528_ & new_n6550_) | (new_n6527_ & (new_n6528_ | new_n6550_));
  assign new_n6599_ = new_n6600_ ^ new_n6607_;
  assign new_n6600_ = ~new_n6601_ ^ new_n6606_;
  assign new_n6601_ = (new_n6602_ | ~new_n6155_) & (~new_n6243_ | ~new_n4019_ | new_n6155_ | new_n5743_ | new_n6605_);
  assign new_n6602_ = new_n5066_ ? new_n6603_ : (new_n3399_ ? ~new_n6604_ : ~new_n6236_);
  assign new_n6603_ = (~new_n5022_ | ~new_n6231_ | new_n4837_) & (new_n6235_ | ~new_n6233_ | ~new_n4837_);
  assign new_n6604_ = new_n4785_ ? new_n5675_ : new_n5802_;
  assign new_n6605_ = ~\i[1187]  & (~\i[1186]  | ~\i[1185] );
  assign new_n6606_ = ~new_n6552_ & (new_n6556_ | ~new_n6238_ | ~new_n6267_);
  assign new_n6607_ = ~new_n6551_ & new_n6557_;
  assign new_n6608_ = (~new_n6562_ & new_n6572_) | (new_n6561_ & (~new_n6562_ | new_n6572_));
  assign \o[31]  = ((new_n6610_ | new_n6611_) & (~new_n6612_ ^ new_n6613_)) | (~new_n6610_ & ~new_n6611_ & (~new_n6612_ ^ ~new_n6613_));
  assign new_n6610_ = ~new_n6576_ & new_n6575_;
  assign new_n6611_ = ~new_n6578_ & new_n6577_;
  assign new_n6612_ = (~new_n6580_ & new_n6608_) | (new_n6579_ & (~new_n6580_ | new_n6608_));
  assign new_n6613_ = new_n6614_ ? (new_n6615_ ^ new_n6626_) : (~new_n6615_ ^ new_n6626_);
  assign new_n6614_ = (~new_n6588_ & new_n6587_) | (~new_n6581_ & (~new_n6588_ | new_n6587_));
  assign new_n6615_ = new_n6616_ ? (new_n6619_ ^ new_n6620_) : (~new_n6619_ ^ new_n6620_);
  assign new_n6616_ = ~new_n6617_ ^ new_n6618_;
  assign new_n6617_ = (new_n6591_ & new_n6592_) | (new_n6590_ & (new_n6591_ | new_n6592_));
  assign new_n6618_ = ~new_n6585_ & new_n6586_;
  assign new_n6619_ = (~new_n6594_ & new_n6593_) | (~new_n6589_ & (~new_n6594_ | new_n6593_));
  assign new_n6620_ = new_n6621_ ? (~new_n6622_ ^ new_n6625_) : (new_n6622_ ^ new_n6625_);
  assign new_n6621_ = (~new_n6599_ & new_n6598_) | (~new_n6595_ & (~new_n6599_ | new_n6598_));
  assign new_n6622_ = new_n6623_ ^ new_n6624_;
  assign new_n6623_ = ~new_n6607_ & new_n6600_;
  assign new_n6624_ = new_n6601_ & new_n6606_;
  assign new_n6625_ = new_n6596_ & new_n6597_;
  assign new_n6626_ = (~new_n6584_ & new_n6583_) | (new_n6582_ & (~new_n6584_ | new_n6583_));
  assign \o[32]  = ~new_n6628_ ^ new_n6629_;
  assign new_n6628_ = (new_n6613_ | new_n6610_ | new_n6611_) & (new_n6612_ | (new_n6613_ & (new_n6610_ | new_n6611_)));
  assign new_n6629_ = new_n6630_ ^ new_n6631_;
  assign new_n6630_ = (~new_n6615_ & new_n6626_) | (new_n6614_ & (~new_n6615_ | new_n6626_));
  assign new_n6631_ = new_n6632_ ? (~new_n6633_ ^ new_n6634_) : (new_n6633_ ^ new_n6634_);
  assign new_n6632_ = (~new_n6620_ & new_n6619_) | (~new_n6616_ & (~new_n6620_ | new_n6619_));
  assign new_n6633_ = new_n6617_ & new_n6618_;
  assign new_n6634_ = ~new_n6635_ ^ new_n6636_;
  assign new_n6635_ = (~new_n6622_ & new_n6625_) | (new_n6621_ & (~new_n6622_ | new_n6625_));
  assign new_n6636_ = ~new_n6624_ & new_n6623_;
  assign \o[33]  = ((new_n6638_ | new_n6639_) & (~new_n6640_ ^ new_n6641_)) | (~new_n6638_ & ~new_n6639_ & (~new_n6640_ ^ ~new_n6641_));
  assign new_n6638_ = ~new_n6629_ & new_n6628_;
  assign new_n6639_ = ~new_n6631_ & new_n6630_;
  assign new_n6640_ = (~new_n6634_ & new_n6633_) | (new_n6632_ & (~new_n6634_ | new_n6633_));
  assign new_n6641_ = new_n6635_ & new_n6636_;
  assign \o[34]  = (new_n6641_ | new_n6638_ | new_n6639_) & (new_n6640_ | (new_n6641_ & (new_n6638_ | new_n6639_)));
  assign \o[35]  = new_n6644_ ^ new_n7024_;
  assign new_n6644_ = new_n6645_ ? (new_n6998_ ^ new_n7009_) : (~new_n6998_ ^ new_n7009_);
  assign new_n6645_ = new_n6646_ ? (new_n6933_ ^ new_n6989_) : (~new_n6933_ ^ new_n6989_);
  assign new_n6646_ = new_n6647_ ? (new_n6800_ ^ new_n6913_) : (~new_n6800_ ^ new_n6913_);
  assign new_n6647_ = new_n6648_ ? (new_n6735_ ^ new_n6787_) : (~new_n6735_ ^ new_n6787_);
  assign new_n6648_ = new_n6649_ ? (new_n6694_ ^ new_n6733_) : (~new_n6694_ ^ new_n6733_);
  assign new_n6649_ = new_n6650_ ? (~new_n6666_ ^ new_n6685_) : (new_n6666_ ^ new_n6685_);
  assign new_n6650_ = ~new_n6651_ & (new_n3624_ | (~new_n6660_ & ~new_n3376_) | (new_n6664_ & new_n6665_ & new_n3376_));
  assign new_n6651_ = new_n3624_ & (new_n6652_ | ~\i[1942]  | ~\i[1943] ) & (new_n6659_ | new_n6657_ | (\i[1942]  & \i[1943] ));
  assign new_n6652_ = new_n4520_ ? (new_n6654_ | (~new_n6656_ & new_n6655_)) : new_n6653_;
  assign new_n6653_ = new_n5717_ ? new_n4837_ : new_n5195_;
  assign new_n6654_ = ~\i[427]  & ~\i[426]  & ~\i[425]  & ~new_n6655_ & ~\i[424] ;
  assign new_n6655_ = ~\i[415]  & ~\i[414]  & ~\i[412]  & ~\i[413] ;
  assign new_n6656_ = ~\i[1715]  & (~\i[1714]  | (~\i[1713]  & ~\i[1712] ));
  assign new_n6657_ = new_n3223_ & ((~new_n4067_ & ~new_n6658_) | (~\i[983]  & new_n6658_ & (~\i[982]  | ~\i[981] )));
  assign new_n6658_ = ~\i[751]  & ~\i[750]  & ~\i[748]  & ~\i[749] ;
  assign new_n6659_ = ~new_n3505_ & ~new_n3470_ & ~new_n3223_;
  assign new_n6660_ = (~new_n6661_ | ~new_n4352_) & (new_n6663_ | ~new_n6662_ | new_n4352_);
  assign new_n6661_ = \i[771]  & \i[770]  & \i[769]  & ~new_n3385_ & \i[768] ;
  assign new_n6662_ = \i[1501]  & new_n4273_ & \i[1500] ;
  assign new_n6663_ = \i[2435]  & \i[2434]  & \i[2432]  & \i[2433] ;
  assign new_n6664_ = \i[1419]  & \i[1418]  & \i[1417]  & ~new_n3323_ & \i[1416] ;
  assign new_n6665_ = ~\i[2287]  & (~\i[2286]  | (~\i[2285]  & ~\i[2284] ));
  assign new_n6666_ = (new_n6674_ | new_n6667_ | ~new_n4380_) & (new_n4380_ | (new_n6684_ ? new_n6681_ : new_n6678_));
  assign new_n6667_ = ~new_n6669_ & (new_n6673_ ? ~new_n6668_ : (new_n6670_ ? new_n6672_ : ~new_n6671_));
  assign new_n6668_ = new_n3467_ ? new_n3889_ : ~new_n4206_;
  assign new_n6669_ = ~\i[655]  & ~\i[654]  & ~\i[652]  & ~\i[653] ;
  assign new_n6670_ = ~\i[1311]  & ~\i[1310]  & ~\i[1308]  & ~\i[1309] ;
  assign new_n6671_ = \i[2034]  & \i[2035]  & (\i[2033]  | \i[2032] );
  assign new_n6672_ = \i[2527]  & (\i[2526]  | \i[2525] );
  assign new_n6673_ = ~\i[1091]  & ~\i[1090]  & ~\i[1088]  & ~\i[1089] ;
  assign new_n6674_ = new_n6669_ & (new_n6677_ ? (~new_n4018_ | ~new_n3437_) : new_n6675_);
  assign new_n6675_ = new_n4433_ ? ~new_n6676_ : ~new_n3618_;
  assign new_n6676_ = new_n3409_ & ~\i[1544]  & ~\i[1545] ;
  assign new_n6677_ = ~\i[1111]  & ~\i[1110]  & ~\i[1108]  & ~\i[1109] ;
  assign new_n6678_ = (new_n3494_ | ~new_n6679_ | ~new_n6680_) & (new_n4392_ | ~new_n6400_ | new_n6680_);
  assign new_n6679_ = new_n4391_ & (\i[1185]  | \i[1184] );
  assign new_n6680_ = ~\i[1423]  & ~\i[1422]  & ~\i[1420]  & ~\i[1421] ;
  assign new_n6681_ = new_n3318_ ? new_n6682_ : ~new_n6683_;
  assign new_n6682_ = \i[1302]  & \i[1303]  & (\i[1301]  | \i[1300] );
  assign new_n6683_ = ~\i[1323]  & ~\i[1321]  & ~\i[1322] ;
  assign new_n6684_ = ~\i[1315]  & ~\i[1314]  & ~\i[1312]  & ~\i[1313] ;
  assign new_n6685_ = (new_n6686_ | ~new_n5698_) & (new_n6692_ | new_n6693_ | new_n3998_ | new_n5698_);
  assign new_n6686_ = new_n6691_ ? ((~new_n6689_ | ~new_n5126_) & (~new_n3555_ | ~new_n6690_ | new_n5126_)) : new_n6687_;
  assign new_n6687_ = (~new_n3342_ | ~new_n3400_ | ~new_n3376_) & (new_n4190_ | ~new_n6688_ | new_n3376_);
  assign new_n6688_ = \i[411]  & \i[410]  & \i[408]  & \i[409] ;
  assign new_n6689_ = new_n5031_ & (\i[765]  | ~new_n4031_);
  assign new_n6690_ = ~\i[1427]  & ~\i[1425]  & ~\i[1426] ;
  assign new_n6691_ = ~\i[1307]  & ~\i[1306]  & ~\i[1304]  & ~\i[1305] ;
  assign new_n6692_ = new_n4445_ & (new_n4810_ ? ~\i[1411]  : new_n4939_);
  assign new_n6693_ = ~new_n4445_ & (\i[1083]  | ~new_n5856_ | (\i[1082]  & (\i[1080]  | \i[1081] )));
  assign new_n6694_ = new_n6695_ ? (new_n6710_ ^ new_n6721_) : (~new_n6710_ ^ new_n6721_);
  assign new_n6695_ = (new_n6700_ | new_n6696_ | ~new_n3905_) & (new_n3905_ | (new_n6708_ ? new_n6704_ : new_n6706_));
  assign new_n6696_ = ~new_n4100_ & ((~new_n6697_ & new_n6699_) | (~new_n4090_ & ~\i[1839]  & ~new_n6699_));
  assign new_n6697_ = ~new_n6698_ & (\i[1038]  | \i[1039]  | ~new_n6067_ | (\i[1037]  & \i[1036] ));
  assign new_n6698_ = ~\i[1375]  & ~\i[1374]  & ~new_n6067_ & ~\i[1373] ;
  assign new_n6699_ = \i[1827]  & (\i[1826]  | (\i[1825]  & \i[1824] ));
  assign new_n6700_ = new_n6701_ & (new_n6703_ | \i[2206]  | \i[2207] );
  assign new_n6701_ = new_n4100_ & (~new_n6702_ | (~new_n5762_ & ~\i[745]  & ~\i[746]  & ~\i[747] ));
  assign new_n6702_ = (\i[2207]  | \i[2206] ) & (~new_n5762_ | (\i[1047]  & (\i[1045]  | \i[1046] )));
  assign new_n6703_ = (~new_n3273_ & ~new_n3448_) | (\i[503]  & new_n3448_ & (\i[502]  | \i[501] ));
  assign new_n6704_ = new_n6440_ ? new_n6705_ : (new_n4067_ ? new_n6424_ : ~new_n4099_);
  assign new_n6705_ = new_n5568_ ? ~\i[1331]  : ~new_n3892_;
  assign new_n6706_ = ~new_n6707_ & (new_n4810_ | ~\i[2834]  | ~\i[2835]  | (~\i[2833]  & ~\i[2832] ));
  assign new_n6707_ = new_n4810_ & (~new_n4275_ | ~new_n4175_) & (~\i[1529]  | ~\i[1530]  | ~\i[1531]  | new_n4175_);
  assign new_n6708_ = new_n6709_ & ~\i[1100]  & ~\i[1101] ;
  assign new_n6709_ = ~\i[1102]  & ~\i[1103] ;
  assign new_n6710_ = new_n3376_ ? ((~new_n6717_ & ~new_n6720_ & new_n5651_) | (~new_n6715_ & ~new_n5651_)) : new_n6711_;
  assign new_n6711_ = (~new_n6712_ | ~new_n6713_) & (new_n5460_ | new_n6714_ | new_n6713_);
  assign new_n6712_ = ~new_n3892_ & ~\i[1223]  & (~\i[1191]  | ~\i[1190]  | ~\i[1189] );
  assign new_n6713_ = ~\i[1303]  & (~\i[1302]  | (~\i[1301]  & ~\i[1300] ));
  assign new_n6714_ = \i[1103]  & (\i[1102]  | (\i[1101]  & \i[1100] ));
  assign new_n6715_ = (~new_n3219_ | new_n5025_ | new_n3364_) & (~new_n3364_ | (new_n6682_ ? new_n6716_ : new_n4220_));
  assign new_n6716_ = \i[2271]  & \i[2270]  & \i[2268]  & \i[2269] ;
  assign new_n6717_ = new_n6718_ & (new_n5176_ ? ~new_n6719_ : (~\i[1719]  | (~\i[1717]  & ~\i[1718] )));
  assign new_n6718_ = \i[1819]  & (\i[1817]  | \i[1818]  | \i[1816] );
  assign new_n6719_ = ~\i[1367]  & ~\i[1366]  & ~\i[1364]  & ~\i[1365] ;
  assign new_n6720_ = ~new_n6535_ & ~new_n6718_ & ~\i[626]  & ~\i[627]  & (~\i[625]  | ~\i[624] );
  assign new_n6721_ = (~new_n6732_ & ~new_n6725_ & new_n3854_) | (~new_n3854_ & (new_n6722_ | (~new_n6730_ & new_n6724_)));
  assign new_n6722_ = \i[651]  & new_n6723_ & ~new_n3771_ & ~new_n6688_;
  assign new_n6723_ = ~new_n6724_ & (\i[650]  | (\i[648]  & \i[649] ));
  assign new_n6724_ = ~\i[1415]  & ~\i[1413]  & ~\i[1414] ;
  assign new_n6725_ = ~new_n3789_ & (new_n6728_ ? (new_n6726_ ? \i[1291]  : new_n6729_) : ~new_n6727_);
  assign new_n6726_ = new_n3556_ & (~\i[1297]  | ~\i[1296] );
  assign new_n6727_ = ~new_n4785_ & \i[1107]  & (\i[1106]  | \i[1105]  | \i[1104] );
  assign new_n6728_ = \i[2639]  & (\i[2637]  | \i[2638]  | \i[2636] );
  assign new_n6729_ = \i[1739]  & (\i[1738]  | \i[1737] );
  assign new_n6730_ = (new_n5826_ | ~new_n4880_ | new_n3259_) & (~new_n3259_ | (new_n3229_ ? ~new_n4881_ : ~new_n6731_));
  assign new_n6731_ = \i[1295]  & (\i[1294]  | \i[1293] );
  assign new_n6732_ = new_n3789_ & ((~new_n5828_ & ~new_n6655_ & new_n5197_) | (~new_n3587_ & new_n3695_ & ~new_n5197_));
  assign new_n6733_ = new_n6734_ & new_n6377_ & new_n5590_ & new_n4946_ & new_n4049_;
  assign new_n6734_ = ~\i[1303]  & ~\i[1301]  & ~\i[1302] ;
  assign new_n6735_ = new_n6736_ ? (~new_n6774_ ^ new_n6733_) : (new_n6774_ ^ new_n6733_);
  assign new_n6736_ = new_n6737_ ? (new_n6749_ ^ new_n6764_) : (~new_n6749_ ^ new_n6764_);
  assign new_n6737_ = ~new_n6738_ & (new_n5576_ | \i[623]  | \i[986]  | \i[987] );
  assign new_n6738_ = new_n5576_ & (new_n6748_ ? new_n6739_ : (new_n6132_ ? new_n6745_ : new_n6746_));
  assign new_n6739_ = new_n6743_ ? (new_n6741_ ? new_n6740_ : ~new_n6742_) : new_n6744_;
  assign new_n6740_ = ~\i[815]  & ~\i[813]  & ~\i[814] ;
  assign new_n6741_ = ~\i[1163]  & (~\i[1162]  | (~\i[1161]  & ~\i[1160] ));
  assign new_n6742_ = \i[1639]  & \i[1638]  & \i[1636]  & \i[1637] ;
  assign new_n6743_ = \i[2439]  & \i[2438]  & \i[2436]  & \i[2437] ;
  assign new_n6744_ = (\i[1549]  | \i[1550]  | \i[1551] ) & (\i[1331]  | \i[1330] );
  assign new_n6745_ = (\i[875]  & (\i[872]  | \i[873]  | \i[874] )) ? ~new_n4379_ : ~new_n4126_;
  assign new_n6746_ = (~new_n6747_ & ~new_n5035_) | (\i[757]  & \i[758]  & \i[759]  & new_n5035_);
  assign new_n6747_ = ~\i[1215]  & ~\i[1213]  & ~\i[1214] ;
  assign new_n6748_ = ~\i[763]  & (~\i[762]  | ~\i[761] );
  assign new_n6749_ = ~new_n6763_ & (new_n6752_ | (new_n6760_ & (~new_n6761_ | new_n6750_)));
  assign new_n6750_ = (\i[1087]  & (\i[1085]  | \i[1086] )) ? ~new_n6751_ : new_n4392_;
  assign new_n6751_ = ~\i[1099]  & (~\i[1097]  | ~\i[1098]  | ~\i[1096] );
  assign new_n6752_ = ~new_n6757_ & (new_n6758_ ? new_n6753_ : (new_n6759_ ? ~new_n6756_ : new_n3373_));
  assign new_n6753_ = (new_n6754_ & new_n6755_) | (\i[871]  & ~new_n6755_ & (\i[870]  | \i[869] ));
  assign new_n6754_ = ~\i[747]  & (~\i[745]  | ~\i[746]  | ~\i[744] );
  assign new_n6755_ = ~\i[1194]  & ~\i[1195]  & (~\i[1193]  | ~\i[1192] );
  assign new_n6756_ = new_n6068_ & (\i[853]  | \i[852] );
  assign new_n6757_ = \i[851]  & \i[850]  & \i[848]  & \i[849] ;
  assign new_n6758_ = \i[859]  & (\i[857]  | \i[858]  | \i[856] );
  assign new_n6759_ = ~\i[950]  & ~\i[951]  & (~\i[949]  | ~\i[948] );
  assign new_n6760_ = new_n6757_ & ((\i[521]  & \i[522]  & \i[523] ) | ~new_n6762_ | new_n6761_);
  assign new_n6761_ = \i[1199]  & (\i[1198]  | \i[1197] );
  assign new_n6762_ = \i[1187]  & \i[1185]  & \i[1186] ;
  assign new_n6763_ = \i[2451]  & \i[2450]  & \i[2448]  & \i[2449] ;
  assign new_n6764_ = (new_n6771_ | new_n6772_ | new_n4929_) & (new_n6767_ | ~new_n4929_ | (new_n6766_ & ~new_n6765_));
  assign new_n6765_ = ~\i[2187]  & ((new_n6354_ & ~new_n4878_) | (\i[1075]  & new_n4878_ & (\i[1074]  | \i[1073] )));
  assign new_n6766_ = \i[2742]  & \i[2743]  & (~\i[2187]  | (new_n4445_ & ~new_n4662_) | (new_n3879_ & new_n4662_));
  assign new_n6767_ = (~new_n6233_ | new_n6769_) & (~\i[2743]  | ~\i[2742] ) & (new_n6768_ | ~new_n6770_ | ~new_n6769_);
  assign new_n6768_ = \i[1379]  & (\i[1378]  | \i[1377] );
  assign new_n6769_ = ~\i[2038]  & ~\i[2039]  & (~\i[2037]  | ~\i[2036] );
  assign new_n6770_ = \i[1831]  & (\i[1830]  | \i[1829] );
  assign new_n6771_ = ~new_n3447_ & ((new_n5632_ & new_n3321_) | (~\i[974]  & ~\i[975]  & new_n3368_ & ~new_n3321_));
  assign new_n6772_ = new_n3447_ & (new_n6773_ | (new_n3574_ & \i[1507] ));
  assign new_n6773_ = \i[1743]  & \i[1742]  & \i[1740]  & \i[1741] ;
  assign new_n6774_ = new_n6785_ ? new_n6775_ : ((new_n6782_ | new_n6784_ | ~new_n6786_) & (~new_n3770_ | new_n6786_));
  assign new_n6775_ = new_n5025_ ? (new_n6519_ ? new_n6780_ : new_n6781_) : new_n6776_;
  assign new_n6776_ = (new_n6777_ & (\i[1946]  | \i[1947] )) | (~\i[1946]  & ~\i[1947]  & (new_n3628_ ? ~new_n5395_ : new_n3339_));
  assign new_n6777_ = (new_n6778_ & (\i[967]  | (new_n4782_ & \i[966] ))) | (~\i[819]  & ~new_n6779_ & ~\i[967]  & (~new_n4782_ | ~\i[966] ));
  assign new_n6778_ = \i[971]  & \i[969]  & \i[970] ;
  assign new_n6779_ = \i[817]  & \i[818] ;
  assign new_n6780_ = (~\i[2631]  & new_n6202_) | (~\i[631]  & ~new_n6202_ & (~\i[630]  | ~\i[629] ));
  assign new_n6781_ = (\i[2405]  | \i[2406]  | \i[2407]  | ~new_n3350_) & (new_n3350_ | (~\i[823]  & ~\i[822] ));
  assign new_n6782_ = (new_n6783_ | ~new_n4862_) & (\i[818]  | \i[819]  | new_n4862_ | (\i[817]  & \i[816] ));
  assign new_n6783_ = \i[619]  & (\i[617]  | \i[618]  | \i[616] );
  assign new_n6784_ = new_n5421_ & (\i[2173]  | \i[2172] );
  assign new_n6785_ = ~\i[2743]  & (~\i[2742]  | (~\i[2741]  & ~\i[2740] ));
  assign new_n6786_ = ~\i[2187]  & (~\i[2185]  | ~\i[2186]  | ~\i[2184] );
  assign new_n6787_ = (new_n6788_ & new_n3273_) | (~new_n6794_ & ~new_n3273_ & (new_n5778_ | new_n6796_));
  assign new_n6788_ = (new_n6789_ & (\i[2073]  | ~new_n3302_)) | (~\i[2073]  & new_n3302_ & (\i[1291]  ? new_n6793_ : new_n6792_));
  assign new_n6789_ = new_n3889_ ? (new_n6790_ ? ~new_n6257_ : new_n6791_) : \i[1535] ;
  assign new_n6790_ = ~\i[535]  & ~\i[534]  & ~\i[532]  & ~\i[533] ;
  assign new_n6791_ = ~\i[1166]  & ~\i[1167]  & (~\i[1165]  | ~\i[1164] );
  assign new_n6792_ = (~\i[1159]  & ~new_n5411_ & new_n3993_) | (~new_n3993_ & (\i[1311]  | \i[1310] ));
  assign new_n6793_ = (new_n5139_ | new_n5215_) & (~\i[532]  | ~\i[533]  | ~\i[534]  | ~\i[535]  | ~new_n5215_);
  assign new_n6794_ = new_n5778_ & (new_n6795_ | new_n4470_) & (new_n4463_ | \i[746]  | \i[747]  | ~new_n4470_);
  assign new_n6795_ = (~new_n5173_ | new_n3404_) & (\i[2742]  | \i[2743]  | ~new_n3404_);
  assign new_n6796_ = new_n6798_ ? new_n6797_ : ((\i[634]  | \i[635]  | ~new_n3351_) & (new_n6799_ | new_n3351_));
  assign new_n6797_ = new_n4071_ ? ~new_n4094_ : (~new_n4330_ | (~\i[1496]  & ~\i[1497] ));
  assign new_n6798_ = ~\i[1495]  & ~\i[1493]  & ~\i[1494] ;
  assign new_n6799_ = ~\i[527]  & ~\i[526]  & ~\i[524]  & ~\i[525] ;
  assign new_n6800_ = new_n6801_ ? (new_n6889_ ^ new_n6903_) : (~new_n6889_ ^ new_n6903_);
  assign new_n6801_ = new_n6802_ ? (~new_n6840_ ^ new_n6877_) : (new_n6840_ ^ new_n6877_);
  assign new_n6802_ = new_n6803_ ? (~new_n6809_ ^ new_n6823_) : (new_n6809_ ^ new_n6823_);
  assign new_n6803_ = (~\i[1138]  & ~\i[1139]  & new_n6804_ & ~\i[1137] ) | (~new_n5567_ & (\i[1137]  | \i[1138]  | \i[1139] ));
  assign new_n6804_ = (\i[2258]  & \i[2259] ) ? ~new_n5030_ : new_n6805_;
  assign new_n6805_ = (new_n6806_ & ~new_n6808_) | (~new_n3447_ & \i[1710]  & \i[1711]  & new_n6808_);
  assign new_n6806_ = new_n6807_ ? ~new_n4162_ : ~\i[1519] ;
  assign new_n6807_ = \i[1403]  & (\i[1401]  | \i[1402]  | \i[1400] );
  assign new_n6808_ = ~\i[1523]  & (~\i[1522]  | (~\i[1521]  & ~\i[1520] ));
  assign new_n6809_ = new_n3502_ ? new_n6810_ : ((~new_n6817_ & new_n5747_) | (~new_n6820_ & ~new_n6821_ & ~new_n5747_));
  assign new_n6810_ = ~new_n6811_ & (new_n5007_ | ((new_n6815_ | new_n3988_) & (new_n4257_ | ~new_n3342_ | ~new_n3988_)));
  assign new_n6811_ = ~new_n6812_ & new_n5007_ & (new_n6814_ | (new_n6447_ & (\i[1061]  | ~new_n4029_)));
  assign new_n6812_ = new_n6814_ & ((new_n6813_ & ~new_n6204_) | (\i[2431]  & new_n6204_ & (\i[2428]  | ~new_n5407_)));
  assign new_n6813_ = ~\i[1303]  & (~\i[1301]  | ~\i[1302]  | ~\i[1300] );
  assign new_n6814_ = \i[851]  & (\i[850]  | (\i[849]  & \i[848] ));
  assign new_n6815_ = (~\i[2266]  & ~\i[2267] ) ? new_n3568_ : ~new_n6816_;
  assign new_n6816_ = \i[626]  & \i[627]  & (\i[625]  | \i[624] );
  assign new_n6817_ = (~\i[1654]  & ~\i[1655]  & new_n6818_ & ~\i[1653] ) | (~new_n6400_ & (\i[1653]  | \i[1654]  | \i[1655] ));
  assign new_n6818_ = (~\i[2042]  | ~\i[2043]  | new_n6819_) & (~\i[1418]  | ~\i[1419]  | ~new_n6819_);
  assign new_n6819_ = ~\i[1639]  & ~\i[1637]  & ~\i[1638] ;
  assign new_n6820_ = \i[615]  & \i[614]  & new_n3515_ & new_n6198_;
  assign new_n6821_ = new_n6822_ & (~\i[1492]  | ~\i[1493]  | ~\i[1494]  | ~\i[1495] );
  assign new_n6822_ = \i[1079]  & (~\i[614]  | ~\i[615] ) & (\i[1078]  | (\i[1077]  & \i[1076] ));
  assign new_n6823_ = new_n6839_ ? new_n6824_ : ((~new_n6834_ & new_n3375_) | (~new_n6837_ & ~new_n6838_ & ~new_n3375_));
  assign new_n6824_ = (~new_n6829_ & ~new_n6832_ & new_n6833_) | (~new_n6833_ & (new_n6827_ | new_n6825_));
  assign new_n6825_ = new_n5750_ & (new_n5842_ ? ~new_n6826_ : (\i[1035]  | (\i[1033]  & \i[1034] )));
  assign new_n6826_ = ~\i[1094]  & ~\i[1095]  & (~\i[1093]  | ~\i[1092] );
  assign new_n6827_ = ~new_n5750_ & ((~new_n6828_ & new_n5646_) | (~\i[1929]  & ~\i[1930]  & ~\i[1931]  & ~new_n5646_));
  assign new_n6828_ = new_n4781_ & (\i[965]  | \i[964] );
  assign new_n6829_ = new_n6831_ & ((new_n4710_ & (new_n3667_ | \i[1070]  | \i[1071] )) | (~\i[1070]  & ~\i[1071]  & new_n6830_ & ~new_n3667_));
  assign new_n6830_ = ~\i[1082]  & ~\i[1083]  & (~\i[1081]  | ~\i[1080] );
  assign new_n6831_ = ~\i[1206]  & ~\i[1207]  & (~\i[1205]  | ~\i[1204] );
  assign new_n6832_ = ~new_n6831_ & ~\i[1651]  & (~\i[1650]  | (~\i[1648]  & ~\i[1649] ));
  assign new_n6833_ = ~\i[982]  & ~\i[983]  & (~\i[981]  | ~\i[980] );
  assign new_n6834_ = ~new_n6836_ & (~new_n6835_ | (~\i[2052]  & ~\i[2053]  & ~\i[2054] ));
  assign new_n6835_ = ~new_n5781_ & \i[2055]  & (~\i[1711]  | ~\i[1710] );
  assign new_n6836_ = \i[1711]  & \i[1710]  & new_n3588_ & new_n3645_;
  assign new_n6837_ = ~\i[1194]  & ~\i[1195]  & \i[963]  & (\i[962]  | \i[961] );
  assign new_n6838_ = \i[987]  & \i[986]  & (\i[1194]  | \i[1195] ) & (\i[984]  | \i[985] );
  assign new_n6839_ = ~\i[639]  & ~\i[638]  & ~\i[636]  & ~\i[637] ;
  assign new_n6840_ = new_n6841_ ? (~new_n6857_ ^ new_n6865_) : (new_n6857_ ^ new_n6865_);
  assign new_n6841_ = ~new_n6842_ & (new_n4272_ | ((new_n6849_ | new_n4371_) & (new_n6847_ | new_n6853_ | ~new_n4371_)));
  assign new_n6842_ = new_n4272_ & (new_n4884_ ? new_n6843_ : (new_n3470_ ? new_n4990_ : new_n6846_));
  assign new_n6843_ = (new_n6844_ | ~new_n4414_ | (~\i[732]  & ~\i[733] )) & (new_n6845_ | new_n4701_ | (new_n4414_ & (\i[732]  | \i[733] )));
  assign new_n6844_ = (\i[2518]  | \i[2519]  | new_n3754_) & (\i[646]  | \i[647]  | ~new_n3754_);
  assign new_n6845_ = ~\i[2186]  & ~\i[2187]  & (~\i[2185]  | ~\i[2184] );
  assign new_n6846_ = ~new_n4094_ & (~\i[1931]  | (~\i[1929]  & ~\i[1930] ));
  assign new_n6847_ = new_n6848_ & (~new_n3376_ | (\i[1933]  & \i[1934]  & \i[1935] ));
  assign new_n6848_ = ~\i[1519]  & (~\i[1517]  | ~\i[1518]  | ~\i[1516] );
  assign new_n6849_ = new_n3477_ ? new_n6852_ : new_n6850_;
  assign new_n6850_ = new_n6851_ ? (~\i[2323]  | (~\i[2321]  & ~\i[2322] )) : new_n6225_;
  assign new_n6851_ = ~\i[943]  & ~\i[941]  & ~\i[942] ;
  assign new_n6852_ = (~\i[713]  & ~\i[714]  & ~\i[715]  & new_n3368_) | (~new_n5719_ & ~new_n3368_);
  assign new_n6853_ = ~new_n6848_ & (new_n6855_ ? (\i[1847]  | new_n6854_) : new_n6856_);
  assign new_n6854_ = \i[1846]  & (\i[1845]  | \i[1844] );
  assign new_n6855_ = ~\i[1411]  & (~\i[1410]  | ~\i[1409] );
  assign new_n6856_ = ~\i[1827]  & (~\i[1825]  | ~\i[1826]  | ~\i[1824] );
  assign new_n6857_ = new_n6864_ ? (new_n6762_ ? new_n6858_ : new_n6860_) : new_n6673_;
  assign new_n6858_ = (~new_n6859_ | ~new_n4257_ | ~new_n3889_) & (new_n3889_ | (\i[1315]  & (\i[1313]  | \i[1314] )));
  assign new_n6859_ = \i[2171]  & \i[2170]  & \i[2168]  & \i[2169] ;
  assign new_n6860_ = new_n5930_ ? new_n6863_ : ((~new_n6862_ | ~new_n4901_) & (new_n6861_ | \i[2055]  | new_n4901_));
  assign new_n6861_ = \i[2054]  & \i[2052]  & \i[2053] ;
  assign new_n6862_ = ~\i[2194]  & ~\i[2195]  & (~\i[2193]  | ~\i[2192] );
  assign new_n6863_ = ~\i[1219]  & ~\i[1218]  & ~\i[1216]  & ~\i[1217] ;
  assign new_n6864_ = ~\i[1107]  & (~\i[1106]  | (~\i[1105]  & ~\i[1104] ));
  assign new_n6865_ = (new_n6871_ | new_n6876_ | ~new_n6225_) & (new_n6225_ | (new_n5079_ ? new_n6874_ : new_n6866_));
  assign new_n6866_ = (\i[1973]  & \i[1974]  & \i[1975] ) ? (new_n6869_ | new_n6870_) : new_n6867_;
  assign new_n6867_ = (~new_n6868_ & (~\i[1269]  | ~\i[1270]  | ~\i[1271] )) | (~new_n3387_ & \i[1269]  & \i[1270]  & \i[1271] );
  assign new_n6868_ = ~\i[2263]  & (~\i[2261]  | ~\i[2262]  | ~\i[2260] );
  assign new_n6869_ = ~\i[2605]  & ~\i[2606]  & ~\i[2607]  & (\i[1059]  | (\i[1058]  & \i[1057] ));
  assign new_n6870_ = ~\i[1059]  & (~\i[1057]  | ~\i[1058] ) & (\i[538]  | \i[539]  | \i[537] );
  assign new_n6871_ = new_n5078_ & ((~new_n6872_ & ~new_n3452_) | (~new_n4402_ & ~new_n6873_ & new_n3452_));
  assign new_n6872_ = new_n3499_ & ~\i[1090]  & ~\i[1091] ;
  assign new_n6873_ = ~\i[751]  & (~\i[749]  | ~\i[750]  | ~\i[748] );
  assign new_n6874_ = new_n6875_ ? new_n3534_ : (~new_n3265_ | (~\i[1494]  & ~\i[1495] ));
  assign new_n6875_ = \i[742]  & \i[743]  & (\i[741]  | \i[740] );
  assign new_n6876_ = ~new_n5078_ & ((new_n3417_ & new_n3477_) | (new_n3432_ & new_n3373_ & ~new_n3477_));
  assign new_n6877_ = new_n6888_ ? new_n6881_ : ((~new_n6886_ & new_n5134_) | (~new_n6883_ & ~new_n6878_ & ~new_n5134_));
  assign new_n6878_ = new_n6879_ & (new_n4470_ ? new_n5693_ : ~new_n6880_);
  assign new_n6879_ = ~\i[2318]  & ~\i[2319]  & (~\i[2317]  | ~\i[2316] );
  assign new_n6880_ = ~\i[650]  & ~\i[651]  & (~\i[649]  | ~\i[648] );
  assign new_n6881_ = new_n5404_ ? ~new_n4288_ : new_n6882_;
  assign new_n6882_ = new_n4759_ ? ((\i[1058]  | \i[1059] ) & (~\i[939]  | ~\i[938] )) : \i[1079] ;
  assign new_n6883_ = ~new_n6879_ & ((new_n6885_ & \i[829] ) ? new_n4268_ : ~new_n6884_);
  assign new_n6884_ = \i[1279]  & (\i[1278]  | (\i[1277]  & \i[1276] ));
  assign new_n6885_ = \i[830]  & \i[831] ;
  assign new_n6886_ = (~new_n6887_ & ~\i[2647]  & new_n6135_) | (~new_n6135_ & (new_n6680_ | new_n3451_));
  assign new_n6887_ = \i[1155]  & \i[1153]  & \i[1154] ;
  assign new_n6888_ = \i[711]  & \i[710]  & \i[708]  & \i[709] ;
  assign new_n6889_ = new_n6785_ ? new_n6890_ : (new_n5626_ ? ~new_n6895_ : ~new_n6900_);
  assign new_n6890_ = (~new_n6893_ | new_n6891_) & (~new_n6894_ | (new_n4463_ ? ~\i[1507]  : new_n3471_));
  assign new_n6891_ = ~new_n5539_ & (new_n6892_ ? ~new_n4976_ : (\i[1183]  | (new_n3720_ & \i[1180] )));
  assign new_n6892_ = new_n3849_ & (~\i[2753]  | ~\i[2752] );
  assign new_n6893_ = new_n4437_ & (new_n5695_ | ~new_n5539_ | (~\i[491]  & (~\i[489]  | ~\i[490] )));
  assign new_n6894_ = ~new_n4437_ & (~\i[2855]  | (~\i[2852]  & ~\i[2853]  & ~\i[2854] ));
  assign new_n6895_ = ~new_n6896_ & (~new_n6899_ | ~new_n4315_ | (\i[1851]  & (\i[1849]  | \i[1850] )));
  assign new_n6896_ = ~new_n4315_ & ((new_n6898_ & new_n6897_) | (~\i[1603]  & ~new_n6897_ & (~\i[1602]  | ~\i[1601] )));
  assign new_n6897_ = ~\i[1987]  & (~\i[1985]  | ~\i[1986]  | ~\i[1984] );
  assign new_n6898_ = ~\i[2498]  & ~\i[2499]  & (~\i[2497]  | ~\i[2496] );
  assign new_n6899_ = ~\i[1494]  & ~\i[1495]  & (~\i[1493]  | ~\i[1492] );
  assign new_n6900_ = (~new_n4659_ | (new_n5006_ ? new_n3342_ : new_n4431_)) & (new_n6902_ | ~new_n6901_ | new_n4659_);
  assign new_n6901_ = ~\i[1098]  & ~\i[1099]  & (~\i[1097]  | ~\i[1096] );
  assign new_n6902_ = ~\i[2071]  & ~\i[2069]  & ~\i[2070] ;
  assign new_n6903_ = (new_n6908_ | new_n6905_ | new_n6377_) & (~new_n6377_ | (~new_n6904_ & (new_n6911_ | new_n5590_)));
  assign new_n6904_ = new_n5590_ & (~new_n4946_ | ~new_n4049_ | ~new_n6734_) & (new_n4353_ | ~new_n4785_ | new_n6734_);
  assign new_n6905_ = ~new_n6734_ & new_n6907_ & (new_n3227_ ? (~\i[955]  | ~new_n3249_) : ~new_n6906_);
  assign new_n6906_ = \i[2747]  & \i[2746]  & \i[2744]  & \i[2745] ;
  assign new_n6907_ = \i[1083]  & (\i[1082]  | \i[1081] );
  assign new_n6908_ = new_n6734_ & ((new_n4939_ & new_n4180_ & new_n6909_) | (~new_n3499_ & ~new_n6910_ & ~new_n6909_));
  assign new_n6909_ = \i[1523]  & \i[1521]  & \i[1522] ;
  assign new_n6910_ = \i[815]  & \i[814]  & \i[812]  & \i[813] ;
  assign new_n6911_ = new_n5065_ ? new_n6387_ : ~new_n6912_;
  assign new_n6912_ = ~\i[2090]  & ~\i[2091]  & (~\i[2089]  | ~\i[2088] );
  assign new_n6913_ = new_n6932_ ? new_n6914_ : ((new_n6927_ | new_n6923_ | ~new_n6808_) & (new_n6928_ | new_n6808_));
  assign new_n6914_ = new_n6922_ ? ((new_n6920_ & ~new_n3729_) | (~new_n5665_ & new_n4078_ & new_n3729_)) : new_n6915_;
  assign new_n6915_ = (new_n6917_ | new_n6919_ | new_n4716_) & (new_n6916_ | new_n6918_ | ~new_n4716_);
  assign new_n6916_ = \i[963]  & new_n3796_ & \i[962] ;
  assign new_n6917_ = ~\i[2399]  & ~\i[2398]  & new_n4755_ & (~\i[2609]  | ~\i[2608] );
  assign new_n6918_ = ~\i[771]  & ~\i[770]  & (~\i[962]  | ~\i[963] ) & (~\i[768]  | ~\i[769] );
  assign new_n6919_ = \i[2647]  & (\i[2398]  | \i[2399] ) & (\i[2646]  | (\i[2645]  & \i[2644] ));
  assign new_n6920_ = ~new_n6921_ & (~\i[1989]  | ~\i[1990]  | ~\i[1991] );
  assign new_n6921_ = \i[878]  & \i[879]  & (\i[877]  | \i[876] );
  assign new_n6922_ = ~\i[2411]  & (~\i[2410]  | ~\i[2409] );
  assign new_n6923_ = new_n4217_ & (new_n6924_ | (~new_n6925_ & ~\i[2509]  & new_n3796_));
  assign new_n6924_ = new_n6925_ & \i[1059]  & (\i[1058]  | \i[1057] );
  assign new_n6925_ = new_n6926_ & (\i[2729]  | \i[2728] );
  assign new_n6926_ = \i[2730]  & \i[2731] ;
  assign new_n6927_ = ~new_n4819_ & ~new_n4217_ & \i[1827]  & (\i[1826]  | \i[1825]  | \i[1824] );
  assign new_n6928_ = (~new_n5654_ & new_n5420_ & new_n6929_) | (~new_n6929_ & (~new_n6931_ | ~new_n6930_));
  assign new_n6929_ = ~\i[1743]  & (~\i[1742]  | (~\i[1741]  & ~\i[1740] ));
  assign new_n6930_ = ~\i[2443]  & (~\i[2442]  | ~\i[2441] );
  assign new_n6931_ = \i[1835]  & \i[1834]  & \i[1832]  & \i[1833] ;
  assign new_n6932_ = \i[2403]  & (\i[2402]  | \i[2401] );
  assign new_n6933_ = new_n6934_ ? (~new_n6960_ ^ new_n6977_) : (new_n6960_ ^ new_n6977_);
  assign new_n6934_ = new_n6935_ ? (new_n6946_ ^ new_n6952_) : (~new_n6946_ ^ new_n6952_);
  assign new_n6935_ = new_n4434_ ? new_n6936_ : ((~new_n6941_ & ~new_n3644_) | (~new_n6945_ & new_n4789_ & new_n3644_));
  assign new_n6936_ = new_n5693_ ? ((new_n6940_ & ~new_n6807_) | (new_n5007_ & new_n4299_ & new_n6807_)) : new_n6937_;
  assign new_n6937_ = ~new_n6938_ & (~new_n4192_ | ((~\i[503]  | ~new_n3873_) & (new_n6939_ | ~\i[1383]  | new_n3873_)));
  assign new_n6938_ = ~new_n4192_ & (new_n4055_ | ~new_n5678_) & (\i[1061]  | \i[1062]  | \i[1063]  | new_n5678_);
  assign new_n6939_ = ~\i[1382]  & ~\i[1380]  & ~\i[1381] ;
  assign new_n6940_ = \i[1943]  & (\i[1942]  | (\i[1941]  & \i[1940] ));
  assign new_n6941_ = (new_n5186_ | ~new_n6944_ | (\i[1195]  & \i[1194] )) & (new_n6943_ | new_n6942_ | new_n6944_);
  assign new_n6942_ = new_n6907_ & (\i[751]  | (\i[749]  & \i[750] ));
  assign new_n6943_ = ~\i[751]  & ~\i[1090]  & ~\i[1091]  & (~\i[750]  | ~\i[749] );
  assign new_n6944_ = \i[2287]  & (\i[2286]  | \i[2285] );
  assign new_n6945_ = ~new_n3675_ & new_n3660_;
  assign new_n6946_ = new_n6864_ ? ((new_n6950_ | new_n6949_ | ~new_n3446_) & (new_n6947_ | new_n3446_)) : new_n5925_;
  assign new_n6947_ = (~new_n3892_ | ~new_n6828_ | new_n6400_) & (~new_n6400_ | (new_n3308_ ? ~new_n6948_ : ~new_n4396_));
  assign new_n6948_ = ~\i[1087]  & ~\i[1086]  & ~\i[1084]  & ~\i[1085] ;
  assign new_n6949_ = new_n3400_ & (new_n3735_ | (\i[1725]  & \i[1726]  & \i[1727] ));
  assign new_n6950_ = ~new_n3400_ & ((~\i[1302]  & ~\i[1303] ) ? ~new_n6951_ : ~new_n6435_);
  assign new_n6951_ = ~\i[1763]  & ~\i[1762]  & ~\i[1760]  & ~\i[1761] ;
  assign new_n6952_ = new_n6959_ ? (new_n6534_ ? ~new_n6953_ : ~new_n6958_) : new_n6955_;
  assign new_n6953_ = (new_n6954_ | new_n5395_) & (new_n5483_ | new_n6385_ | ~new_n5395_);
  assign new_n6954_ = new_n5675_ & (\i[963]  | (\i[962]  & (\i[961]  | \i[960] )));
  assign new_n6955_ = new_n4859_ ? ((new_n6957_ & new_n6472_) | (~new_n6956_ & new_n3556_ & ~new_n6472_)) : ~new_n3555_;
  assign new_n6956_ = ~\i[2163]  & ~\i[2162]  & ~\i[2160]  & ~\i[2161] ;
  assign new_n6957_ = \i[2067]  & \i[2522]  & \i[2523]  & (\i[2521]  | \i[2520] );
  assign new_n6958_ = ~\i[1325]  & ~\i[1326]  & ~\i[1327]  & (new_n5134_ | new_n3461_);
  assign new_n6959_ = ~\i[643]  & (~\i[641]  | ~\i[642]  | ~\i[640] );
  assign new_n6960_ = new_n4960_ ? new_n6961_ : (new_n6974_ | (~new_n6969_ & ~new_n6673_));
  assign new_n6961_ = (new_n6965_ & new_n5568_) | (~new_n6962_ & ~new_n6967_ & ~new_n5568_);
  assign new_n6962_ = new_n6963_ & (new_n3239_ | \i[2715]  | (\i[2714]  & (\i[2712]  | \i[2713] )));
  assign new_n6963_ = ~new_n6964_ & (~\i[1527]  | ~new_n3239_ | (~\i[1524]  & ~\i[1525]  & ~\i[1526] ));
  assign new_n6964_ = ~\i[1427]  & (~\i[1426]  | (~\i[1425]  & ~\i[1424] ));
  assign new_n6965_ = (~new_n6830_ & ~new_n6966_ & new_n4818_) | (~new_n4818_ & (\i[1187]  | new_n5804_));
  assign new_n6966_ = ~\i[971]  & (~\i[969]  | ~\i[970]  | ~\i[968] );
  assign new_n6967_ = new_n6964_ & ((new_n6968_ & ~new_n3899_) | (~\i[1439]  & new_n3899_ & (~\i[1438]  | ~\i[1437] )));
  assign new_n6968_ = \i[2087]  & \i[2086]  & \i[2084]  & \i[2085] ;
  assign new_n6969_ = new_n6973_ ? new_n6970_ : (new_n6972_ ? \i[2439]  : new_n6912_);
  assign new_n6970_ = new_n6971_ ? ~new_n5721_ : new_n6443_;
  assign new_n6971_ = ~\i[1423]  & (~\i[1422]  | (~\i[1421]  & ~\i[1420] ));
  assign new_n6972_ = ~\i[763]  & (~\i[761]  | ~\i[762]  | ~\i[760] );
  assign new_n6973_ = \i[963]  & \i[961]  & \i[962] ;
  assign new_n6974_ = new_n6673_ & (new_n4695_ | ~new_n4380_ | ~new_n6975_) & (new_n6976_ | new_n3741_ | new_n6975_);
  assign new_n6975_ = ~\i[1095]  & ~\i[1094]  & ~\i[1092]  & ~\i[1093] ;
  assign new_n6976_ = ~\i[979]  & (~\i[977]  | ~\i[978]  | ~\i[976] );
  assign new_n6977_ = new_n3996_ ? ((new_n6987_ | new_n6988_ | ~new_n6534_) & (new_n6983_ | new_n6534_)) : new_n6978_;
  assign new_n6978_ = ~new_n6979_ & (new_n3726_ | new_n6980_ | ~new_n6519_ | ~new_n3568_);
  assign new_n6979_ = new_n6980_ & (new_n6982_ | new_n3405_) & (new_n6981_ | new_n5443_ | \i[607]  | ~new_n3405_);
  assign new_n6980_ = ~\i[974]  & ~\i[975]  & (~\i[973]  | ~\i[972] );
  assign new_n6981_ = \i[606]  & \i[604]  & \i[605] ;
  assign new_n6982_ = ~\i[987]  & ~\i[986]  & ~\i[984]  & ~\i[985] ;
  assign new_n6983_ = \i[639]  ? new_n6984_ : (new_n6975_ ? new_n6986_ : ~new_n6320_);
  assign new_n6984_ = (~new_n6985_ | ~new_n3760_) & (~\i[2499]  | new_n3760_ | (~\i[2498]  & (~\i[2496]  | ~\i[2497] )));
  assign new_n6985_ = \i[850]  & \i[851]  & (\i[849]  | \i[848] );
  assign new_n6986_ = \i[995]  & (\i[994]  | \i[993] );
  assign new_n6987_ = ~new_n4060_ & ((~new_n3400_ & ~new_n6839_) | (~\i[1093]  & ~\i[1094]  & ~\i[1095]  & new_n6839_));
  assign new_n6988_ = new_n4060_ & (new_n4231_ | new_n3615_) & (\i[1061]  | \i[1062]  | \i[1063]  | ~new_n3615_);
  assign new_n6989_ = (new_n6997_ | (\i[419]  ? ~new_n6996_ : new_n6990_)) & (new_n6763_ | ~new_n6992_ | ~new_n6997_);
  assign new_n6990_ = ~new_n6991_ & ((~\i[1030]  & ~\i[1031] ) | new_n4667_ | ~new_n4273_);
  assign new_n6991_ = ~new_n4273_ & new_n6171_ & (\i[411]  | (\i[408]  & \i[409]  & \i[410] ));
  assign new_n6992_ = (~new_n3539_ | (~\i[547]  & (~\i[545]  | ~\i[546] ))) & (new_n6995_ | new_n6993_ | \i[547]  | (\i[545]  & \i[546] ));
  assign new_n6993_ = ~\i[2187]  & ~\i[2186]  & ~new_n6994_ & ~\i[2185] ;
  assign new_n6994_ = ~\i[2847]  & ~\i[2845]  & ~\i[2846] ;
  assign new_n6995_ = \i[415]  & \i[414]  & \i[413]  & new_n6994_ & \i[412] ;
  assign new_n6996_ = new_n3437_ & (\i[2415]  | \i[2414] );
  assign new_n6997_ = \i[1942]  & \i[1943]  & (\i[1941]  | \i[1940] );
  assign new_n6998_ = (~new_n7004_ & ~new_n7007_ & ~new_n6198_) | (new_n6198_ & (new_n6982_ ? new_n7003_ : new_n6999_));
  assign new_n6999_ = ~new_n7000_ & (~new_n7002_ | (~\i[1311]  & (~\i[1308]  | ~\i[1309]  | ~\i[1310] )));
  assign new_n7000_ = \i[2603]  & \i[2602]  & \i[2601]  & ~new_n7001_ & ~new_n3858_;
  assign new_n7001_ = \i[1189]  & new_n3499_ & \i[1188] ;
  assign new_n7002_ = new_n3858_ & ~\i[1439]  & ~\i[1438]  & ~\i[1436]  & ~\i[1437] ;
  assign new_n7003_ = new_n6799_ ? ~new_n6863_ : (new_n3415_ ? new_n4717_ : ~new_n4396_);
  assign new_n7004_ = ~new_n7006_ & ~new_n7005_ & new_n4884_ & (~new_n4788_ | (\i[1078]  & \i[1079] ));
  assign new_n7005_ = \i[1079]  & \i[1078]  & (\i[1503]  | (\i[1501]  & \i[1502] ));
  assign new_n7006_ = ~\i[1207]  & ~\i[1205]  & ~\i[1206] ;
  assign new_n7007_ = ~new_n4884_ & ~new_n5843_ & ~new_n7008_ & (\i[955]  | (\i[1494]  & \i[1495] ));
  assign new_n7008_ = \i[955]  & (~\i[631]  | (~\i[629]  & ~\i[630]  & ~\i[628] ));
  assign new_n7009_ = new_n6073_ ? new_n7019_ : ((new_n7017_ | new_n7013_ | ~new_n6708_) & (new_n7010_ | new_n6708_));
  assign new_n7010_ = new_n6427_ ? ~new_n7012_ : ~new_n7011_;
  assign new_n7011_ = ~new_n4424_ & \i[1223]  & (\i[1222]  | (\i[1220]  & \i[1221] ));
  assign new_n7012_ = new_n4175_ & ~\i[1551]  & ~\i[1550]  & ~\i[1548]  & ~\i[1549] ;
  assign new_n7013_ = ~new_n7014_ & new_n3445_;
  assign new_n7014_ = new_n7015_ ? (~\i[1331]  & (~\i[1328]  | ~\i[1329]  | ~\i[1330] )) : ~new_n7016_;
  assign new_n7015_ = ~\i[762]  & ~\i[763]  & (~\i[761]  | ~\i[760] );
  assign new_n7016_ = ~\i[987]  & ~\i[985]  & ~\i[986] ;
  assign new_n7017_ = ~new_n3445_ & ((~\i[1218]  & ~\i[1219]  & new_n6135_) | (~new_n7018_ & ~new_n6135_));
  assign new_n7018_ = new_n4068_ & (~\i[1201]  | ~\i[1200] );
  assign new_n7019_ = new_n7023_ ? ((new_n7020_ | ~new_n3436_) & (new_n3881_ | ~new_n4020_ | new_n3436_)) : new_n7021_;
  assign new_n7020_ = new_n3898_ & ~\i[870]  & ~\i[871] ;
  assign new_n7021_ = (new_n3663_ | new_n6297_ | \i[1175] ) & (\i[1079]  | ~new_n7022_ | ~\i[1175] );
  assign new_n7022_ = ~\i[1099]  & ~\i[1098]  & ~\i[1096]  & ~\i[1097] ;
  assign new_n7023_ = ~\i[1191]  & (~\i[1189]  | ~\i[1190]  | ~\i[1188] );
  assign new_n7024_ = new_n4701_ ? new_n7029_ : ((new_n7025_ | new_n4958_ | ~new_n4190_) & (new_n7026_ | new_n4190_));
  assign new_n7025_ = (~new_n3854_ | new_n5733_) & (\i[2622]  | \i[2623]  | ~new_n5733_ | (\i[2621]  & \i[2620] ));
  assign new_n7026_ = new_n3278_ ? (new_n7028_ ? new_n6459_ : ~\i[1331] ) : new_n7027_;
  assign new_n7027_ = (~new_n4981_ | \i[1851] ) & (~\i[692]  | ~\i[693]  | ~\i[694]  | ~\i[695]  | ~\i[1851] );
  assign new_n7028_ = ~\i[1419]  & ~\i[1418]  & ~\i[1416]  & ~\i[1417] ;
  assign new_n7029_ = (new_n3496_ | new_n5240_ | new_n5483_ | ~new_n7032_) & (new_n7030_ | new_n7032_);
  assign new_n7030_ = (~new_n7031_ | ~new_n3401_) & (~\i[2762]  | ~\i[2763]  | new_n3401_ | new_n6986_ | ~\i[2761] );
  assign new_n7031_ = ~\i[2091]  & ~\i[2090]  & ~\i[2088]  & ~\i[2089] ;
  assign new_n7032_ = ~\i[1319]  & ~\i[1318]  & ~\i[1316]  & ~\i[1317] ;
  assign \o[36]  = new_n7034_ ? (new_n7035_ ^ new_n7036_) : (~new_n7035_ ^ new_n7036_);
  assign new_n7034_ = ~new_n6644_ & ~new_n7024_;
  assign new_n7035_ = (~new_n6998_ & ~new_n7009_) | (new_n6645_ & (~new_n6998_ | ~new_n7009_));
  assign new_n7036_ = new_n7037_ ? (~new_n7038_ ^ new_n7129_) : (new_n7038_ ^ new_n7129_);
  assign new_n7037_ = (~new_n6933_ & new_n6989_) | (new_n6646_ & (~new_n6933_ | new_n6989_));
  assign new_n7038_ = new_n7039_ ? (new_n7040_ ^ new_n7122_) : (~new_n7040_ ^ new_n7122_);
  assign new_n7039_ = (~new_n6913_ & new_n6800_) | (new_n6647_ & (~new_n6913_ | new_n6800_));
  assign new_n7040_ = new_n7041_ ? (new_n7042_ ^ new_n7101_) : (~new_n7042_ ^ new_n7101_);
  assign new_n7041_ = (~new_n6787_ & new_n6735_) | (new_n6648_ & (~new_n6787_ | new_n6735_));
  assign new_n7042_ = new_n7043_ ? (new_n7044_ ^ new_n7082_) : (~new_n7044_ ^ new_n7082_);
  assign new_n7043_ = (new_n6694_ & new_n6733_) | (~new_n6649_ & (new_n6694_ | new_n6733_));
  assign new_n7044_ = new_n7045_ ? (new_n7066_ ^ new_n7067_) : (~new_n7066_ ^ new_n7067_);
  assign new_n7045_ = new_n7046_ ? (new_n7052_ ^ new_n7060_) : (~new_n7052_ ^ new_n7060_);
  assign new_n7046_ = ~new_n6651_ & (new_n3624_ | (~new_n7047_ & ~new_n3376_) | (~new_n7049_ & new_n3376_));
  assign new_n7047_ = (new_n7048_ | new_n4352_) & (~new_n3385_ | ~new_n3502_ | ~new_n4352_);
  assign new_n7048_ = (~new_n6662_ & ~new_n6663_) | (~\i[1271]  & new_n6663_ & (~\i[1270]  | ~\i[1269] ));
  assign new_n7049_ = (new_n7050_ | new_n7051_ | new_n6665_) & (~new_n6665_ | (~new_n6664_ & (~new_n4148_ | ~new_n3323_)));
  assign new_n7050_ = ~\i[1107]  & (~\i[1105]  | ~\i[1106]  | ~\i[1104] );
  assign new_n7051_ = ~\i[1195]  & (~\i[1194]  | ~\i[1193] );
  assign new_n7052_ = new_n4701_ ? new_n7053_ : (~new_n4190_ | (~new_n7057_ & ~new_n7059_));
  assign new_n7053_ = new_n7032_ ? new_n7054_ : ((new_n7056_ | ~new_n3401_) & (~new_n3609_ | ~new_n6986_ | new_n3401_));
  assign new_n7054_ = new_n3496_ ? (new_n5013_ ? ~new_n5842_ : ~new_n4316_) : new_n7055_;
  assign new_n7055_ = new_n5240_ ? new_n6708_ : ~new_n5483_;
  assign new_n7056_ = new_n7031_ ? new_n5133_ : ~\i[2255] ;
  assign new_n7057_ = new_n4958_ & (new_n4689_ | new_n7058_) & (\i[1333]  | \i[1334]  | \i[1335]  | ~new_n7058_);
  assign new_n7058_ = ~\i[2155]  & ~\i[2154]  & ~\i[2152]  & ~\i[2153] ;
  assign new_n7059_ = ~new_n4958_ & new_n5733_ & ((\i[2620]  & \i[2621] ) | \i[2623]  | \i[2622] );
  assign new_n7060_ = new_n6073_ ? new_n7061_ : ((~new_n7013_ & new_n6708_) | (~new_n7064_ & ~new_n7065_ & ~new_n6708_));
  assign new_n7061_ = (new_n7062_ | new_n7023_) & (new_n3436_ | ~new_n3351_ | ~new_n3881_ | ~new_n7023_);
  assign new_n7062_ = (~new_n6948_ | ~new_n6297_ | \i[1175] ) & (new_n7022_ | \i[1652]  | ~new_n7063_ | ~\i[1175] );
  assign new_n7063_ = ~\i[1655]  & ~\i[1653]  & ~\i[1654] ;
  assign new_n7064_ = ~new_n6427_ & new_n4424_ & (\i[1219]  | (\i[1216]  & \i[1217]  & \i[1218] ));
  assign new_n7065_ = new_n6427_ & ~\i[1551]  & ~\i[1550]  & ~\i[1549]  & ~new_n4175_ & ~\i[1548] ;
  assign new_n7066_ = (~new_n6666_ & ~new_n6685_) | (~new_n6650_ & (~new_n6666_ | ~new_n6685_));
  assign new_n7067_ = new_n7068_ ^ new_n7075_;
  assign new_n7068_ = (new_n7069_ & new_n4380_) | (~new_n7073_ & ~new_n4380_ & (new_n6684_ | new_n7072_));
  assign new_n7069_ = (new_n7070_ | ~new_n6669_) & (~new_n3467_ | ~new_n3889_ | ~new_n6673_ | new_n6669_);
  assign new_n7070_ = (new_n6675_ | new_n6677_) & (new_n4018_ | new_n7071_ | ~new_n6677_);
  assign new_n7071_ = ~\i[1107]  & ~\i[1106]  & ~\i[1104]  & ~\i[1105] ;
  assign new_n7072_ = (~new_n3384_ | ~new_n4392_ | new_n6680_) & (~new_n6680_ | (new_n6679_ ? ~new_n3494_ : new_n6314_));
  assign new_n7073_ = new_n6684_ & new_n3318_ & ~new_n6682_ & ~new_n7074_;
  assign new_n7074_ = \i[531]  & \i[529]  & \i[530] ;
  assign new_n7075_ = (~new_n5698_ | (new_n6691_ ? new_n7076_ : new_n7077_)) & (new_n7078_ | new_n7081_ | new_n5698_);
  assign new_n7076_ = (new_n5031_ | ~new_n3618_ | ~new_n5126_) & (new_n5126_ | (new_n3555_ ? ~new_n6690_ : ~new_n5006_));
  assign new_n7077_ = (new_n6709_ | ~new_n4190_ | new_n3376_) & (~new_n3376_ | (new_n3400_ ? ~new_n3342_ : new_n6864_));
  assign new_n7078_ = new_n3998_ & (new_n5842_ ? (new_n3462_ ? ~new_n4804_ : new_n7080_) : ~new_n7079_);
  assign new_n7079_ = (new_n3318_ | new_n3313_) & (\i[1090]  | \i[1091]  | ~new_n3313_);
  assign new_n7080_ = ~\i[1067]  & (~\i[1066]  | (~\i[1065]  & ~\i[1064] ));
  assign new_n7081_ = ~new_n3998_ & (new_n6693_ | (new_n4445_ & (new_n4810_ ? \i[1411]  : new_n4939_)));
  assign new_n7082_ = new_n7083_ ? (~new_n7084_ ^ new_n7100_) : (new_n7084_ ^ new_n7100_);
  assign new_n7083_ = (new_n6710_ & new_n6721_) | (~new_n6695_ & (new_n6710_ | new_n6721_));
  assign new_n7084_ = new_n7085_ ? (new_n7093_ ^ new_n7099_) : (~new_n7093_ ^ new_n7099_);
  assign new_n7085_ = new_n6198_ ? (new_n6982_ ? new_n7092_ : new_n7086_) : new_n7088_;
  assign new_n7086_ = ~new_n7087_ & ((\i[1308]  & \i[1309]  & \i[1310] ) | \i[1311]  | ~new_n7002_);
  assign new_n7087_ = ~new_n3858_ & ~\i[1535]  & new_n7001_ & (~\i[1534]  | ~\i[1533] );
  assign new_n7088_ = new_n4884_ ? new_n7089_ : (new_n5843_ ? new_n7091_ : ~new_n7008_);
  assign new_n7089_ = new_n7006_ ? ((\i[1214]  | \i[1215]  | ~new_n3695_) & (~new_n7090_ | new_n3695_)) : ~new_n7005_;
  assign new_n7090_ = ~\i[1411]  & (~\i[1410]  | (~\i[1409]  & ~\i[1408] ));
  assign new_n7091_ = (new_n5762_ | ~new_n4781_ | ~new_n4782_) & (~\i[658]  | ~\i[659]  | (new_n4781_ & new_n4782_));
  assign new_n7092_ = (new_n6863_ | ~new_n6288_ | ~new_n6799_) & (~new_n3415_ | ~new_n4717_ | new_n6799_);
  assign new_n7093_ = (new_n7094_ | new_n3854_) & (new_n5828_ | new_n6655_ | ~new_n5197_ | ~new_n3789_ | ~new_n3854_);
  assign new_n7094_ = new_n6724_ ? new_n7097_ : ((new_n7095_ | ~new_n3771_) & (~new_n6688_ | ~new_n7098_ | new_n3771_));
  assign new_n7095_ = (~new_n4884_ & ~new_n7096_) | (~\i[1327]  & new_n7096_ & (~\i[1326]  | ~\i[1325] ));
  assign new_n7096_ = ~\i[2151]  & (~\i[2150]  | (~\i[2149]  & ~\i[2148] ));
  assign new_n7097_ = (~new_n5011_ | ~new_n5826_ | new_n3259_) & (new_n3229_ | new_n6731_ | ~new_n3259_);
  assign new_n7098_ = \i[963]  & (\i[961]  | \i[962]  | \i[960] );
  assign new_n7099_ = ~new_n4100_ & new_n3905_ & ((new_n6698_ & new_n6699_) | (~new_n4090_ & ~\i[1839]  & ~new_n6699_));
  assign new_n7100_ = (new_n6749_ & new_n6764_) | (new_n6737_ & (new_n6749_ | new_n6764_));
  assign new_n7101_ = new_n7102_ ? (~new_n7103_ ^ new_n7121_) : (new_n7103_ ^ new_n7121_);
  assign new_n7102_ = (~new_n6877_ & new_n6840_) | (new_n6802_ & (~new_n6877_ | new_n6840_));
  assign new_n7103_ = new_n7104_ ? (new_n7112_ ^ new_n7113_) : (~new_n7112_ ^ new_n7113_);
  assign new_n7104_ = new_n7105_ ? (new_n7107_ ^ new_n7111_) : (~new_n7107_ ^ new_n7111_);
  assign new_n7105_ = (new_n7106_ | new_n6932_) & (new_n4716_ | new_n6922_ | ~new_n6919_ | ~new_n6932_);
  assign new_n7106_ = (~new_n4217_ | ~new_n6924_ | ~new_n6808_) & (new_n5543_ | new_n6929_ | new_n6930_ | new_n6808_);
  assign new_n7107_ = (new_n7108_ | new_n4929_) & (new_n4878_ | ~new_n6354_ | ~new_n7110_ | ~new_n4929_);
  assign new_n7108_ = (new_n7109_ | ~new_n3447_) & (new_n3321_ | new_n3368_ | \i[974]  | \i[975]  | new_n3447_);
  assign new_n7109_ = ~new_n6773_ & (\i[1507]  | ~new_n3574_);
  assign new_n7110_ = \i[2743]  & ~\i[2187]  & \i[2742] ;
  assign new_n7111_ = new_n6743_ & new_n6748_ & new_n5576_ & ~new_n6741_ & ~new_n6742_;
  assign new_n7112_ = (~new_n6823_ & new_n6809_) | (~new_n6803_ & (~new_n6823_ | new_n6809_));
  assign new_n7113_ = new_n7114_ ? (new_n7116_ ^ new_n7117_) : (~new_n7116_ ^ new_n7117_);
  assign new_n7114_ = (new_n7115_ | ~new_n3376_) & (new_n5460_ | new_n6713_ | new_n6714_ | ~new_n6688_ | new_n3376_);
  assign new_n7115_ = (~new_n6720_ | ~new_n5651_) & (new_n3364_ | ~new_n3219_ | ~new_n5025_ | new_n5651_);
  assign new_n7116_ = (new_n6763_ | new_n6992_ | ~new_n6997_) & (new_n6997_ | (\i[419]  ? new_n6996_ : new_n6991_));
  assign new_n7117_ = (new_n7118_ | new_n4960_) & (new_n4818_ | ~new_n7120_ | ~new_n4960_);
  assign new_n7118_ = (~new_n6975_ | ~new_n7119_ | ~new_n6673_) & (~new_n5721_ | ~new_n6973_ | ~new_n6971_ | new_n6673_);
  assign new_n7119_ = new_n3790_ & new_n4695_;
  assign new_n7120_ = new_n5804_ & new_n5568_ & (\i[1323]  | (\i[1321]  & \i[1322] ));
  assign new_n7121_ = (~new_n6774_ & new_n6733_) | (~new_n6736_ & (~new_n6774_ | new_n6733_));
  assign new_n7122_ = new_n7123_ ? (~new_n7124_ ^ new_n7128_) : (new_n7124_ ^ new_n7128_);
  assign new_n7123_ = (~new_n6889_ & ~new_n6903_) | (~new_n6801_ & (~new_n6889_ | ~new_n6903_));
  assign new_n7124_ = new_n7125_ ? (new_n7126_ ^ new_n7127_) : (~new_n7126_ ^ new_n7127_);
  assign new_n7125_ = (~new_n6857_ & new_n6865_) | (~new_n6841_ & (~new_n6857_ | new_n6865_));
  assign new_n7126_ = ~new_n4437_ & new_n6785_ & \i[2855]  & (\i[2854]  | \i[2853]  | \i[2852] );
  assign new_n7127_ = new_n3726_ & ~new_n6980_ & ~new_n6198_ & ~new_n4816_ & ~new_n3996_;
  assign new_n7128_ = (~new_n6946_ & ~new_n6952_) | (new_n6935_ & (~new_n6946_ | ~new_n6952_));
  assign new_n7129_ = (~new_n6960_ & ~new_n6977_) | (~new_n6934_ & (~new_n6960_ | ~new_n6977_));
  assign \o[37]  = ~new_n7131_ ^ new_n7132_;
  assign new_n7131_ = (~new_n7036_ & new_n7035_) | (new_n7034_ & (~new_n7036_ | new_n7035_));
  assign new_n7132_ = new_n7133_ ^ new_n7134_;
  assign new_n7133_ = (~new_n7038_ & new_n7129_) | (new_n7037_ & (~new_n7038_ | new_n7129_));
  assign new_n7134_ = new_n7135_ ? (~new_n7136_ ^ new_n7163_) : (new_n7136_ ^ new_n7163_);
  assign new_n7135_ = (~new_n7040_ & ~new_n7122_) | (new_n7039_ & (~new_n7040_ | ~new_n7122_));
  assign new_n7136_ = new_n7137_ ? (new_n7138_ ^ new_n7159_) : (~new_n7138_ ^ new_n7159_);
  assign new_n7137_ = (~new_n7042_ & ~new_n7101_) | (new_n7041_ & (~new_n7042_ | ~new_n7101_));
  assign new_n7138_ = new_n7139_ ? (new_n7140_ ^ new_n7155_) : (~new_n7140_ ^ new_n7155_);
  assign new_n7139_ = (~new_n7044_ & ~new_n7082_) | (new_n7043_ & (~new_n7044_ | ~new_n7082_));
  assign new_n7140_ = new_n7141_ ? (new_n7144_ ^ new_n7145_) : (~new_n7144_ ^ new_n7145_);
  assign new_n7141_ = ~new_n7142_ ^ new_n7143_;
  assign new_n7142_ = (~new_n7052_ & ~new_n7060_) | (new_n7046_ & (~new_n7052_ | ~new_n7060_));
  assign new_n7143_ = (~new_n7093_ & new_n7099_) | (~new_n7085_ & (~new_n7093_ | new_n7099_));
  assign new_n7144_ = (~new_n7067_ & new_n7066_) | (~new_n7045_ & (~new_n7067_ | new_n7066_));
  assign new_n7145_ = new_n7146_ ^ new_n7147_;
  assign new_n7146_ = new_n7068_ & new_n7075_;
  assign new_n7147_ = new_n7148_ ? (new_n7153_ ^ new_n7154_) : (~new_n7153_ ^ new_n7154_);
  assign new_n7148_ = new_n4380_ ? new_n7149_ : new_n7151_;
  assign new_n7149_ = (new_n7150_ | new_n6669_) & (new_n6677_ | ~new_n6676_ | ~new_n4433_ | ~new_n6669_);
  assign new_n7150_ = (~new_n6670_ | ~new_n6672_ | new_n6673_) & (~new_n6673_ | (new_n3467_ ? ~new_n3889_ : ~new_n4206_));
  assign new_n7151_ = ~new_n7152_ & (new_n6684_ | ~new_n3494_ | ~new_n6680_ | ~new_n6679_);
  assign new_n7152_ = new_n6684_ & new_n3318_ & (new_n6682_ ? ~new_n5530_ : ~new_n7074_);
  assign new_n7153_ = \i[1943]  & \i[1942]  & new_n3624_ & new_n4520_ & new_n6654_;
  assign new_n7154_ = new_n7080_ & new_n3998_ & new_n5842_ & ~new_n5698_ & ~new_n3462_;
  assign new_n7155_ = new_n7156_ ? (new_n7157_ ^ new_n7158_) : (~new_n7157_ ^ new_n7158_);
  assign new_n7156_ = (~new_n7084_ & new_n7100_) | (new_n7083_ & (~new_n7084_ | new_n7100_));
  assign new_n7157_ = (~new_n7113_ & new_n7112_) | (~new_n7104_ & (~new_n7113_ | new_n7112_));
  assign new_n7158_ = (~new_n7117_ & new_n7116_) | (~new_n7114_ & (~new_n7117_ | new_n7116_));
  assign new_n7159_ = new_n7160_ ? (new_n7161_ ^ new_n7162_) : (~new_n7161_ ^ new_n7162_);
  assign new_n7160_ = (~new_n7103_ & new_n7121_) | (new_n7102_ & (~new_n7103_ | new_n7121_));
  assign new_n7161_ = (new_n7126_ & new_n7127_) | (new_n7125_ & (new_n7126_ | new_n7127_));
  assign new_n7162_ = (~new_n7107_ & new_n7111_) | (~new_n7105_ & (~new_n7107_ | new_n7111_));
  assign new_n7163_ = (~new_n7124_ & new_n7128_) | (new_n7123_ & (~new_n7124_ | new_n7128_));
  assign \o[38]  = ((new_n7165_ | new_n7166_) & (~new_n7167_ ^ ~new_n7168_)) | (~new_n7165_ & ~new_n7166_ & (~new_n7167_ ^ new_n7168_));
  assign new_n7165_ = ~new_n7132_ & new_n7131_;
  assign new_n7166_ = ~new_n7134_ & new_n7133_;
  assign new_n7167_ = (~new_n7136_ & new_n7163_) | (new_n7135_ & (~new_n7136_ | new_n7163_));
  assign new_n7168_ = new_n7169_ ? (~new_n7170_ ^ new_n7179_) : (new_n7170_ ^ new_n7179_);
  assign new_n7169_ = (~new_n7138_ & ~new_n7159_) | (new_n7137_ & (~new_n7138_ | ~new_n7159_));
  assign new_n7170_ = new_n7171_ ? (~new_n7172_ ^ new_n7178_) : (new_n7172_ ^ new_n7178_);
  assign new_n7171_ = (~new_n7140_ & ~new_n7155_) | (new_n7139_ & (~new_n7140_ | ~new_n7155_));
  assign new_n7172_ = new_n7173_ ? (~new_n7174_ ^ new_n7177_) : (new_n7174_ ^ new_n7177_);
  assign new_n7173_ = (~new_n7145_ & new_n7144_) | (~new_n7141_ & (~new_n7145_ | new_n7144_));
  assign new_n7174_ = new_n7175_ ^ new_n7176_;
  assign new_n7175_ = ~new_n7146_ & new_n7147_;
  assign new_n7176_ = (new_n7153_ & new_n7154_) | (~new_n7148_ & (new_n7153_ | new_n7154_));
  assign new_n7177_ = new_n7142_ & new_n7143_;
  assign new_n7178_ = (new_n7157_ & new_n7158_) | (new_n7156_ & (new_n7157_ | new_n7158_));
  assign new_n7179_ = (new_n7161_ & new_n7162_) | (new_n7160_ & (new_n7161_ | new_n7162_));
  assign \o[39]  = ~new_n7181_ ^ new_n7182_;
  assign new_n7181_ = (new_n7167_ | (~new_n7168_ & (new_n7166_ | new_n7165_))) & (new_n7166_ | new_n7165_ | ~new_n7168_);
  assign new_n7182_ = new_n7183_ ^ new_n7184_;
  assign new_n7183_ = (~new_n7170_ & new_n7179_) | (new_n7169_ & (~new_n7170_ | new_n7179_));
  assign new_n7184_ = ~new_n7185_ ^ new_n7186_;
  assign new_n7185_ = (~new_n7172_ & new_n7178_) | (new_n7171_ & (~new_n7172_ | new_n7178_));
  assign new_n7186_ = ~new_n7187_ ^ new_n7188_;
  assign new_n7187_ = (~new_n7174_ & new_n7177_) | (new_n7173_ & (~new_n7174_ | new_n7177_));
  assign new_n7188_ = ~new_n7175_ & ~new_n7176_;
  assign \o[40]  = ((new_n7190_ | new_n7191_) & (~new_n7192_ ^ new_n7193_)) | (~new_n7190_ & ~new_n7191_ & (~new_n7192_ ^ ~new_n7193_));
  assign new_n7190_ = ~new_n7182_ & new_n7181_;
  assign new_n7191_ = ~new_n7184_ & new_n7183_;
  assign new_n7192_ = new_n7185_ & new_n7186_;
  assign new_n7193_ = ~new_n7188_ & new_n7187_;
  assign \o[41]  = (new_n7193_ | new_n7190_ | new_n7191_) & (new_n7192_ | (new_n7193_ & (new_n7190_ | new_n7191_)));
  assign \o[42]  = new_n7196_ ? (new_n7506_ ^ new_n7518_) : (~new_n7506_ ^ new_n7518_);
  assign new_n7196_ = new_n7197_ ? (~new_n7447_ ^ new_n7490_) : (new_n7447_ ^ new_n7490_);
  assign new_n7197_ = new_n7198_ ? (~new_n7340_ ^ new_n7433_) : (new_n7340_ ^ new_n7433_);
  assign new_n7198_ = new_n7199_ ? (new_n7261_ ^ new_n7333_) : (~new_n7261_ ^ new_n7333_);
  assign new_n7199_ = new_n7200_ ? (~new_n7243_ ^ new_n7254_) : (new_n7243_ ^ new_n7254_);
  assign new_n7200_ = new_n7201_ ? (~new_n7217_ ^ new_n7228_) : (new_n7217_ ^ new_n7228_);
  assign new_n7201_ = (~new_n7215_ & ~new_n7202_ & new_n4074_) | (~new_n4074_ & (new_n7216_ ? new_n7207_ : new_n7210_));
  assign new_n7202_ = ~new_n7206_ & (new_n6726_ ? (new_n3375_ ? ~new_n7205_ : new_n5062_) : new_n7203_);
  assign new_n7203_ = (new_n7204_ | ~\i[2057]  | ~\i[2058]  | ~\i[2059] ) & (~\i[2051]  | ~new_n6442_ | (\i[2057]  & \i[2058]  & \i[2059] ));
  assign new_n7204_ = new_n4674_ & ~\i[2408]  & ~\i[2409] ;
  assign new_n7205_ = ~\i[2494]  & ~\i[2495]  & (~\i[2493]  | ~\i[2492] );
  assign new_n7206_ = \i[1091]  & (\i[1090]  | \i[1089] );
  assign new_n7207_ = (new_n7208_ | ~new_n3994_ | (\i[1836]  & \i[1837] )) & (~new_n6773_ | ~new_n4247_ | (new_n3994_ & (~\i[1836]  | ~\i[1837] )));
  assign new_n7208_ = new_n5034_ ? (\i[395]  | (\i[393]  & \i[394] )) : new_n7209_;
  assign new_n7209_ = ~\i[939]  & (~\i[937]  | ~\i[938]  | ~\i[936] );
  assign new_n7210_ = \i[1715]  ? ~new_n7211_ : (new_n7214_ ? new_n4433_ : new_n3795_);
  assign new_n7211_ = ~new_n7212_ & ~new_n7213_;
  assign new_n7212_ = \i[835]  & (\i[833]  | \i[834]  | \i[832] );
  assign new_n7213_ = \i[1171]  & (\i[1169]  | \i[1170]  | \i[1168] );
  assign new_n7214_ = \i[2099]  & (\i[2098]  | \i[2097] );
  assign new_n7215_ = new_n7206_ & ((~new_n6062_ & ~new_n6762_) | (~\i[2434]  & ~\i[2435]  & new_n6762_));
  assign new_n7216_ = ~\i[403]  & (~\i[402]  | (~\i[401]  & ~\i[400] ));
  assign new_n7217_ = \i[1839]  ? ((new_n7222_ | ~new_n7227_) & (new_n7224_ | new_n7226_ | new_n7227_)) : new_n7218_;
  assign new_n7218_ = new_n3253_ ? (new_n3340_ ? new_n7219_ : new_n7221_) : new_n7220_;
  assign new_n7219_ = (new_n6729_ | ~new_n4696_) & (~new_n3397_ | ~\i[1710]  | ~\i[1711]  | new_n4696_);
  assign new_n7220_ = (new_n3273_ | ~new_n6535_ | new_n3854_) & (~new_n3854_ | (new_n6956_ ? new_n5588_ : ~new_n4805_));
  assign new_n7221_ = (\i[1851]  & (\i[1849]  | \i[1850] )) ? ~new_n4238_ : new_n5031_;
  assign new_n7222_ = (~new_n7223_ | new_n4750_) & (new_n5717_ | ~new_n4938_ | ~new_n4750_);
  assign new_n7223_ = \i[2513]  & \i[2514]  & \i[2515]  & (~\i[1667]  | ~\i[1666]  | ~\i[1665] );
  assign new_n7224_ = ~new_n3988_ & new_n7225_ & \i[1427]  & (\i[1426]  | \i[1425]  | \i[1424] );
  assign new_n7225_ = ~\i[1307]  & (~\i[1305]  | ~\i[1306]  | ~\i[1304] );
  assign new_n7226_ = new_n6288_ & ~\i[395]  & ~\i[394]  & ~\i[393]  & ~new_n7225_ & ~\i[392] ;
  assign new_n7227_ = ~\i[2407]  & ~\i[2406]  & ~\i[2404]  & ~\i[2405] ;
  assign new_n7228_ = (new_n7233_ | new_n7241_ | ~new_n4018_) & (new_n4018_ | (new_n6313_ ? new_n7236_ : new_n7229_));
  assign new_n7229_ = (~new_n7230_ | ~new_n7231_) & (new_n7232_ | \i[485]  | \i[486]  | \i[487]  | new_n7231_);
  assign new_n7230_ = ~new_n5957_ & ~\i[2403]  & (~\i[2402]  | ~\i[2401] );
  assign new_n7231_ = ~\i[967]  & ~new_n4782_ & ~\i[966] ;
  assign new_n7232_ = \i[2111]  & (\i[2110]  | (\i[2109]  & \i[2108] ));
  assign new_n7233_ = new_n7234_ & ((~\i[523]  & (~\i[521]  | ~\i[522] )) ? new_n6361_ : new_n7235_);
  assign new_n7234_ = ~\i[1284]  & ~\i[1285]  & new_n4235_ & (\i[715]  | \i[714] );
  assign new_n7235_ = ~\i[2215]  & ~\i[2214]  & ~\i[2212]  & ~\i[2213] ;
  assign new_n7236_ = new_n7239_ ? new_n7237_ : (new_n3677_ ? new_n3585_ : ~new_n7240_);
  assign new_n7237_ = new_n6808_ ? (\i[1963]  | (\i[1961]  & \i[1962] )) : new_n7238_;
  assign new_n7238_ = \i[655]  & (\i[653]  | \i[654]  | \i[652] );
  assign new_n7239_ = \i[1295]  & (\i[1294]  | (\i[1293]  & \i[1292] ));
  assign new_n7240_ = ~\i[371]  & ~\i[370]  & ~\i[368]  & ~\i[369] ;
  assign new_n7241_ = ~\i[714]  & ~\i[715]  & (new_n7242_ ? ~\i[1191]  : (\i[607]  | \i[606] ));
  assign new_n7242_ = ~\i[1207]  & (~\i[1206]  | (~\i[1205]  & ~\i[1204] ));
  assign new_n7243_ = (new_n7244_ & ~new_n3340_) | (~new_n7249_ & new_n3340_ & (~new_n3763_ | new_n7251_));
  assign new_n7244_ = new_n4389_ ? new_n7245_ : (new_n5100_ ? new_n7248_ : ~new_n7247_);
  assign new_n7245_ = (~new_n5184_ & ~new_n7246_) | (\i[2519]  & new_n7246_ & (\i[2518]  | \i[2517] ));
  assign new_n7246_ = \i[2275]  & (\i[2274]  | (\i[2273]  & \i[2272] ));
  assign new_n7247_ = (\i[1605]  & \i[1606]  & \i[1607] ) ? (~\i[1642]  | ~\i[1643] ) : new_n5827_;
  assign new_n7248_ = \i[2431]  & \i[2430]  & ~new_n4877_ & new_n4153_;
  assign new_n7249_ = new_n7250_ & ((~\i[2077]  & new_n5078_) ? new_n6257_ : ~new_n3458_);
  assign new_n7250_ = ~new_n3763_ & \i[1731]  & (\i[1730]  | (\i[1728]  & \i[1729] ));
  assign new_n7251_ = new_n7252_ ? new_n7253_ : ((~new_n6132_ & new_n5802_) | (~\i[638]  & ~\i[639]  & ~new_n5802_));
  assign new_n7252_ = \i[1967]  & \i[1965]  & \i[1966] ;
  assign new_n7253_ = ~\i[1767]  & ~\i[1766]  & ~\i[1835]  & (~\i[1834]  | ~\i[1833]  | ~\i[1832] );
  assign new_n7254_ = new_n3309_ ? new_n7255_ : ((~new_n7260_ & new_n4111_) | (~new_n7259_ & ~new_n7257_ & ~new_n4111_));
  assign new_n7255_ = (~new_n4848_ | ~new_n6415_ | new_n6098_) & (~new_n6098_ | (new_n4291_ ? ~new_n4946_ : new_n7256_));
  assign new_n7256_ = new_n3736_ & (~\i[2303]  | (~\i[2300]  & ~\i[2301]  & ~\i[2302] ));
  assign new_n7257_ = new_n7258_ & \i[2278]  & \i[2279]  & (\i[1715]  | (\i[1714]  & new_n3526_));
  assign new_n7258_ = \i[1275]  & (\i[1274]  | \i[1273] );
  assign new_n7259_ = ~new_n7258_ & (new_n4216_ ? new_n4662_ : new_n5670_);
  assign new_n7260_ = \i[1203]  & (\i[1202]  | (\i[1201]  & \i[1200] ));
  assign new_n7261_ = new_n7262_ ? (~new_n7299_ ^ new_n7326_) : (new_n7299_ ^ new_n7326_);
  assign new_n7262_ = new_n7263_ ? (~new_n7276_ ^ new_n7288_) : (new_n7276_ ^ new_n7288_);
  assign new_n7263_ = new_n7275_ ? (new_n4206_ ? new_n7270_ : ~new_n7273_) : new_n7264_;
  assign new_n7264_ = new_n5456_ ? (new_n7267_ | (~new_n7268_ & ~new_n7269_ & new_n3722_)) : new_n7265_;
  assign new_n7265_ = (new_n7266_ | ~new_n5237_) & (~new_n5429_ | ~new_n6110_ | new_n5237_);
  assign new_n7266_ = (\i[487]  | \i[486]  | ~new_n5743_) & (~\i[967]  | new_n5743_ | (~\i[966]  & ~\i[965] ));
  assign new_n7267_ = ~new_n3722_ & ~new_n5588_ & (~new_n4337_ | (\i[2064]  & \i[2065] ));
  assign new_n7268_ = ~\i[1819]  & (~\i[1817]  | ~\i[1818]  | ~\i[1816] );
  assign new_n7269_ = ~\i[2183]  & (~\i[2182]  | ~\i[2181] );
  assign new_n7270_ = new_n5038_ ? new_n7271_ : (new_n3998_ ? new_n7272_ : ~new_n4732_);
  assign new_n7271_ = ~new_n5616_ & (\i[2317]  | \i[2318]  | \i[2319] );
  assign new_n7272_ = ~\i[1099]  & ~\i[1097]  & ~\i[1098] ;
  assign new_n7273_ = (new_n7274_ | (new_n6005_ ? ~new_n5048_ : ~new_n4190_)) & (new_n6729_ | \i[1179]  | ~new_n7274_);
  assign new_n7274_ = ~\i[2303]  & ~\i[2301]  & ~\i[2302] ;
  assign new_n7275_ = \i[2179]  & (\i[2178]  | \i[2177] );
  assign new_n7276_ = (new_n7285_ | ~new_n7286_) & (new_n7277_ | ~new_n7287_);
  assign new_n7277_ = (~\i[2498]  & ~\i[2499]  & new_n7281_ & ~\i[2497] ) | (~new_n7284_ & ~new_n7278_ & (\i[2497]  | \i[2498]  | \i[2499] ));
  assign new_n7278_ = ~new_n7280_ & (new_n5925_ ? new_n5698_ : ~new_n7279_);
  assign new_n7279_ = ~\i[750]  & ~\i[751]  & (~\i[749]  | ~\i[748] );
  assign new_n7280_ = ~\i[1827]  & ~\i[1825]  & ~\i[1826] ;
  assign new_n7281_ = (~new_n7204_ | (new_n7282_ ? ~new_n7283_ : ~new_n5102_)) & (~new_n4774_ | ~new_n3289_ | new_n7204_);
  assign new_n7282_ = ~\i[1551]  & (~\i[1550]  | (~\i[1549]  & ~\i[1548] ));
  assign new_n7283_ = ~\i[2299]  & (~\i[2297]  | ~\i[2298]  | ~\i[2296] );
  assign new_n7284_ = ~new_n6403_ & ~\i[666]  & ~\i[667]  & new_n7280_ & (~\i[665]  | ~\i[664] );
  assign new_n7285_ = \i[875]  & \i[874]  & \i[873]  & \i[872]  & ~new_n4244_ & new_n4149_;
  assign new_n7286_ = ~new_n7287_ & (~\i[652]  | ~\i[653]  | ~\i[654]  | ~\i[655] );
  assign new_n7287_ = ~\i[2743]  & ~\i[2742]  & ~\i[2740]  & ~\i[2741] ;
  assign new_n7288_ = ~new_n7289_ & (~new_n4084_ | (~new_n7291_ & (new_n7296_ | new_n7298_ | new_n3274_)));
  assign new_n7289_ = ~new_n4084_ & ~new_n7290_ & (~\i[659]  | (~\i[658]  & (~\i[657]  | ~\i[656] )));
  assign new_n7290_ = \i[635]  & \i[634]  & \i[633]  & \i[632]  & new_n3455_ & new_n3512_;
  assign new_n7291_ = new_n3274_ & ((new_n7293_ & new_n6519_ & ~new_n7292_) | (new_n7292_ & (~new_n7295_ | ~new_n7294_)));
  assign new_n7292_ = ~\i[1611]  & (~\i[1610]  | ~\i[1609] );
  assign new_n7293_ = ~\i[1939]  & (~\i[1938]  | (~\i[1937]  & ~\i[1936] ));
  assign new_n7294_ = ~\i[1554]  & ~\i[1555]  & (~\i[1553]  | ~\i[1552] );
  assign new_n7295_ = ~\i[1414]  & ~\i[1415]  & (~\i[1413]  | ~\i[1412] );
  assign new_n7296_ = new_n5223_ & (new_n6658_ ? ~new_n7297_ : (\i[1527]  | (\i[1525]  & \i[1526] )));
  assign new_n7297_ = \i[1066]  & \i[1067]  & (\i[1065]  | \i[1064] );
  assign new_n7298_ = ~new_n5223_ & ~new_n3996_ & ~\i[759]  & (~\i[758]  | (~\i[756]  & ~\i[757] ));
  assign new_n7299_ = ~new_n7300_ ^ new_n7314_;
  assign new_n7300_ = new_n5507_ ? ((~new_n7311_ & new_n7313_) | (~new_n7308_ & ~new_n7310_ & ~new_n7313_)) : new_n7301_;
  assign new_n7301_ = ~new_n7302_ & (new_n7303_ | (~new_n7306_ & (new_n6790_ | (~new_n7307_ & new_n3278_))));
  assign new_n7302_ = new_n7303_ & (new_n3394_ ? new_n7304_ : (new_n4704_ ? new_n3735_ : new_n4809_));
  assign new_n7303_ = new_n3416_ & (~\i[969]  | ~\i[968] );
  assign new_n7304_ = (new_n7305_ | ~new_n3393_) & (\i[1550]  | \i[1551]  | new_n3393_);
  assign new_n7305_ = ~\i[1727]  & (~\i[1726]  | (~\i[1725]  & ~\i[1724] ));
  assign new_n7306_ = new_n6790_ & ~\i[663]  & ~\i[662]  & ~\i[660]  & ~\i[661] ;
  assign new_n7307_ = ~\i[1195]  & ~\i[1193]  & ~\i[1194] ;
  assign new_n7308_ = new_n7309_ & (new_n3399_ ? ~new_n6292_ : new_n6655_);
  assign new_n7309_ = \i[1943]  & (\i[1942]  | \i[1941] );
  assign new_n7310_ = ~new_n7309_ & (~new_n3761_ | (~\i[415]  & (~\i[414]  | (~\i[412]  & ~\i[413] ))));
  assign new_n7311_ = (new_n5440_ | ~new_n7312_ | (\i[2282]  & \i[2283] )) & (~\i[2282]  | ~\i[2283]  | new_n3322_ | new_n4291_);
  assign new_n7312_ = \i[1550]  & \i[1551]  & (\i[1549]  | \i[1548] );
  assign new_n7313_ = ~\i[539]  & (~\i[537]  | ~\i[538]  | ~\i[536] );
  assign new_n7314_ = new_n4809_ ? new_n7315_ : ((~new_n7321_ & new_n3415_) | (~new_n7324_ & ~new_n7325_ & ~new_n3415_));
  assign new_n7315_ = ~new_n7316_ & (new_n7319_ | new_n7320_ | ~new_n5733_);
  assign new_n7316_ = new_n7319_ & (~new_n6155_ | new_n7318_ | ~new_n6655_) & (~new_n7317_ | ~new_n6948_ | new_n6655_);
  assign new_n7317_ = \i[2379]  & (\i[2378]  | (\i[2377]  & \i[2376] ));
  assign new_n7318_ = ~\i[267]  & ~\i[266]  & ~\i[264]  & ~\i[265] ;
  assign new_n7319_ = ~\i[279]  & ~\i[278]  & ~\i[276]  & ~\i[277] ;
  assign new_n7320_ = ~\i[959]  & ~\i[957]  & ~\i[958] ;
  assign new_n7321_ = new_n3369_ ? new_n4222_ : (new_n7322_ ? new_n7323_ : new_n5827_);
  assign new_n7322_ = \i[1267]  & (\i[1266]  | \i[1265] );
  assign new_n7323_ = ~\i[1630]  & ~\i[1631]  & (~\i[1629]  | ~\i[1628] );
  assign new_n7324_ = new_n4018_ & (\i[394]  | \i[395]  | (~new_n6976_ & (~\i[392]  | ~\i[393] )));
  assign new_n7325_ = new_n3587_ & ~new_n3400_ & ~new_n4018_;
  assign new_n7326_ = (~\i[1078]  & ~\i[1079] ) ? new_n7327_ : (new_n4195_ ? new_n7331_ : ~new_n4166_);
  assign new_n7327_ = ~new_n7328_ & (~new_n7330_ | (~\i[2295]  & (~\i[2294]  | ~\i[2293] )));
  assign new_n7328_ = ~\i[714]  & ~\i[715]  & ((~new_n7329_ & ~\i[871] ) | (new_n4265_ & new_n4304_ & \i[871] ));
  assign new_n7329_ = (new_n4046_ & new_n4674_) | (new_n4199_ & ~new_n4674_ & (~\i[2061]  | ~\i[2060] ));
  assign new_n7330_ = ~new_n4167_ & ~\i[730]  & ~\i[731]  & (\i[715]  | \i[714] );
  assign new_n7331_ = (~new_n6119_ | ~new_n6155_ | ~new_n3494_) & (new_n7332_ | ~\i[1171]  | new_n3494_);
  assign new_n7332_ = ~\i[1170]  & (~\i[1169]  | ~\i[1168] );
  assign new_n7333_ = new_n3512_ & (new_n7334_ | (~new_n5387_ & ~new_n7339_ & (\i[1611]  | new_n7337_)));
  assign new_n7334_ = new_n5387_ & (new_n7336_ ? (~new_n5062_ | (~\i[1302]  & ~\i[1303] )) : new_n7335_);
  assign new_n7335_ = (new_n5397_ & new_n5431_) | (\i[503]  & ~new_n5431_ & (\i[502]  | \i[501] ));
  assign new_n7336_ = ~\i[1627]  & (~\i[1625]  | ~\i[1626]  | ~\i[1624] );
  assign new_n7337_ = (new_n4057_ & ~new_n7338_) | (~\i[723]  & new_n7338_ & (~\i[722]  | ~\i[721] ));
  assign new_n7338_ = \i[951]  & (\i[949]  | \i[950]  | \i[948] );
  assign new_n7339_ = \i[1611]  & ~new_n6884_ & ~\i[1839] ;
  assign new_n7340_ = new_n7341_ ? (~new_n7407_ ^ new_n7419_) : (new_n7407_ ^ new_n7419_);
  assign new_n7341_ = new_n7342_ ? (~new_n7375_ ^ new_n7397_) : (new_n7375_ ^ new_n7397_);
  assign new_n7342_ = new_n7343_ ? (~new_n7355_ ^ new_n7366_) : (new_n7355_ ^ new_n7366_);
  assign new_n7343_ = new_n7354_ ? ((~new_n6235_ & new_n7352_) | (~new_n3683_ & ~new_n7349_)) : new_n7344_;
  assign new_n7344_ = (new_n7345_ & ~\i[1660]  & ~\i[1661]  & ~\i[1662]  & ~\i[1663] ) | (~new_n5152_ & (\i[1660]  | \i[1661]  | \i[1662]  | \i[1663] ));
  assign new_n7345_ = (\i[2627]  & (\i[2625]  | \i[2626] )) ? new_n7346_ : new_n7347_;
  assign new_n7346_ = (new_n5544_ | ~new_n3998_) & (~\i[514]  | ~\i[515]  | new_n3998_);
  assign new_n7347_ = new_n3479_ ? new_n7348_ : (\i[1403]  | (\i[1401]  & \i[1402] ));
  assign new_n7348_ = ~\i[2402]  & ~\i[2403]  & (~\i[2401]  | ~\i[2400] );
  assign new_n7349_ = (new_n3450_ | new_n6813_ | \i[1063]  | (\i[1061]  & \i[1062] )) & (new_n7350_ | (~\i[1063]  & (~\i[1061]  | ~\i[1062] )));
  assign new_n7350_ = new_n7214_ ? ~new_n7351_ : (\i[2063]  | (\i[2061]  & \i[2062] ));
  assign new_n7351_ = ~\i[2307]  & (~\i[2306]  | ~\i[2305] );
  assign new_n7352_ = new_n3683_ & new_n3799_ & ~\i[1773]  & ~new_n7353_ & ~\i[1772] ;
  assign new_n7353_ = \i[1610]  & \i[1611] ;
  assign new_n7354_ = \i[1839]  & (\i[1838]  | (\i[1837]  & \i[1836] ));
  assign new_n7355_ = (new_n7365_ | ~new_n3259_ | new_n6098_) & (~new_n6098_ | (~new_n7361_ & (new_n7275_ | new_n7356_)));
  assign new_n7356_ = new_n7358_ ? (new_n7359_ ? new_n7360_ : ~new_n4681_) : new_n7357_;
  assign new_n7357_ = (\i[1083]  | \i[1082]  | new_n3340_) & (\i[2521]  | \i[2522]  | \i[2523]  | ~new_n3340_);
  assign new_n7358_ = ~\i[2167]  & (~\i[2166]  | (~\i[2165]  & ~\i[2164] ));
  assign new_n7359_ = ~\i[2159]  & (~\i[2158]  | ~\i[2157] );
  assign new_n7360_ = ~\i[2175]  & (~\i[2173]  | ~\i[2174]  | ~\i[2172] );
  assign new_n7361_ = new_n7275_ & (new_n7364_ ? new_n7362_ : new_n7363_);
  assign new_n7362_ = new_n7283_ ? (\i[2287]  | (\i[2285]  & \i[2286] )) : ~\i[1067] ;
  assign new_n7363_ = (~new_n4060_ & new_n3399_) | (\i[1763]  & ~new_n3399_ & (\i[1762]  | \i[1761] ));
  assign new_n7364_ = \i[2207]  & (\i[2206]  | \i[2205] );
  assign new_n7365_ = ~new_n6348_ & (~\i[2169]  | ~\i[2170]  | ~\i[2171] );
  assign new_n7366_ = new_n3781_ ? new_n7373_ : (new_n4947_ ? new_n7368_ : new_n7367_);
  assign new_n7367_ = (new_n7227_ | ~new_n6713_ | ~new_n3502_) & (new_n5842_ | ~new_n6784_ | new_n3502_);
  assign new_n7368_ = (~\i[2303]  & (~\i[2301]  | ~\i[2302] )) ? new_n7371_ : new_n7369_;
  assign new_n7369_ = new_n4654_ ? ~new_n7370_ : (~\i[847]  & (~\i[844]  | ~\i[845]  | ~\i[846] ));
  assign new_n7370_ = ~\i[2639]  & ~\i[2637]  & ~\i[2638] ;
  assign new_n7371_ = (~\i[606]  & ~\i[607] ) ? ~new_n6672_ : ~new_n7372_;
  assign new_n7372_ = \i[1383]  & (\i[1382]  | (\i[1381]  & \i[1380] ));
  assign new_n7373_ = (new_n4147_ & new_n6198_ & \i[635] ) | (~\i[635]  & (~new_n7374_ | ~new_n6929_));
  assign new_n7374_ = \i[1938]  & \i[1939]  & (\i[1937]  | \i[1936] );
  assign new_n7375_ = new_n7376_ ? (new_n7382_ ^ new_n7391_) : (~new_n7382_ ^ new_n7391_);
  assign new_n7376_ = (new_n7377_ & ~\i[2604]  & ~\i[2605]  & ~\i[2606]  & ~\i[2607] ) | (~new_n7381_ & (\i[2604]  | \i[2605]  | \i[2606]  | \i[2607] ));
  assign new_n7377_ = (new_n7378_ | \i[2742]  | \i[2743] ) & (~\i[2395]  | ~\i[2393]  | ~\i[2394]  | (~\i[2742]  & ~\i[2743] ));
  assign new_n7378_ = (new_n7379_ | \i[834]  | \i[835]  | new_n7380_) & (~new_n7380_ | (~new_n4947_ & new_n3997_));
  assign new_n7379_ = ~\i[1287]  & (~\i[1286]  | (~\i[1285]  & ~\i[1284] ));
  assign new_n7380_ = ~\i[1071]  & ~\i[1069]  & ~\i[1070] ;
  assign new_n7381_ = \i[1979]  & \i[1978]  & \i[1976]  & \i[1977] ;
  assign new_n7382_ = new_n5007_ ? ((~new_n7388_ & ~new_n7272_ & new_n3375_) | (~new_n7390_ & ~new_n3375_)) : new_n7383_;
  assign new_n7383_ = new_n7386_ ? new_n7384_ : ((new_n7387_ | ~new_n4141_) & (~new_n7380_ | ~new_n4018_ | new_n4141_));
  assign new_n7384_ = new_n6081_ ? ~new_n7385_ : (~\i[1091]  & (~\i[1088]  | ~\i[1089]  | ~\i[1090] ));
  assign new_n7385_ = ~\i[1415]  & (~\i[1413]  | ~\i[1414]  | ~\i[1412] );
  assign new_n7386_ = ~\i[1403]  & ~\i[1401]  & ~\i[1402] ;
  assign new_n7387_ = \i[1633]  & \i[1634]  & \i[1635]  & (\i[1411]  | \i[1410] );
  assign new_n7388_ = (\i[2427]  & (\i[2425]  | \i[2426] )) ? new_n6683_ : new_n7389_;
  assign new_n7389_ = \i[1263]  & (\i[1262]  | (\i[1261]  & \i[1260] ));
  assign new_n7390_ = (new_n3458_ | new_n3502_) & (new_n3304_ | new_n6672_ | ~new_n3502_);
  assign new_n7391_ = ~new_n7395_ & ~new_n7392_ & (~\i[2495]  | (~\i[2494]  & (~\i[2493]  | ~\i[2492] )));
  assign new_n7392_ = ~new_n7394_ & (new_n7393_ | (~new_n6385_ & (new_n4121_ ? ~new_n5695_ : ~\i[427] )));
  assign new_n7393_ = new_n6385_ & (new_n5733_ | new_n4809_) & (\i[2752]  | \i[2753]  | ~new_n3849_ | ~new_n4809_);
  assign new_n7394_ = \i[646]  & \i[647]  & (\i[645]  | \i[644] );
  assign new_n7395_ = new_n7394_ & (new_n5611_ ? (new_n5738_ ? new_n4192_ : new_n7396_) : new_n3308_);
  assign new_n7396_ = ~\i[2511]  & (~\i[2509]  | ~\i[2510]  | ~\i[2508] );
  assign new_n7397_ = new_n7275_ ? new_n7398_ : (new_n3399_ ? new_n7406_ : new_n7403_);
  assign new_n7398_ = new_n4035_ ? new_n3659_ : (new_n4701_ ? new_n7399_ : new_n7400_);
  assign new_n7399_ = (~\i[1723]  & (~\i[1721]  | ~\i[1722] )) ? ~new_n4098_ : ~new_n5651_;
  assign new_n7400_ = (~new_n7401_ | ~new_n7402_) & (\i[1066]  | \i[1067]  | new_n7402_ | (\i[1065]  & \i[1064] ));
  assign new_n7401_ = ~\i[2383]  & ~\i[2382]  & ~\i[2380]  & ~\i[2381] ;
  assign new_n7402_ = ~\i[943]  & (~\i[942]  | (~\i[941]  & ~\i[940] ));
  assign new_n7403_ = new_n4134_ ? (new_n4286_ ? ~new_n7405_ : new_n6324_) : new_n7404_;
  assign new_n7404_ = (~\i[1279]  | ~\i[1278]  | new_n7225_) & (\i[494]  | \i[495]  | \i[493]  | ~new_n7225_);
  assign new_n7405_ = ~\i[1171]  & (~\i[1170]  | ~\i[1169] );
  assign new_n7406_ = ~\i[1998]  & ~\i[1999]  & new_n4469_ & (~\i[1041]  | ~\i[1040]  | ~new_n6525_);
  assign new_n7407_ = (new_n7416_ | new_n7417_ | new_n4368_) & (new_n7408_ | new_n7414_ | ~new_n4368_);
  assign new_n7408_ = ~\i[2051]  & ~new_n7409_ & ~new_n6442_;
  assign new_n7409_ = ~new_n7410_ & ((\i[2157]  & \i[2158]  & \i[2159] ) | new_n7413_ | ~new_n7412_);
  assign new_n7410_ = (\i[1947]  | (\i[1945]  & \i[1946] )) & (new_n4119_ ? ~new_n5483_ : new_n7411_);
  assign new_n7411_ = ~\i[2291]  & (~\i[2289]  | ~\i[2290]  | ~\i[2288] );
  assign new_n7412_ = ~new_n3431_ & ~\i[1947]  & (~\i[1946]  | ~\i[1945] );
  assign new_n7413_ = \i[2167]  & \i[2164]  & ~\i[2166]  & \i[2165] ;
  assign new_n7414_ = \i[2535]  & \i[2534]  & \i[2533]  & \i[2532]  & ~new_n3573_ & new_n7415_;
  assign new_n7415_ = (\i[2051]  | new_n6442_) & (~new_n5740_ | (~\i[2217]  & ~\i[2216] ));
  assign new_n7416_ = ~new_n3619_ & ((new_n3254_ & new_n6951_ & ~new_n3394_) | (~new_n5404_ & new_n3586_ & new_n3394_));
  assign new_n7417_ = new_n3619_ & ((new_n5087_ & \i[1407]  & new_n7418_) | (new_n3504_ & new_n4018_ & ~new_n7418_));
  assign new_n7418_ = \i[1738]  & \i[1739]  & (\i[1737]  | \i[1736] );
  assign new_n7419_ = (~new_n7420_ & ~new_n7424_ & new_n7432_) | (~new_n7432_ & (new_n7428_ | (~new_n7431_ & new_n5563_)));
  assign new_n7420_ = new_n7422_ & (~new_n4678_ | new_n7421_);
  assign new_n7421_ = \i[967]  & (\i[966]  | new_n4782_);
  assign new_n7422_ = ~new_n7209_ & (new_n4678_ | new_n7423_ | ~new_n4393_);
  assign new_n7423_ = \i[1311]  & (\i[1310]  | (\i[1309]  & \i[1308] ));
  assign new_n7424_ = new_n7425_ & (\i[385]  | \i[386]  | \i[387]  | ~new_n7426_ | ~new_n6813_);
  assign new_n7425_ = new_n7209_ & (new_n7426_ | new_n7427_ | (~\i[819]  & (~\i[816]  | ~new_n6779_)));
  assign new_n7426_ = ~\i[1203]  & (~\i[1201]  | ~\i[1202]  | ~\i[1200] );
  assign new_n7427_ = \i[1651]  & (\i[1650]  | (\i[1649]  & \i[1648] ));
  assign new_n7428_ = ~new_n5563_ & ((~new_n4041_ & ~new_n4851_ & new_n7429_) | (new_n7430_ & ~new_n7429_));
  assign new_n7429_ = new_n6085_ & (~\i[845]  | ~\i[844] );
  assign new_n7430_ = ~new_n4942_ & \i[1499]  & (~\i[827]  | (~\i[825]  & ~\i[826] ));
  assign new_n7431_ = (new_n6117_ | new_n5422_ | ~new_n6862_) & (~new_n3223_ | new_n6862_ | (~\i[391]  & ~\i[390] ));
  assign new_n7432_ = ~\i[719]  & ~\i[717]  & ~\i[718] ;
  assign new_n7433_ = new_n4409_ ? new_n7434_ : (~new_n7440_ & (new_n7445_ | ~new_n3637_ | ~new_n7446_));
  assign new_n7434_ = new_n3342_ ? (\i[1295]  ? new_n7438_ : new_n7439_) : new_n7435_;
  assign new_n7435_ = (~new_n7436_ | ~new_n3299_ | new_n5472_) & (~new_n5472_ | (new_n6167_ ? ~new_n7437_ : new_n3439_));
  assign new_n7436_ = ~\i[2411]  & (~\i[2410]  | (~\i[2409]  & ~\i[2408] ));
  assign new_n7437_ = \i[1615]  & (\i[1614]  | (\i[1613]  & \i[1612] ));
  assign new_n7438_ = (~new_n3462_ | new_n3585_) & (~\i[2517]  | ~\i[2518]  | ~\i[2519]  | ~new_n3585_);
  assign new_n7439_ = (~new_n3889_ | \i[607] ) & (\i[1394]  | \i[1395]  | ~\i[607]  | (\i[1393]  & \i[1392] ));
  assign new_n7440_ = new_n7443_ & (~new_n7441_ | (~\i[2531]  & (~\i[2530]  | (~\i[2528]  & ~\i[2529] ))));
  assign new_n7441_ = ~new_n7442_ & (~\i[519]  | (~\i[518]  & (~\i[517]  | ~\i[516] )));
  assign new_n7442_ = ~\i[2639]  & ~\i[2638]  & ~\i[2636]  & ~\i[2637] ;
  assign new_n7443_ = ~new_n3637_ & (\i[2059]  | ~new_n7444_ | ~\i[1535]  | ~new_n7442_);
  assign new_n7444_ = (~\i[2058]  | (~\i[2056]  & ~\i[2057] )) & (\i[1534]  | (\i[1533]  & \i[1532] ));
  assign new_n7445_ = new_n3562_ ? ~new_n5497_ : (~\i[663]  & (~\i[660]  | ~\i[661]  | ~\i[662] ));
  assign new_n7446_ = ~\i[1327]  & (~\i[1325]  | ~\i[1326]  | ~\i[1324] );
  assign new_n7447_ = new_n7448_ ? (new_n7474_ ^ new_n7485_) : (~new_n7474_ ^ new_n7485_);
  assign new_n7448_ = new_n7449_ ? (~new_n7457_ ^ new_n7465_) : (new_n7457_ ^ new_n7465_);
  assign new_n7449_ = (~\i[1551]  & (~\i[1548]  | ~\i[1549]  | ~\i[1550] )) ? new_n7450_ : ~new_n7456_;
  assign new_n7450_ = new_n6670_ ? (~new_n7455_ & (~new_n6726_ | ~new_n5845_ | ~new_n6683_)) : new_n7451_;
  assign new_n7451_ = ~new_n7453_ & (~new_n7452_ | (\i[1616]  & \i[1617]  & \i[1618]  & \i[1619] ));
  assign new_n7452_ = ~new_n6288_ & (\i[1408]  | \i[1409]  | \i[1410]  | \i[1411] );
  assign new_n7453_ = new_n6288_ & new_n7454_ & \i[951]  & (\i[950]  | \i[949] );
  assign new_n7454_ = \i[2283]  & \i[2282]  & \i[2280]  & \i[2281] ;
  assign new_n7455_ = ~new_n6726_ & ~new_n3585_ & \i[2395]  & (\i[2394]  | \i[2393]  | \i[2392] );
  assign new_n7456_ = new_n4288_ & ((~\i[1721]  & ~\i[1720] ) | ~\i[1723]  | ~\i[1722] );
  assign new_n7457_ = new_n7464_ ? ((new_n7462_ | new_n7353_) & (new_n4355_ | ~new_n6826_ | ~new_n7353_)) : new_n7458_;
  assign new_n7458_ = (new_n3273_ | (new_n4393_ ? ~new_n7460_ : ~new_n7459_)) & (~new_n7461_ | ~new_n4779_ | ~new_n3273_);
  assign new_n7459_ = ~new_n6459_ & (\i[1715]  | (\i[1712]  & \i[1713]  & \i[1714] ));
  assign new_n7460_ = (~new_n4060_ | ~new_n4235_) & (\i[734]  | \i[735]  | new_n4235_);
  assign new_n7461_ = (\i[1063]  | (\i[1062]  & \i[1061] )) & (~new_n3670_ | (\i[1940]  & \i[1941] ));
  assign new_n7462_ = ~new_n7463_ & ((\i[2298]  & \i[2299] ) | new_n6138_ | ~new_n5845_);
  assign new_n7463_ = ~new_n6168_ & \i[1615]  & \i[2298]  & \i[2299]  & (\i[1614]  | \i[1613] );
  assign new_n7464_ = \i[1838]  & \i[1839] ;
  assign new_n7465_ = (~new_n7472_ & ~new_n7466_ & ~new_n3726_) | (new_n3726_ & (new_n7469_ | (~new_n7467_ & new_n5437_)));
  assign new_n7466_ = ~new_n6655_ & (new_n5763_ ? (new_n4395_ | (\i[1618]  & \i[1619] )) : ~new_n6122_);
  assign new_n7467_ = ~new_n7468_ & (\i[1607]  | ~new_n6413_ | ~new_n4147_);
  assign new_n7468_ = ~new_n6413_ & (\i[1603]  ? (~\i[523]  | (~\i[521]  & ~\i[522] )) : new_n4875_);
  assign new_n7469_ = new_n7470_ & (new_n6325_ | (~new_n7394_ & ~\i[519] ) | (~new_n7471_ & \i[519] ));
  assign new_n7470_ = ~new_n5437_ & (\i[2551]  | ~new_n6325_ | (\i[2550]  & (\i[2548]  | \i[2549] )));
  assign new_n7471_ = \i[2179]  & (\i[2178]  | (\i[2177]  & \i[2176] ));
  assign new_n7472_ = new_n6655_ & (~new_n3532_ | \i[1667]  | ~new_n3638_) & (new_n5115_ | new_n7473_ | new_n3638_);
  assign new_n7473_ = ~\i[2438]  & ~\i[2439] ;
  assign new_n7474_ = new_n5048_ ? (new_n4060_ ? new_n7479_ : new_n7475_) : new_n7484_;
  assign new_n7475_ = new_n6413_ ? ~new_n7478_ : new_n7476_;
  assign new_n7476_ = (new_n7477_ | ~new_n3377_) & (\i[737]  | \i[738]  | \i[739]  | new_n3377_);
  assign new_n7477_ = \i[2634]  & \i[2635]  & (\i[2633]  | \i[2632] );
  assign new_n7478_ = (~\i[1169]  | ~\i[1170]  | ~\i[1171]  | \i[951] ) & (~\i[951]  | (\i[635]  & \i[634] ));
  assign new_n7479_ = new_n7483_ ? new_n7480_ : new_n7482_;
  assign new_n7480_ = (~new_n3779_ | new_n7481_) & (~\i[511]  | ~new_n7481_ | (~\i[510]  & (~\i[508]  | ~\i[509] )));
  assign new_n7481_ = ~\i[531]  & (~\i[530]  | ~\i[529] );
  assign new_n7482_ = new_n3340_ ? (~\i[2067]  & (~\i[2064]  | ~\i[2065]  | ~\i[2066] )) : \i[611] ;
  assign new_n7483_ = ~\i[2422]  & ~\i[2423]  & (~\i[2421]  | ~\i[2420] );
  assign new_n7484_ = (~new_n5567_ | ~new_n4149_ | ~new_n3717_) & (~new_n3462_ | ~\i[2310]  | ~\i[2311]  | new_n3717_);
  assign new_n7485_ = new_n3512_ & ((~new_n7489_ & ~new_n7240_) | (~new_n7488_ & new_n7240_ & (new_n6243_ | new_n7486_)));
  assign new_n7486_ = new_n4521_ ? ~new_n5541_ : new_n7487_;
  assign new_n7487_ = ~\i[1259]  & ~\i[1258]  & ~\i[1256]  & ~\i[1257] ;
  assign new_n7488_ = new_n7294_ & new_n6243_ & (~\i[2295]  | (~\i[2292]  & ~\i[2293]  & ~\i[2294] ));
  assign new_n7489_ = (\i[501]  | \i[502]  | \i[503]  | ~new_n3627_) & (new_n4939_ | new_n3627_);
  assign new_n7490_ = new_n7505_ ? new_n7491_ : (~new_n7497_ & (new_n7502_ | ~new_n7501_ | ~new_n7504_));
  assign new_n7491_ = new_n3760_ ? (new_n7495_ | (~new_n7496_ & new_n4779_ & new_n3313_)) : new_n7492_;
  assign new_n7492_ = new_n5125_ ? new_n7493_ : ((~\i[1434]  & ~\i[1435] ) ? ~new_n5056_ : ~new_n7380_);
  assign new_n7493_ = new_n7494_ ? new_n5030_ : (\i[723]  | (\i[721]  & \i[722] ));
  assign new_n7494_ = ~\i[2415]  & (~\i[2413]  | ~\i[2414]  | ~\i[2412] );
  assign new_n7495_ = ~new_n3313_ & new_n7028_ & (~\i[2527]  | ~\i[2526] );
  assign new_n7496_ = ~\i[2403]  & ~\i[2401]  & ~\i[2402] ;
  assign new_n7497_ = ~new_n7501_ & ((~new_n3585_ & ~new_n7498_ & \i[1303] ) | (~\i[1303]  & (~new_n7500_ | new_n7499_)));
  assign new_n7498_ = \i[1390]  & \i[1391]  & (\i[1389]  | \i[1388] );
  assign new_n7499_ = ~\i[423]  & (~\i[422]  | (~\i[421]  & ~\i[420] ));
  assign new_n7500_ = \i[2494]  & \i[2495]  & (\i[2493]  | \i[2492] );
  assign new_n7501_ = ~\i[531]  & ~\i[530]  & ~\i[528]  & ~\i[529] ;
  assign new_n7502_ = new_n7503_ & \i[1663]  & (\i[1662]  | \i[1661]  | \i[1660] );
  assign new_n7503_ = ~\i[655]  & (~\i[654]  | ~\i[653] );
  assign new_n7504_ = ~\i[471]  & (~\i[470]  | (~\i[469]  & ~\i[468] ));
  assign new_n7505_ = ~\i[967]  & ~\i[965]  & ~\i[966] ;
  assign new_n7506_ = new_n7517_ ? new_n7512_ : ((~\i[2502]  & ~\i[2503] ) ? new_n7507_ : new_n7510_);
  assign new_n7507_ = (new_n7508_ & ~new_n5635_) | (~new_n7509_ & new_n5635_ & (new_n3997_ | (~\i[1946]  & ~\i[1947] )));
  assign new_n7508_ = (~new_n5495_ & ~\i[536]  & ~\i[537]  & ~\i[538]  & ~\i[539] ) | (~new_n5703_ & (\i[536]  | \i[537]  | \i[538]  | \i[539] ));
  assign new_n7509_ = ~\i[1658]  & ~\i[1659]  & ~\i[1946]  & ~\i[1947]  & (~\i[1657]  | ~\i[1656] );
  assign new_n7510_ = (~new_n6204_ | ~\i[2499]  | ~new_n5049_) & (new_n7511_ | new_n5049_ | (~new_n6673_ & ~new_n5856_));
  assign new_n7511_ = new_n6673_ & ((\i[525]  & \i[524] ) | \i[527]  | \i[526] );
  assign new_n7512_ = (new_n4046_ | new_n7513_ | new_n7516_) & (~new_n7516_ | (new_n3289_ ? new_n7515_ : new_n7514_));
  assign new_n7513_ = (~\i[534]  & ~\i[535] ) ? (~\i[390]  | ~\i[391] ) : new_n3690_;
  assign new_n7514_ = new_n6778_ ? (~\i[535]  | (~\i[533]  & ~\i[534] )) : new_n3659_;
  assign new_n7515_ = (\i[1946]  & \i[1947] ) ? new_n4390_ : ~new_n6718_;
  assign new_n7516_ = \i[2283]  & (\i[2282]  | (\i[2281]  & \i[2280] ));
  assign new_n7517_ = ~\i[2175]  & (~\i[2174]  | ~\i[2173] );
  assign new_n7518_ = (new_n3619_ & (new_n3716_ ? new_n7523_ : new_n7525_)) | (~new_n7521_ & ~new_n7519_ & ~new_n3619_);
  assign new_n7519_ = ~new_n3400_ & new_n6676_ & (new_n7520_ ? new_n4018_ : ~new_n6655_);
  assign new_n7520_ = ~\i[427]  & (~\i[426]  | ~\i[425] );
  assign new_n7521_ = new_n3400_ & ((new_n7522_ & ~new_n6975_) | (~new_n4391_ & ~new_n4809_ & new_n6975_));
  assign new_n7522_ = ~new_n7294_ & (~\i[1201]  | ~\i[1202]  | ~\i[1203] );
  assign new_n7523_ = (new_n3779_ & (~new_n7353_ | ~new_n5066_)) | (~new_n6132_ & new_n7524_ & ~new_n3779_);
  assign new_n7524_ = ~\i[539]  & (~\i[538]  | (~\i[537]  & ~\i[536] ));
  assign new_n7525_ = (new_n7527_ | new_n7528_ | new_n7526_) & (~new_n3618_ | ~new_n5526_ | ~new_n7526_);
  assign new_n7526_ = \i[1951]  & \i[1949]  & \i[1950] ;
  assign new_n7527_ = \i[1551]  & (\i[1549]  | \i[1550]  | \i[1548] );
  assign new_n7528_ = ~\i[430]  & ~\i[431] ;
  assign \o[43]  = new_n7530_ ^ new_n7624_;
  assign new_n7530_ = new_n7531_ ? (~new_n7622_ ^ new_n7623_) : (new_n7622_ ^ new_n7623_);
  assign new_n7531_ = new_n7532_ ? (~new_n7611_ ^ new_n7612_) : (new_n7611_ ^ new_n7612_);
  assign new_n7532_ = new_n7533_ ? (~new_n7588_ ^ new_n7589_) : (new_n7588_ ^ new_n7589_);
  assign new_n7533_ = new_n7534_ ? (~new_n7571_ ^ new_n7587_) : (new_n7571_ ^ new_n7587_);
  assign new_n7534_ = new_n7535_ ? (new_n7556_ ^ new_n7557_) : (~new_n7556_ ^ new_n7557_);
  assign new_n7535_ = new_n7536_ ? (new_n7545_ ^ new_n7553_) : (~new_n7545_ ^ new_n7553_);
  assign new_n7536_ = (new_n7537_ & new_n5507_) | (~new_n7542_ & ~new_n5507_ & (~new_n7543_ | (~new_n3278_ & ~new_n7307_)));
  assign new_n7537_ = (new_n7538_ | ~new_n7313_) & (new_n7308_ | new_n7313_ | (~new_n7309_ & (new_n3761_ | new_n7541_)));
  assign new_n7538_ = (new_n7539_ & (~\i[2282]  | ~\i[2283] )) | (\i[2282]  & \i[2283]  & (new_n3322_ ? new_n7540_ : new_n4291_));
  assign new_n7539_ = (~new_n6240_ | ~new_n5440_) & (~\i[1550]  | ~\i[1551]  | new_n5440_ | (~\i[1549]  & ~\i[1548] ));
  assign new_n7540_ = ~\i[1439]  & ~\i[1437]  & ~\i[1438] ;
  assign new_n7541_ = ~\i[2319]  & ~\i[2318]  & ~\i[2316]  & ~\i[2317] ;
  assign new_n7542_ = new_n7303_ & (~new_n7305_ | ~new_n3393_ | ~new_n3394_) & (~new_n3735_ | ~new_n4704_ | new_n3394_);
  assign new_n7543_ = ~new_n6790_ & ~new_n7303_ & ~new_n7544_;
  assign new_n7544_ = new_n7307_ & (\i[656]  | \i[657]  | \i[658]  | \i[659] );
  assign new_n7545_ = (~new_n7549_ & ~new_n7546_ & ~new_n7517_) | (new_n7517_ & (new_n7516_ ? new_n7552_ : new_n7550_));
  assign new_n7546_ = ~\i[2502]  & ~\i[2503]  & (new_n5635_ ? ~new_n7509_ : (new_n7548_ | new_n7547_));
  assign new_n7547_ = new_n5703_ & (\i[536]  | \i[537]  | \i[538]  | \i[539] );
  assign new_n7548_ = ~\i[539]  & ~\i[538]  & ~\i[537]  & ~new_n5495_ & ~\i[536] ;
  assign new_n7549_ = (\i[2502]  | \i[2503] ) & ((new_n7511_ & ~new_n5049_) | (~\i[2499]  & new_n6204_ & new_n5049_));
  assign new_n7550_ = new_n4046_ ? (new_n4805_ ? new_n7269_ : ~new_n4398_) : ~new_n7551_;
  assign new_n7551_ = new_n3690_ & (\i[535]  | \i[534] );
  assign new_n7552_ = (~new_n4390_ | ~\i[1946]  | ~\i[1947]  | ~new_n3289_) & (~new_n3659_ | new_n6778_ | new_n3289_);
  assign new_n7553_ = (new_n7282_ | ~new_n7554_) & (~new_n7286_ | ~new_n4149_ | ~new_n4244_ | ~new_n7555_);
  assign new_n7554_ = new_n7287_ & new_n5102_ & new_n7204_ & ~\i[2499]  & ~\i[2497]  & ~\i[2498] ;
  assign new_n7555_ = ~\i[2199]  & ~\i[2197]  & ~\i[2198] ;
  assign new_n7556_ = ~new_n7314_ & new_n7300_;
  assign new_n7557_ = ~new_n7558_ ^ new_n7566_;
  assign new_n7558_ = new_n3619_ ? new_n7559_ : ((new_n7564_ | ~new_n3400_) & (~new_n7563_ | new_n7562_));
  assign new_n7559_ = new_n3716_ ? ((new_n7524_ | new_n3779_) & (\i[987]  | ~new_n7560_ | ~new_n3779_)) : new_n7561_;
  assign new_n7560_ = ~new_n5066_ & (~\i[984]  | ~\i[985]  | ~\i[986] );
  assign new_n7561_ = (new_n5526_ | ~new_n5007_ | ~new_n7526_) & (new_n7526_ | (new_n7527_ ? ~new_n3523_ : new_n7528_));
  assign new_n7562_ = ~new_n6676_ & (new_n6240_ ? ~new_n4742_ : (~\i[399]  | (~\i[397]  & ~\i[398] )));
  assign new_n7563_ = ~new_n3400_ & (~new_n6676_ | (~new_n7520_ & new_n6655_));
  assign new_n7564_ = (~new_n6684_ | ~new_n7294_ | new_n6975_) & (~new_n6975_ | (new_n4391_ ? ~new_n7565_ : ~new_n4809_));
  assign new_n7565_ = ~\i[1075]  & (~\i[1074]  | ~\i[1073] );
  assign new_n7566_ = ~new_n7567_ & (~new_n7570_ | (new_n3369_ & (new_n4222_ | new_n3467_)));
  assign new_n7567_ = new_n4809_ & (new_n7319_ ? ~new_n7568_ : (new_n7320_ ? new_n4946_ : ~new_n5733_));
  assign new_n7568_ = new_n6655_ ? (new_n7318_ ? new_n6307_ : ~new_n6155_) : new_n7569_;
  assign new_n7569_ = new_n6948_ ? new_n7317_ : ~new_n3998_;
  assign new_n7570_ = ~new_n4809_ & new_n3415_ & (new_n3369_ | (~new_n7323_ & new_n7322_));
  assign new_n7571_ = new_n7572_ ? (new_n7573_ ^ new_n7586_) : (~new_n7573_ ^ new_n7586_);
  assign new_n7572_ = (~new_n7217_ & ~new_n7228_) | (~new_n7201_ & (~new_n7217_ | ~new_n7228_));
  assign new_n7573_ = new_n7574_ ? (new_n7581_ ^ new_n7584_) : (~new_n7581_ ^ new_n7584_);
  assign new_n7574_ = new_n7505_ ? new_n7575_ : ((new_n7580_ | new_n7501_) & (new_n7579_ | ~new_n7504_ | ~new_n7501_));
  assign new_n7575_ = ~new_n7576_ & ((~new_n5030_ & new_n5125_ & new_n7494_) | new_n3760_ | new_n7578_);
  assign new_n7576_ = new_n7577_ & (~new_n3313_ | ((~new_n7496_ | ~new_n4779_) & (~\i[986]  | ~\i[987]  | new_n4779_)));
  assign new_n7577_ = new_n3760_ & (new_n7028_ | new_n3313_ | (\i[483]  & (\i[481]  | \i[482] )));
  assign new_n7578_ = new_n5056_ & ~\i[1435]  & ~new_n5125_ & ~\i[1434] ;
  assign new_n7579_ = ~new_n7502_ & (new_n7503_ | ~new_n6155_);
  assign new_n7580_ = (~new_n7498_ | new_n3585_ | ~\i[1303] ) & (\i[1303]  | (new_n7500_ ? new_n7499_ : ~new_n4119_));
  assign new_n7581_ = (new_n6413_ | ~new_n7583_ | ~new_n7477_ | ~new_n5048_) & (~new_n3717_ | new_n7582_ | new_n5048_);
  assign new_n7582_ = (~new_n4219_ | ~new_n5567_ | ~new_n4149_) & (~new_n3879_ | ~new_n4716_ | new_n4149_);
  assign new_n7583_ = ~new_n4060_ & new_n3377_;
  assign new_n7584_ = new_n4084_ & (new_n7585_ | (~new_n7294_ & new_n3274_ & new_n7292_ & new_n4028_));
  assign new_n7585_ = new_n3996_ & ~new_n7240_ & ~new_n3274_ & ~new_n5223_;
  assign new_n7586_ = (new_n7276_ & new_n7288_) | (~new_n7263_ & (new_n7276_ | new_n7288_));
  assign new_n7587_ = (~new_n7299_ & ~new_n7326_) | (~new_n7262_ & (~new_n7299_ | ~new_n7326_));
  assign new_n7588_ = (~new_n7261_ & new_n7333_) | (~new_n7199_ & (~new_n7261_ | new_n7333_));
  assign new_n7589_ = new_n7590_ ? (new_n7591_ ^ new_n7592_) : (~new_n7591_ ^ new_n7592_);
  assign new_n7590_ = (~new_n7243_ & ~new_n7254_) | (~new_n7200_ & (~new_n7243_ | ~new_n7254_));
  assign new_n7591_ = (~new_n7375_ & ~new_n7397_) | (~new_n7342_ & (~new_n7375_ | ~new_n7397_));
  assign new_n7592_ = new_n7593_ ? (new_n7603_ ^ new_n7610_) : (~new_n7603_ ^ new_n7610_);
  assign new_n7593_ = new_n7594_ ? (new_n7599_ ^ new_n7601_) : (~new_n7599_ ^ new_n7601_);
  assign new_n7594_ = new_n7275_ ? ((~new_n5038_ & ~new_n7598_ & new_n4206_) | (~new_n7273_ & ~new_n4206_)) : new_n7595_;
  assign new_n7595_ = ~new_n7596_ & (new_n5456_ | (new_n7266_ & new_n5237_) | (~\i[851]  & new_n7597_ & ~new_n5237_));
  assign new_n7596_ = ~new_n7267_ & new_n5456_ & (~new_n3722_ | (~\i[1423]  & new_n7268_) | (new_n7269_ & ~new_n7268_));
  assign new_n7597_ = ~new_n5429_ & (~\i[848]  | ~\i[849]  | ~\i[850] );
  assign new_n7598_ = new_n3998_ ? ~new_n7272_ : new_n4732_;
  assign new_n7599_ = \i[1839]  & ~new_n7600_ & new_n7227_;
  assign new_n7600_ = (~new_n5717_ | ~new_n4938_ | ~new_n4750_) & (~\i[1665]  | ~\i[1666]  | ~\i[1667]  | new_n4750_);
  assign new_n7601_ = ~new_n7602_ & (new_n4409_ | new_n7446_ | ~new_n5022_ | ~new_n3637_);
  assign new_n7602_ = new_n4409_ & new_n3299_ & ~new_n7436_ & ~new_n3342_ & ~new_n5472_;
  assign new_n7603_ = new_n7604_ ? (new_n7608_ ^ new_n7609_) : (~new_n7608_ ^ new_n7609_);
  assign new_n7604_ = new_n4018_ ? new_n7606_ : (new_n6313_ ? new_n7605_ : ~new_n7229_);
  assign new_n7605_ = new_n7239_ ? ~new_n7237_ : (new_n3677_ ? ~new_n3585_ : new_n7240_);
  assign new_n7606_ = ~new_n7607_ & (\i[523]  | ~new_n6361_ | ~new_n7234_ | (\i[522]  & \i[521] ));
  assign new_n7607_ = ~\i[714]  & ~\i[715]  & (new_n7242_ ? ~\i[1191]  : (\i[607]  | \i[606] ));
  assign new_n7608_ = new_n3512_ & new_n4939_ & ~new_n3627_ & ~new_n7240_;
  assign new_n7609_ = new_n3619_ & new_n3504_ & new_n4018_ & ~new_n4368_ & ~new_n7418_;
  assign new_n7610_ = (~new_n7382_ & new_n7391_) | (~new_n7376_ & (~new_n7382_ | new_n7391_));
  assign new_n7611_ = (~new_n7340_ & ~new_n7433_) | (~new_n7198_ & (~new_n7340_ | ~new_n7433_));
  assign new_n7612_ = new_n7613_ ? (new_n7614_ ^ new_n7621_) : (~new_n7614_ ^ new_n7621_);
  assign new_n7613_ = (~new_n7407_ & ~new_n7419_) | (~new_n7341_ & (~new_n7407_ | ~new_n7419_));
  assign new_n7614_ = new_n7615_ ? (~new_n7616_ ^ new_n7619_) : (new_n7616_ ^ new_n7619_);
  assign new_n7615_ = (~new_n7355_ & ~new_n7366_) | (~new_n7343_ & (~new_n7355_ | ~new_n7366_));
  assign new_n7616_ = (new_n4074_ | (new_n7216_ ? ~new_n7207_ : new_n7618_)) & (new_n7215_ | new_n7617_ | ~new_n4074_);
  assign new_n7617_ = ~new_n7206_ & (new_n6726_ ? (new_n3375_ ? ~new_n7205_ : new_n5062_) : new_n7203_);
  assign new_n7618_ = (new_n7211_ | ~\i[1715] ) & (new_n7214_ | ~new_n3795_ | \i[1715] );
  assign new_n7619_ = (~new_n7422_ & ~new_n7424_ & new_n7432_) | (~new_n7432_ & (new_n7620_ | new_n7428_));
  assign new_n7620_ = ~new_n6862_ & new_n3223_ & new_n5563_ & (\i[391]  | \i[390] );
  assign new_n7621_ = (~new_n7457_ & ~new_n7465_) | (~new_n7449_ & (~new_n7457_ | ~new_n7465_));
  assign new_n7622_ = (~new_n7447_ & ~new_n7490_) | (~new_n7197_ & (~new_n7447_ | ~new_n7490_));
  assign new_n7623_ = (~new_n7474_ & new_n7485_) | (~new_n7448_ & (~new_n7474_ | new_n7485_));
  assign new_n7624_ = (~new_n7506_ & ~new_n7518_) | (~new_n7196_ & (~new_n7506_ | ~new_n7518_));
  assign \o[44]  = ~new_n7626_ ^ new_n7627_;
  assign new_n7626_ = new_n7530_ & new_n7624_;
  assign new_n7627_ = new_n7628_ ^ new_n7629_;
  assign new_n7628_ = (new_n7622_ & new_n7623_) | (new_n7531_ & (new_n7622_ | new_n7623_));
  assign new_n7629_ = new_n7630_ ? (~new_n7631_ ^ new_n7660_) : (new_n7631_ ^ new_n7660_);
  assign new_n7630_ = (new_n7611_ & new_n7612_) | (new_n7532_ & (new_n7611_ | new_n7612_));
  assign new_n7631_ = new_n7632_ ? (new_n7633_ ^ new_n7656_) : (~new_n7633_ ^ new_n7656_);
  assign new_n7632_ = (new_n7588_ & new_n7589_) | (new_n7533_ & (new_n7588_ | new_n7589_));
  assign new_n7633_ = new_n7634_ ? (new_n7635_ ^ new_n7652_) : (~new_n7635_ ^ new_n7652_);
  assign new_n7634_ = (new_n7571_ & new_n7587_) | (new_n7534_ & (new_n7571_ | new_n7587_));
  assign new_n7635_ = new_n7636_ ? (new_n7637_ ^ new_n7640_) : (~new_n7637_ ^ new_n7640_);
  assign new_n7636_ = (~new_n7556_ & new_n7557_) | (new_n7535_ & (~new_n7556_ | new_n7557_));
  assign new_n7637_ = ~new_n7638_ ^ new_n7639_;
  assign new_n7638_ = (~new_n7545_ & ~new_n7553_) | (~new_n7536_ & (~new_n7545_ | ~new_n7553_));
  assign new_n7639_ = (~new_n7581_ & new_n7584_) | (~new_n7574_ & (~new_n7581_ | new_n7584_));
  assign new_n7640_ = new_n7641_ ? (~new_n7642_ ^ new_n7649_) : (new_n7642_ ^ new_n7649_);
  assign new_n7641_ = new_n7558_ & new_n7566_;
  assign new_n7642_ = ~new_n7643_ ^ new_n7647_;
  assign new_n7643_ = new_n4809_ ? ((new_n7646_ | ~new_n7319_) & (~new_n4946_ | ~new_n7320_ | new_n7319_)) : new_n7644_;
  assign new_n7644_ = (~new_n6976_ | ~new_n7645_) & (~new_n3369_ | ~new_n3415_ | (new_n4222_ & ~new_n3611_));
  assign new_n7645_ = ~new_n3415_ & ~\i[394]  & ~\i[395]  & new_n4018_ & (~\i[393]  | ~\i[392] );
  assign new_n7646_ = (new_n7318_ | ~new_n6155_ | ~new_n6655_) & (new_n7317_ | ~new_n6948_ | new_n6655_);
  assign new_n7647_ = ~new_n3619_ & (new_n7648_ | (new_n7563_ & (new_n6676_ | (~new_n4742_ & new_n6240_))));
  assign new_n7648_ = \i[1203]  & \i[1202]  & \i[1201]  & new_n3400_ & ~new_n6975_ & ~new_n7294_;
  assign new_n7649_ = (new_n7650_ & (new_n7504_ | new_n7505_ | ~new_n7501_)) | (~new_n7504_ & ~new_n7505_ & new_n7501_ & ~new_n7650_);
  assign new_n7650_ = ~new_n7651_ & (new_n7303_ | new_n5507_ | new_n7306_ | (~new_n6790_ & ~new_n7544_));
  assign new_n7651_ = new_n5507_ & new_n7309_ & new_n6655_ & ~new_n3399_ & ~new_n7313_;
  assign new_n7652_ = new_n7653_ ? (new_n7654_ ^ new_n7655_) : (~new_n7654_ ^ new_n7655_);
  assign new_n7653_ = (~new_n7573_ & new_n7586_) | (new_n7572_ & (~new_n7573_ | new_n7586_));
  assign new_n7654_ = (new_n7603_ & new_n7610_) | (new_n7593_ & (new_n7603_ | new_n7610_));
  assign new_n7655_ = (~new_n7601_ & new_n7599_) | (new_n7594_ & (~new_n7601_ | new_n7599_));
  assign new_n7656_ = new_n7657_ ? (~new_n7658_ ^ new_n7659_) : (new_n7658_ ^ new_n7659_);
  assign new_n7657_ = (~new_n7592_ & new_n7591_) | (new_n7590_ & (~new_n7592_ | new_n7591_));
  assign new_n7658_ = (~new_n7616_ & new_n7619_) | (new_n7615_ & (~new_n7616_ | new_n7619_));
  assign new_n7659_ = (~new_n7608_ & ~new_n7609_) | (new_n7604_ & (~new_n7608_ | ~new_n7609_));
  assign new_n7660_ = (~new_n7614_ & new_n7621_) | (new_n7613_ & (~new_n7614_ | new_n7621_));
  assign \o[45]  = ((new_n7662_ | new_n7663_) & (~new_n7664_ ^ new_n7665_)) | (~new_n7662_ & ~new_n7663_ & (~new_n7664_ ^ ~new_n7665_));
  assign new_n7662_ = ~new_n7627_ & new_n7626_;
  assign new_n7663_ = ~new_n7629_ & new_n7628_;
  assign new_n7664_ = (~new_n7631_ & new_n7660_) | (new_n7630_ & (~new_n7631_ | new_n7660_));
  assign new_n7665_ = new_n7666_ ? (new_n7667_ ^ new_n7677_) : (~new_n7667_ ^ new_n7677_);
  assign new_n7666_ = (~new_n7633_ & ~new_n7656_) | (new_n7632_ & (~new_n7633_ | ~new_n7656_));
  assign new_n7667_ = new_n7668_ ? (~new_n7669_ ^ new_n7676_) : (new_n7669_ ^ new_n7676_);
  assign new_n7668_ = (~new_n7635_ & ~new_n7652_) | (new_n7634_ & (~new_n7635_ | ~new_n7652_));
  assign new_n7669_ = new_n7670_ ? (~new_n7671_ ^ new_n7675_) : (new_n7671_ ^ new_n7675_);
  assign new_n7670_ = (~new_n7637_ & ~new_n7640_) | (new_n7636_ & (~new_n7637_ | ~new_n7640_));
  assign new_n7671_ = new_n7672_ ? (~new_n7673_ ^ new_n7674_) : (new_n7673_ ^ new_n7674_);
  assign new_n7672_ = (~new_n7642_ & ~new_n7649_) | (~new_n7641_ & (~new_n7642_ | ~new_n7649_));
  assign new_n7673_ = ~new_n7647_ & new_n7643_;
  assign new_n7674_ = new_n7501_ & ~new_n7505_ & ~new_n7650_ & ~new_n7504_;
  assign new_n7675_ = new_n7638_ & new_n7639_;
  assign new_n7676_ = (new_n7654_ & new_n7655_) | (new_n7653_ & (new_n7654_ | new_n7655_));
  assign new_n7677_ = (~new_n7659_ & new_n7658_) | (new_n7657_ & (~new_n7659_ | new_n7658_));
  assign \o[46]  = ~new_n7679_ ^ new_n7680_;
  assign new_n7679_ = (new_n7665_ | new_n7662_ | new_n7663_) & (new_n7664_ | (new_n7665_ & (new_n7662_ | new_n7663_)));
  assign new_n7680_ = new_n7681_ ^ new_n7682_;
  assign new_n7681_ = (~new_n7667_ & new_n7677_) | (new_n7666_ & (~new_n7667_ | new_n7677_));
  assign new_n7682_ = new_n7683_ ^ new_n7684_;
  assign new_n7683_ = (~new_n7669_ & new_n7676_) | (new_n7668_ & (~new_n7669_ | new_n7676_));
  assign new_n7684_ = ~new_n7685_ ^ new_n7686_;
  assign new_n7685_ = (~new_n7671_ & new_n7675_) | (new_n7670_ & (~new_n7671_ | new_n7675_));
  assign new_n7686_ = (~new_n7673_ & new_n7674_) | (new_n7672_ & (~new_n7673_ | new_n7674_));
  assign \o[47]  = ((new_n7688_ | new_n7689_) & (~new_n7690_ ^ new_n7691_)) | (~new_n7688_ & ~new_n7689_ & (~new_n7690_ ^ ~new_n7691_));
  assign new_n7688_ = ~new_n7680_ & new_n7679_;
  assign new_n7689_ = ~new_n7682_ & new_n7681_;
  assign new_n7690_ = ~new_n7684_ & new_n7683_;
  assign new_n7691_ = new_n7685_ & new_n7686_;
  assign \o[48]  = (new_n7691_ | new_n7688_ | new_n7689_) & (new_n7690_ | (new_n7691_ & (new_n7688_ | new_n7689_)));
  assign \o[49]  = new_n7694_ ^ new_n8000_;
  assign new_n7694_ = new_n7695_ ? (~new_n7787_ ^ new_n7990_) : (new_n7787_ ^ new_n7990_);
  assign new_n7695_ = new_n7696_ ? (~new_n7763_ ^ new_n7776_) : (new_n7763_ ^ new_n7776_);
  assign new_n7696_ = new_n7697_ ? (new_n7738_ ^ new_n7747_) : (~new_n7738_ ^ new_n7747_);
  assign new_n7697_ = new_n7698_ ? (~new_n7723_ ^ new_n7735_) : (new_n7723_ ^ new_n7735_);
  assign new_n7698_ = new_n7699_ ? (new_n7706_ ^ new_n7715_) : (~new_n7706_ ^ new_n7715_);
  assign new_n7699_ = (~\i[2170]  & ~\i[2171] ) ? (~new_n7704_ & ~new_n4304_) : new_n7700_;
  assign new_n7700_ = new_n7703_ ? ((new_n7701_ & ~new_n4231_) | (new_n6155_ & new_n7426_ & new_n4231_)) : ~new_n7702_;
  assign new_n7701_ = ~new_n4190_ & ~new_n5820_;
  assign new_n7702_ = (\i[1878]  | \i[1879]  | new_n5396_) & (~new_n3477_ | (~\i[2161]  & ~\i[2160] ));
  assign new_n7703_ = ~\i[1939]  & (~\i[1937]  | ~\i[1938]  | ~\i[1936] );
  assign new_n7704_ = (new_n7705_ | new_n5721_) & (~new_n3731_ | ~new_n3843_ | ~new_n5721_);
  assign new_n7705_ = (\i[2291]  & (\i[2289]  | \i[2290] )) ? ~new_n6154_ : new_n3437_;
  assign new_n7706_ = new_n7713_ ? (new_n7712_ ? ~new_n7707_ : ~new_n7710_) : ~new_n7714_;
  assign new_n7707_ = (new_n7708_ | new_n3905_) & (new_n7709_ | ~new_n4236_ | ~new_n3905_);
  assign new_n7708_ = ~new_n5636_ & ~\i[1535]  & (~\i[1534]  | ~\i[1533]  | ~\i[1532] );
  assign new_n7709_ = new_n4120_ & (~\i[825]  | ~\i[824] );
  assign new_n7710_ = new_n7471_ ? (~new_n5262_ & (\i[1057]  | \i[1058]  | \i[1059] )) : new_n7711_;
  assign new_n7711_ = ~\i[2322]  & ~\i[2323]  & (~\i[2321]  | ~\i[2320] );
  assign new_n7712_ = ~\i[815]  & (~\i[813]  | ~\i[814]  | ~\i[812] );
  assign new_n7713_ = ~\i[2547]  & (~\i[2545]  | ~\i[2546]  | ~\i[2544] );
  assign new_n7714_ = \i[1259]  & (\i[1258]  | \i[1257] );
  assign new_n7715_ = (new_n7716_ | ~new_n7712_) & (new_n7721_ | ~new_n4100_ | ~new_n7722_ | new_n7712_);
  assign new_n7716_ = (~new_n4679_ | ~new_n7720_ | ~new_n7555_) & (new_n7717_ | new_n7719_ | new_n7555_);
  assign new_n7717_ = new_n4247_ & (new_n7718_ | (\i[1260]  & \i[1261]  & \i[1262]  & \i[1263] ));
  assign new_n7718_ = \i[1874]  & \i[1875]  & (\i[1873]  | \i[1872] );
  assign new_n7719_ = ~new_n4247_ & ((\i[2085]  & \i[2086] ) | \i[2087]  | (\i[1147]  & \i[1146] ));
  assign new_n7720_ = \i[818]  & \i[819]  & (\i[817]  | \i[816] );
  assign new_n7721_ = \i[2087]  & (\i[2086]  | (\i[2085]  & \i[2084] ));
  assign new_n7722_ = ~\i[1759]  & ~\i[1757]  & ~\i[1758] ;
  assign new_n7723_ = new_n5422_ ? (new_n7732_ | (~new_n7724_ & ~\i[1841]  & new_n4109_)) : new_n7727_;
  assign new_n7724_ = new_n6848_ ? (~new_n7726_ & (~new_n7258_ | ~\i[1166]  | ~\i[1167] )) : new_n7725_;
  assign new_n7725_ = ~new_n3548_ & ~\i[1142]  & ~\i[1143]  & (~\i[1141]  | ~\i[1140] );
  assign new_n7726_ = ~\i[831]  & ~\i[830]  & (~\i[1166]  | ~\i[1167] ) & (~\i[828]  | ~\i[829] );
  assign new_n7727_ = (new_n7728_ | new_n7731_) & (new_n6719_ | ~new_n7731_ | (new_n4701_ ? new_n4453_ : \i[1887] ));
  assign new_n7728_ = (new_n4681_ | new_n7730_ | ~\i[1055] ) & (\i[1055]  | (new_n7729_ ? new_n6214_ : ~new_n5082_));
  assign new_n7729_ = \i[1747]  & \i[1745]  & \i[1746] ;
  assign new_n7730_ = \i[815]  & (\i[814]  | (\i[813]  & \i[812] ));
  assign new_n7731_ = ~\i[1395]  & ~\i[1393]  & ~\i[1394] ;
  assign new_n7732_ = (new_n7734_ | ~\i[2279] ) & (\i[1841]  | ~new_n4109_) & (new_n6525_ | ~new_n7733_ | \i[2279] );
  assign new_n7733_ = ~\i[1031]  & ~\i[1030]  & ~\i[1028]  & ~\i[1029] ;
  assign new_n7734_ = ~\i[1619]  & (~\i[1618]  | ~\i[1617] );
  assign new_n7735_ = ~new_n7737_ & ~\i[2315]  & ((new_n7736_ & ~\i[927] ) | (~new_n4100_ & new_n6452_ & \i[927] ));
  assign new_n7736_ = ~new_n4105_ & \i[1623]  & (\i[1622]  | \i[1621]  | \i[1620] );
  assign new_n7737_ = \i[2655]  & (\i[2653]  | \i[2654]  | \i[2652] );
  assign new_n7738_ = ~new_n7739_ & (~new_n3652_ | (new_n7745_ & (new_n5957_ | ~new_n4659_ | ~new_n6061_)));
  assign new_n7739_ = ~new_n3652_ & ~new_n7740_ & (~new_n7742_ | (new_n7743_ & (~new_n7744_ | new_n6110_)));
  assign new_n7740_ = new_n7714_ & ((new_n7741_ & ~new_n5316_) | (new_n7360_ & new_n5316_ & (\i[2631]  | \i[2630] )));
  assign new_n7741_ = \i[1027]  & \i[1025]  & \i[1026] ;
  assign new_n7742_ = ~new_n7714_ & (new_n7743_ | ~new_n6901_ | (\i[2991]  & (\i[2989]  | \i[2990] )));
  assign new_n7743_ = \i[2199]  & \i[2198]  & \i[2196]  & \i[2197] ;
  assign new_n7744_ = ~\i[1731]  & ~\i[1729]  & ~\i[1730] ;
  assign new_n7745_ = new_n7746_ & (new_n4659_ | ~new_n6407_ | ~new_n3771_ | ~\i[1285] );
  assign new_n7746_ = ~\i[511]  & ~\i[510]  & ~\i[508]  & ~\i[509] ;
  assign new_n7747_ = new_n7762_ ? (new_n3349_ ? new_n7757_ : new_n7759_) : new_n7748_;
  assign new_n7748_ = new_n7754_ ? ((~new_n7753_ & ~new_n7755_) | (~new_n7756_ & new_n6073_ & new_n7755_)) : new_n7749_;
  assign new_n7749_ = (new_n7752_ | new_n7751_) & (\i[1407]  | ~new_n7750_ | ~new_n7751_ | (\i[1406]  & \i[1405] ));
  assign new_n7750_ = ~\i[1951]  & (~\i[1950]  | (~\i[1949]  & ~\i[1948] ));
  assign new_n7751_ = ~\i[1627]  & ~\i[1626]  & ~\i[1624]  & ~\i[1625] ;
  assign new_n7752_ = (~\i[1077]  | ~\i[1078]  | ~\i[1079] ) & (~\i[1045]  | ~\i[1046]  | ~\i[1047] );
  assign new_n7753_ = (~\i[1099]  & (~\i[1097]  | ~\i[1098] )) ? new_n3696_ : new_n7744_;
  assign new_n7754_ = \i[1071]  & (\i[1069]  | \i[1070]  | \i[1068] );
  assign new_n7755_ = ~\i[1322]  & ~\i[1323]  & (~\i[1321]  | ~\i[1320] );
  assign new_n7756_ = ~\i[1399]  & (~\i[1397]  | ~\i[1398]  | ~\i[1396] );
  assign new_n7757_ = (new_n7758_ | ~new_n3368_) & (~\i[1847]  | new_n3368_ | (~\i[1846]  & (~\i[1844]  | ~\i[1845] )));
  assign new_n7758_ = (~new_n7487_ | ~new_n3659_) & (~\i[2613]  | ~\i[2614]  | ~\i[2615]  | new_n3659_);
  assign new_n7759_ = (new_n7760_ | ~new_n6240_) & (new_n7761_ | ~new_n4470_ | new_n6240_);
  assign new_n7760_ = new_n4788_ & (~\i[1255]  | (~\i[1254]  & (~\i[1253]  | ~\i[1252] )));
  assign new_n7761_ = ~\i[2735]  & (~\i[2734]  | (~\i[2733]  & ~\i[2732] ));
  assign new_n7762_ = ~\i[1067]  & (~\i[1065]  | ~\i[1066]  | ~\i[1064] );
  assign new_n7763_ = (new_n7775_ & (new_n5032_ ? ~new_n7764_ : ~new_n7768_)) | (~new_n7771_ & ~new_n7774_ & ~new_n7775_);
  assign new_n7764_ = new_n7731_ ? (new_n7766_ ? new_n4167_ : new_n7767_) : new_n7765_;
  assign new_n7765_ = (~\i[739]  | new_n6680_) & (\i[1258]  | \i[1259]  | ~new_n6680_ | (\i[1257]  & \i[1256] ));
  assign new_n7766_ = ~\i[1075]  & (~\i[1073]  | ~\i[1074]  | ~\i[1072] );
  assign new_n7767_ = ~\i[1547]  & (~\i[1546]  | ~\i[1545] );
  assign new_n7768_ = (~new_n5316_ | new_n4430_ | ~new_n7769_) & (new_n7769_ | (new_n4050_ ? new_n3445_ : ~new_n7770_));
  assign new_n7769_ = \i[2875]  & (\i[2873]  | \i[2874]  | \i[2872] );
  assign new_n7770_ = ~\i[2855]  & (~\i[2854]  | ~\i[2853] );
  assign new_n7771_ = new_n7772_ & ~new_n7773_ & new_n5440_;
  assign new_n7772_ = new_n4018_ & (\i[2741]  | \i[2742]  | \i[2743] );
  assign new_n7773_ = \i[727]  & (\i[726]  | \i[725] );
  assign new_n7774_ = ~new_n5440_ & new_n4973_ & (\i[1663]  | \i[1662]  | \i[1661] );
  assign new_n7775_ = ~\i[635]  & ~\i[633]  & ~\i[634] ;
  assign new_n7776_ = new_n7785_ & ((~new_n7777_ & new_n7786_) | (~new_n7782_ & ~new_n7784_ & ~new_n7786_));
  assign new_n7777_ = (new_n7423_ | ~new_n4019_ | new_n7780_) & (new_n7778_ | ~new_n7780_ | (new_n7781_ & ~new_n7779_));
  assign new_n7778_ = new_n7779_ & (\i[2865]  | \i[2866]  | \i[2867] );
  assign new_n7779_ = ~\i[1955]  & (~\i[1954]  | (~\i[1953]  & ~\i[1952] ));
  assign new_n7780_ = ~\i[1399]  & (~\i[1398]  | (~\i[1397]  & ~\i[1396] ));
  assign new_n7781_ = ~\i[1631]  & (~\i[1630]  | (~\i[1629]  & ~\i[1628] ));
  assign new_n7782_ = new_n4075_ & (new_n4659_ ? new_n7783_ : ~new_n7733_);
  assign new_n7783_ = ~\i[2423]  & ~\i[2421]  & ~\i[2422] ;
  assign new_n7784_ = ~new_n4075_ & ~new_n4069_ & ~\i[811]  & (~\i[810]  | (~\i[808]  & ~\i[809] ));
  assign new_n7785_ = ~\i[503]  & ~\i[502]  & ~\i[500]  & ~\i[501] ;
  assign new_n7786_ = ~\i[1735]  & ~\i[1734]  & ~\i[1732]  & ~\i[1733] ;
  assign new_n7787_ = new_n7788_ ? (~new_n7865_ ^ new_n7977_) : (new_n7865_ ^ new_n7977_);
  assign new_n7788_ = new_n7789_ ? (~new_n7844_ ^ new_n7852_) : (new_n7844_ ^ new_n7852_);
  assign new_n7789_ = new_n7790_ ? (new_n7815_ ^ new_n7735_) : (~new_n7815_ ^ new_n7735_);
  assign new_n7790_ = new_n7791_ ? (new_n7798_ ^ new_n7807_) : (~new_n7798_ ^ new_n7807_);
  assign new_n7791_ = (\i[1279]  & (\i[1276]  | \i[1277]  | \i[1278] )) ? new_n7795_ : new_n7792_;
  assign new_n7792_ = \i[1283]  ? new_n7794_ : ((~new_n4317_ & ~new_n4678_ & new_n4780_) | (~new_n7793_ & ~new_n4780_));
  assign new_n7793_ = new_n5423_ ? new_n7305_ : ~new_n5769_;
  assign new_n7794_ = new_n4805_ ? ~new_n3275_ : (~\i[2735]  | (~\i[2733]  & ~\i[2734] ));
  assign new_n7795_ = ~new_n7796_ & (new_n7797_ | ((~new_n3593_ | new_n3898_) & (new_n3490_ | new_n4651_ | ~new_n3898_)));
  assign new_n7796_ = new_n7797_ & (new_n7260_ | new_n3549_ | ~new_n4966_) & (~new_n5625_ | new_n3540_ | new_n4966_);
  assign new_n7797_ = ~\i[1623]  & (~\i[1622]  | (~\i[1621]  & ~\i[1620] ));
  assign new_n7798_ = \i[2315]  ? (new_n7804_ | (~new_n7744_ & new_n5843_ & new_n7806_)) : new_n7799_;
  assign new_n7799_ = new_n7762_ ? new_n7800_ : ((~new_n7385_ & ~new_n3550_ & new_n4195_) | (~new_n7803_ & ~new_n4195_));
  assign new_n7800_ = (new_n4029_ & (~\i[1060]  | ~\i[1061] )) ? new_n7802_ : new_n7801_;
  assign new_n7801_ = new_n5156_ ? ~new_n4211_ : new_n3437_;
  assign new_n7802_ = \i[1047]  ? ~new_n4317_ : new_n4062_;
  assign new_n7803_ = ~\i[1811]  & (~\i[1810]  | ~\i[1809] );
  assign new_n7804_ = ~new_n5664_ & ~new_n7806_ & ((\i[2758]  & \i[2759] ) ? ~new_n3233_ : ~new_n7805_);
  assign new_n7805_ = \i[1767]  & (\i[1766]  | (\i[1765]  & \i[1764] ));
  assign new_n7806_ = \i[2095]  & \i[2094]  & \i[2092]  & \i[2093] ;
  assign new_n7807_ = new_n7775_ ? new_n7808_ : ((new_n4390_ | new_n6074_ | ~\i[727] ) & (new_n7814_ | \i[727] ));
  assign new_n7808_ = new_n7555_ ? (new_n7809_ | (~new_n4141_ & new_n4132_ & new_n5763_)) : new_n7811_;
  assign new_n7809_ = new_n4141_ & ((~new_n7810_ & ~new_n4803_) | (~\i[1423]  & new_n4803_ & (~\i[1422]  | ~\i[1421] )));
  assign new_n7810_ = \i[2415]  & (\i[2414]  | (\i[2413]  & \i[2412] ));
  assign new_n7811_ = new_n7712_ ? (new_n4247_ ? new_n7812_ : new_n3624_) : new_n7813_;
  assign new_n7812_ = \i[1707]  & \i[1706]  & \i[1704]  & \i[1705] ;
  assign new_n7813_ = ~\i[1135]  & (~\i[1133]  | ~\i[1134]  | ~\i[1132] );
  assign new_n7814_ = new_n4301_ & new_n5005_;
  assign new_n7815_ = new_n7816_ ? (~new_n7825_ ^ new_n7834_) : (new_n7825_ ^ new_n7834_);
  assign new_n7816_ = new_n4020_ ? new_n7817_ : (\i[2323]  ? ~new_n7821_ : new_n7822_);
  assign new_n7817_ = new_n5256_ ? ~new_n7818_ : ((~new_n7820_ | ~new_n3741_) & (~new_n4724_ | ~new_n6773_ | new_n3741_));
  assign new_n7818_ = new_n7819_ & \i[2855]  & (~\i[1846]  | ~\i[1847] ) & (\i[2853]  | \i[2854] );
  assign new_n7819_ = new_n4335_ & (~\i[705]  | ~\i[704] );
  assign new_n7820_ = \i[1843]  & (~\i[1642]  | ~\i[1643]  | ~\i[1641] );
  assign new_n7821_ = ~new_n5794_ & new_n5230_ & ((~\i[2764]  & ~\i[2765] ) | ~\i[2767]  | ~\i[2766] );
  assign new_n7822_ = (new_n7824_ | ~new_n3510_ | ~new_n7823_) & (new_n4070_ | ~\i[2615]  | new_n7823_);
  assign new_n7823_ = \i[2279]  & (\i[2278]  | \i[2277] );
  assign new_n7824_ = \i[2607]  & (\i[2606]  | \i[2605] );
  assign new_n7825_ = new_n4968_ ? new_n7830_ : ((~\i[2602]  & ~\i[2603] ) ? ~new_n7826_ : new_n7833_);
  assign new_n7826_ = (~\i[831]  & (~\i[830]  | (~\i[828]  & ~\i[829] ))) ? new_n7828_ : new_n7827_;
  assign new_n7827_ = (~new_n5035_ & (~\i[973]  | ~\i[974]  | ~\i[975] )) | (~new_n7734_ & \i[973]  & \i[974]  & \i[975] );
  assign new_n7828_ = ~\i[702]  & ~\i[703]  & new_n7829_ & (~\i[701]  | ~\i[700] );
  assign new_n7829_ = ~\i[2947]  & ~\i[2946]  & ~\i[2944]  & ~\i[2945] ;
  assign new_n7830_ = (new_n7831_ | new_n6225_) & (new_n5051_ | new_n6910_ | \i[1422]  | \i[1423]  | ~new_n6225_);
  assign new_n7831_ = (~new_n5448_ & \i[2394]  & \i[2395]  & new_n5480_) | (~new_n5480_ & (new_n7832_ | ~new_n5726_));
  assign new_n7832_ = \i[947]  & (\i[946]  | (\i[945]  & \i[944] ));
  assign new_n7833_ = ~\i[647]  & ~\i[645]  & ~\i[646] ;
  assign new_n7834_ = ~new_n7838_ & (new_n7835_ | ~new_n4661_ | (new_n6393_ & (new_n7839_ | new_n7841_)));
  assign new_n7835_ = new_n7836_ & (new_n7837_ | ~new_n3778_ | (new_n5843_ & (\i[2042]  | \i[2043] )));
  assign new_n7836_ = ~new_n6393_ & ((new_n3268_ & (~\i[2510]  | ~\i[2511] )) | new_n3778_ | (~new_n4973_ & \i[2510]  & \i[2511] ));
  assign new_n7837_ = ~\i[2042]  & ~\i[2043]  & \i[1487]  & (\i[1486]  | \i[1485] );
  assign new_n7838_ = ~new_n4661_ & ((~new_n5822_ & ~new_n6971_ & ~new_n5665_) | (~\i[715]  & new_n4071_ & new_n5665_));
  assign new_n7839_ = new_n7840_ & (new_n3613_ ? ~new_n6151_ : ~new_n5413_);
  assign new_n7840_ = \i[2183]  & \i[2182]  & \i[2180]  & \i[2181] ;
  assign new_n7841_ = ~new_n7840_ & ((~new_n6361_ & new_n7843_) | (~\i[2824]  & ~\i[2825]  & new_n7842_ & ~new_n7843_));
  assign new_n7842_ = ~\i[2826]  & ~\i[2827] ;
  assign new_n7843_ = \i[2839]  & (\i[2837]  | \i[2838]  | \i[2836] );
  assign new_n7844_ = ~new_n7850_ & (~new_n7851_ | new_n7845_ | (~new_n7823_ & ~new_n7848_ & new_n4070_));
  assign new_n7845_ = ~new_n7846_ & new_n7823_ & (~new_n7824_ | (~\i[1203]  & new_n4062_) | (new_n7386_ & ~new_n4062_));
  assign new_n7846_ = ~new_n7824_ & ~new_n7847_ & (new_n3572_ | (\i[2211]  & (\i[2210]  | \i[2209] )));
  assign new_n7847_ = \i[2195]  & \i[2194]  & new_n3572_ & \i[2193] ;
  assign new_n7848_ = (~\i[2952]  & ~\i[2953]  & ~\i[2954]  & ~\i[2955]  & new_n4719_) | (new_n7849_ & ~new_n4719_);
  assign new_n7849_ = \i[1511]  & (\i[1510]  | \i[1509] );
  assign new_n7850_ = ~new_n7851_ & (~new_n4110_ | (~\i[1081]  & ~\i[1082]  & ~\i[1083] ));
  assign new_n7851_ = ~\i[2711]  & (~\i[2710]  | ~\i[2709] );
  assign new_n7852_ = new_n7864_ ? ((~new_n4994_ & new_n7863_) | (\i[2307]  & ~new_n7853_)) : new_n7856_;
  assign new_n7853_ = (new_n7854_ | \i[2974]  | \i[2975] ) & (new_n7855_ | new_n7274_ | (~\i[2974]  & ~\i[2975] ));
  assign new_n7854_ = new_n6306_ ? new_n5041_ : new_n7464_;
  assign new_n7855_ = ~\i[2311]  & (~\i[2310]  | (~\i[2309]  & ~\i[2308] ));
  assign new_n7856_ = (new_n7860_ | new_n7862_ | ~new_n7783_) & (new_n7857_ | new_n7859_ | new_n7783_);
  assign new_n7857_ = new_n5262_ & ((~\i[1261]  & ~\i[1262]  & ~\i[1263]  & new_n7858_) | (~new_n7517_ & ~new_n7858_));
  assign new_n7858_ = ~\i[1978]  & ~\i[1979]  & (~\i[1977]  | ~\i[1976] );
  assign new_n7859_ = ~new_n6910_ & ~new_n5262_ & ~new_n3565_;
  assign new_n7860_ = new_n7861_ & ~new_n3606_ & ~new_n3686_;
  assign new_n7861_ = \i[827]  & (\i[826]  | (\i[825]  & \i[824] ));
  assign new_n7862_ = ~new_n7861_ & new_n5428_ & (\i[2183]  | (\i[2180]  & \i[2181]  & \i[2182] ));
  assign new_n7863_ = ~new_n3782_ & ~\i[2307]  & (~\i[2207]  | ~\i[2206] );
  assign new_n7864_ = \i[2867]  & (\i[2865]  | \i[2866]  | \i[2864] );
  assign new_n7865_ = new_n7866_ ? (new_n7910_ ^ new_n7972_) : (~new_n7910_ ^ new_n7972_);
  assign new_n7866_ = new_n7867_ ? (new_n7896_ ^ new_n7906_) : (~new_n7896_ ^ new_n7906_);
  assign new_n7867_ = new_n7868_ ? (new_n7880_ ^ new_n7891_) : (~new_n7880_ ^ new_n7891_);
  assign new_n7868_ = ~new_n7869_ & (~new_n7775_ | (~new_n7877_ & (~new_n7875_ | new_n7874_)));
  assign new_n7869_ = (new_n7873_ | new_n4046_ | (new_n4078_ & \i[1957] )) & ~new_n7775_ & (new_n7870_ | ~new_n4078_ | ~\i[1957] );
  assign new_n7870_ = ~new_n7871_ & (~new_n7872_ | (\i[823]  & (\i[820]  | \i[821]  | \i[822] )));
  assign new_n7871_ = ~new_n4234_ & (new_n6074_ | ~\i[2731]  | (~\i[2730]  & (~\i[2728]  | ~\i[2729] )));
  assign new_n7872_ = new_n4234_ & (~\i[2736]  | ~\i[2737]  | ~\i[2738]  | ~\i[2739] );
  assign new_n7873_ = \i[1658]  & \i[1659]  & (\i[1657]  | \i[1656] );
  assign new_n7874_ = new_n4110_ & new_n3604_ & ~\i[2266]  & ~\i[2267] ;
  assign new_n7875_ = new_n5051_ & (~new_n7876_ | (\i[1884]  & \i[1885]  & \i[1886]  & \i[1887] ));
  assign new_n7876_ = ~\i[2708]  & ~\i[2709]  & ~\i[2710]  & ~\i[2711]  & (\i[2267]  | \i[2266] );
  assign new_n7877_ = ~new_n5051_ & (new_n7878_ ? (new_n4781_ | new_n4402_) : ~new_n7879_);
  assign new_n7878_ = \i[811]  & \i[810]  & \i[808]  & \i[809] ;
  assign new_n7879_ = ~\i[1099]  & ~\i[2886]  & ~\i[2887]  & (~\i[1098]  | ~\i[1097] );
  assign new_n7880_ = (new_n7884_ & ~\i[2315] ) | (~new_n7881_ & \i[2315]  & (~new_n7886_ | (~new_n7889_ & ~new_n7887_)));
  assign new_n7881_ = ~new_n3775_ & (~new_n7882_ | (\i[2223]  & (\i[2220]  | \i[2221]  | \i[2222] )));
  assign new_n7882_ = ~new_n7883_ & ~\i[803]  & (~\i[802]  | (~\i[800]  & ~\i[801] ));
  assign new_n7883_ = new_n6300_ & (\i[1541]  | \i[1540] );
  assign new_n7884_ = new_n7737_ ? ~new_n4058_ : (\i[927]  ? new_n7885_ : new_n7736_);
  assign new_n7885_ = (~\i[855]  | ~new_n4100_ | (~\i[854]  & (~\i[852]  | ~\i[853] ))) & (new_n6452_ | new_n4100_);
  assign new_n7886_ = new_n3775_ & (~new_n7888_ | ~new_n7887_ | (~\i[1626]  & (~\i[1624]  | ~\i[1625] )));
  assign new_n7887_ = \i[1983]  & (\i[1981]  | \i[1982]  | \i[1980] );
  assign new_n7888_ = ~\i[919]  & \i[1627]  & (~\i[918]  | ~\i[917] );
  assign new_n7889_ = (new_n5566_ | ~new_n7890_) & (\i[1475]  | new_n7890_ | (\i[1474]  & (\i[1472]  | \i[1473] )));
  assign new_n7890_ = \i[2759]  & \i[2757]  & \i[2758] ;
  assign new_n7891_ = new_n7785_ & (new_n5896_ ? (~\i[1939]  | new_n7894_) : new_n7892_);
  assign new_n7892_ = (new_n7893_ | (new_n5845_ ? ~new_n3432_ : new_n6543_)) & (~new_n4520_ | new_n3455_ | ~new_n7893_);
  assign new_n7893_ = ~\i[2519]  & (~\i[2518]  | (~\i[2517]  & ~\i[2516] ));
  assign new_n7894_ = ~new_n7895_ & (new_n5737_ | (\i[933]  & \i[934]  & \i[935] ));
  assign new_n7895_ = \i[933]  & \i[934]  & \i[935]  & (~\i[829]  | ~\i[828]  | ~new_n6885_);
  assign new_n7896_ = (~new_n7903_ & ~new_n7897_ & ~new_n7905_) | (new_n7905_ & (new_n6278_ ? ~new_n7901_ : ~new_n7899_));
  assign new_n7897_ = new_n7898_ & new_n7893_ & \i[2411]  & (\i[2410]  | \i[2409] );
  assign new_n7898_ = \i[1743]  & \i[1742]  & new_n4449_ & \i[1741] ;
  assign new_n7899_ = (new_n7900_ & ~new_n3524_) | (~new_n4132_ & new_n5778_ & new_n3524_);
  assign new_n7900_ = \i[2731]  & \i[2729]  & \i[2730]  & (\i[2849]  | \i[2848]  | ~new_n5624_);
  assign new_n7901_ = new_n7849_ ? new_n7902_ : ((~\i[2974]  & ~\i[2975]  & new_n4521_) | (new_n3275_ & ~new_n4521_));
  assign new_n7902_ = ~new_n3490_ & (\i[1039]  | (\i[1038]  & (\i[1037]  | \i[1036] )));
  assign new_n7903_ = new_n7904_ & \i[819]  & \i[818]  & ~new_n4666_ & ~\i[943] ;
  assign new_n7904_ = (~\i[942]  | ~\i[940]  | ~\i[941] ) & (~\i[2411]  | (~\i[2410]  & ~\i[2409] ));
  assign new_n7905_ = \i[2191]  & \i[2190]  & \i[2188]  & \i[2189] ;
  assign new_n7906_ = ~new_n7838_ & (~new_n4661_ | ((new_n7839_ | new_n7909_ | ~new_n6393_) & (new_n7907_ | new_n6393_)));
  assign new_n7907_ = new_n3778_ ? new_n7908_ : ((\i[2510]  & \i[2511] ) ? ~new_n4973_ : new_n3268_);
  assign new_n7908_ = (new_n5843_ & (\i[2042]  | \i[2043] )) | (\i[1487]  & ~\i[2042]  & ~\i[2043]  & (\i[1486]  | \i[1485] ));
  assign new_n7909_ = ~new_n7840_ & (new_n7843_ | (~\i[2824]  & ~\i[2825]  & new_n7842_));
  assign new_n7910_ = new_n7911_ ? (~new_n7943_ ^ new_n7906_) : (new_n7943_ ^ new_n7906_);
  assign new_n7911_ = new_n7912_ ? (~new_n7921_ ^ new_n7934_) : (new_n7921_ ^ new_n7934_);
  assign new_n7912_ = new_n6354_ ? new_n7913_ : ((new_n7916_ | ~new_n4074_) & (~new_n7918_ | ~\i[2735]  | new_n4074_));
  assign new_n7913_ = new_n5625_ ? new_n7914_ : ((new_n7915_ | ~new_n3594_) & (new_n5648_ | ~new_n4915_ | new_n3594_));
  assign new_n7914_ = (\i[2718]  | \i[2719]  | ~new_n4162_) & (new_n4162_ | (new_n3985_ ? ~new_n3993_ : ~new_n7080_));
  assign new_n7915_ = new_n3492_ ? new_n4437_ : new_n6605_;
  assign new_n7916_ = (~new_n6361_ | ~new_n7541_ | new_n4309_) & (~new_n4965_ | ~new_n7917_ | ~new_n4309_);
  assign new_n7917_ = \i[2723]  & \i[2722]  & \i[2720]  & \i[2721] ;
  assign new_n7918_ = new_n7920_ & new_n7919_ & (\i[2734]  | \i[2733]  | \i[2732] );
  assign new_n7919_ = ~\i[2714]  & ~\i[2715]  & (~\i[2713]  | ~\i[2712] );
  assign new_n7920_ = \i[2071]  & \i[2070]  & \i[2068]  & \i[2069] ;
  assign new_n7921_ = new_n7933_ ? new_n7922_ : ((new_n7926_ | new_n7930_ | ~new_n5625_) & (new_n7927_ | new_n5625_));
  assign new_n7922_ = new_n5571_ ? (new_n7925_ | (~new_n5316_ & new_n6740_)) : new_n7923_;
  assign new_n7923_ = (~new_n7924_ | ~new_n4317_) & (new_n4890_ | ~new_n5625_ | new_n4317_);
  assign new_n7924_ = ~\i[1835]  & (~\i[1834]  | (~\i[1833]  & ~\i[1832] ));
  assign new_n7925_ = ~\i[2975]  & ~\i[2974]  & ~\i[2972]  & ~\i[2973] ;
  assign new_n7926_ = new_n4109_ & ~new_n4131_ & ~new_n3650_;
  assign new_n7927_ = (new_n7928_ | new_n7929_) & (new_n4463_ | new_n4065_ | ~new_n7929_);
  assign new_n7928_ = ~\i[927]  & ~\i[926]  & (~\i[1259]  | (~\i[1256]  & ~\i[1257]  & ~\i[1258] ));
  assign new_n7929_ = ~\i[1383]  & ~\i[1381]  & ~\i[1382] ;
  assign new_n7930_ = ~new_n4109_ & (new_n7931_ ? (\i[1527]  | (\i[1525]  & \i[1526] )) : ~new_n7932_);
  assign new_n7931_ = ~\i[931]  & (~\i[930]  | (~\i[929]  & ~\i[928] ));
  assign new_n7932_ = ~\i[1095]  & (~\i[1094]  | (~\i[1093]  & ~\i[1092] ));
  assign new_n7933_ = ~\i[2963]  & ~\i[2962]  & ~\i[2960]  & ~\i[2961] ;
  assign new_n7934_ = new_n3299_ ? new_n7938_ : ((new_n7935_ | ~new_n4985_) & (~new_n6892_ | ~new_n7942_ | new_n4985_));
  assign new_n7935_ = (~new_n7936_ | new_n3756_) & (~new_n4373_ | ~new_n7746_ | ~new_n3756_);
  assign new_n7936_ = \i[1659]  & \i[1658]  & new_n7937_ & \i[1657] ;
  assign new_n7937_ = ~\i[851]  & \i[1656]  & (~\i[850]  | ~\i[849] );
  assign new_n7938_ = (new_n7939_ | new_n7941_ | new_n5625_) & (new_n6519_ | ~new_n5625_ | (new_n5684_ & ~new_n5066_));
  assign new_n7939_ = ~new_n3221_ & (~new_n7940_ | (\i[1619]  & (\i[1618]  | (\i[1616]  & \i[1617] ))));
  assign new_n7940_ = \i[1475]  & (\i[1474]  | (\i[1473]  & \i[1472] ));
  assign new_n7941_ = ~new_n4373_ & new_n3221_ & (~\i[2071]  | ~\i[2070] );
  assign new_n7942_ = new_n7890_ & (\i[621]  | ~new_n5675_);
  assign new_n7943_ = new_n7944_ ? (~new_n7957_ ^ new_n7966_) : (new_n7957_ ^ new_n7966_);
  assign new_n7944_ = new_n5436_ ? (new_n4819_ ? new_n7951_ : new_n7955_) : new_n7945_;
  assign new_n7945_ = new_n5626_ ? new_n7946_ : ((new_n7949_ | new_n7950_) & (~new_n3775_ | ~new_n4779_ | ~new_n7950_));
  assign new_n7946_ = (new_n4036_ | ~new_n6252_ | ~new_n4664_) & (new_n7947_ | ~new_n7948_ | new_n4664_);
  assign new_n7947_ = \i[822]  & \i[823]  & (\i[821]  | \i[820] );
  assign new_n7948_ = \i[927]  & \i[926]  & \i[924]  & \i[925] ;
  assign new_n7949_ = (new_n7770_ | new_n3326_) & (~\i[2641]  | ~\i[2642]  | ~\i[2643]  | ~new_n3326_);
  assign new_n7950_ = ~\i[1739]  & (~\i[1738]  | (~\i[1737]  & ~\i[1736] ));
  assign new_n7951_ = new_n7954_ ? (new_n5684_ ? ~new_n7555_ : ~new_n6120_) : new_n7952_;
  assign new_n7952_ = ~new_n7953_ & (~\i[1035]  | ~\i[2191]  | (~\i[1034]  & (~\i[1033]  | ~\i[1032] )));
  assign new_n7953_ = ~\i[2191]  & (~\i[2879]  | (~\i[2877]  & ~\i[2878] ));
  assign new_n7954_ = ~\i[2435]  & (~\i[2434]  | ~\i[2433] );
  assign new_n7955_ = (~new_n7956_ | ~new_n6473_) & (new_n4425_ | ~\i[2487]  | new_n6473_ | (~\i[2486]  & ~\i[2485] ));
  assign new_n7956_ = (\i[1039]  | (\i[1038]  & \i[1037] )) & (~\i[827]  | ~\i[826] );
  assign new_n7957_ = (new_n7963_ | new_n7965_ | new_n3549_) & (new_n7958_ | new_n7962_ | ~new_n3549_);
  assign new_n7958_ = new_n4206_ & (new_n4768_ ? (new_n3988_ ? new_n7961_ : new_n5513_) : ~new_n7959_);
  assign new_n7959_ = (new_n3749_ | ~new_n7960_) & (\i[2841]  | \i[2842]  | \i[2843]  | new_n7960_);
  assign new_n7960_ = \i[2715]  & (\i[2714]  | (\i[2713]  & \i[2712] ));
  assign new_n7961_ = ~\i[2063]  & (~\i[2062]  | (~\i[2061]  & ~\i[2060] ));
  assign new_n7962_ = ~new_n4206_ & (new_n6899_ ? new_n3555_ : (new_n3451_ ? new_n3564_ : ~new_n6001_));
  assign new_n7963_ = (new_n4147_ | ~new_n4661_ | ~new_n7964_) & (~new_n3258_ | new_n7964_ | (\i[1847]  & \i[1846] ));
  assign new_n7964_ = ~\i[735]  & (~\i[734]  | ~\i[733] );
  assign new_n7965_ = ~\i[1646]  & ~\i[1647]  & (~\i[1645]  | ~\i[1644] );
  assign new_n7966_ = new_n4063_ & (new_n6839_ ? ~new_n7967_ : ~new_n7970_);
  assign new_n7967_ = (~new_n7968_ | ~new_n3365_ | new_n7235_) & (~new_n7235_ | (new_n7969_ ? new_n4093_ : ~new_n5571_));
  assign new_n7968_ = ~\i[2995]  & ~\i[2994]  & ~\i[2992]  & ~\i[2993] ;
  assign new_n7969_ = \i[1087]  & \i[1085]  & \i[1086] ;
  assign new_n7970_ = (new_n7971_ | new_n4147_) & (\i[1399]  | ~new_n4147_ | (\i[1415]  & (\i[1413]  | \i[1414] )));
  assign new_n7971_ = ~\i[2255]  & ~\i[2254]  & ~\i[2253]  & ~\i[594]  & ~\i[595] ;
  assign new_n7972_ = new_n3735_ & (new_n3275_ ? ~new_n7973_ : (\i[1607]  ? ~new_n7975_ : ~new_n7976_));
  assign new_n7973_ = new_n4340_ ? ((\i[1398]  | \i[1399]  | ~new_n5138_) & (~new_n7961_ | new_n5138_)) : new_n7974_;
  assign new_n7974_ = new_n4437_ ? ~new_n6966_ : (~new_n3771_ | (~\i[1284]  & ~\i[1285] ));
  assign new_n7975_ = new_n5041_ ? (~\i[1623]  | (~\i[1621]  & ~\i[1622] )) : ~new_n4086_;
  assign new_n7976_ = (new_n3241_ | new_n3243_) & (~\i[1734]  | ~\i[1735]  | ~new_n3243_);
  assign new_n7977_ = (new_n7978_ & new_n7762_) | (~new_n7983_ & ~new_n7762_ & (~new_n4195_ | (~new_n7987_ & ~new_n7988_)));
  assign new_n7978_ = (new_n7979_ | new_n6446_) & (new_n4735_ | ~new_n6446_ | (new_n7982_ ? new_n7770_ : ~new_n3775_));
  assign new_n7979_ = (~\i[1051]  & (~\i[1049]  | ~\i[1050] )) ? new_n7981_ : ~new_n7980_;
  assign new_n7980_ = \i[2871]  & new_n3664_ & \i[2870] ;
  assign new_n7981_ = new_n4207_ ? ~new_n4703_ : ~new_n7372_;
  assign new_n7982_ = ~\i[1879]  & (~\i[1878]  | ~new_n5396_);
  assign new_n7983_ = ~new_n4195_ & (new_n7986_ ? ~new_n7984_ : (new_n7985_ | new_n7744_));
  assign new_n7984_ = (~\i[807]  & \i[2102]  & \i[2103]  & (~\i[806]  | ~\i[805] )) | (new_n5522_ & (~\i[2102]  | ~\i[2103] ));
  assign new_n7985_ = \i[2171]  & (\i[2169]  | \i[2170]  | \i[2168] );
  assign new_n7986_ = \i[1635]  & (\i[1633]  | \i[1634]  | \i[1632] );
  assign new_n7987_ = (\i[590]  | \i[591]  | (\i[2734]  & \i[2735] )) & ~new_n6906_ & (~new_n4953_ | ~\i[2734]  | ~\i[2735] );
  assign new_n7988_ = new_n7989_ & new_n4369_ & new_n6906_;
  assign new_n7989_ = ~\i[1863]  & (~\i[1862]  | (~\i[1861]  & ~\i[1860] ));
  assign new_n7990_ = (new_n7994_ | ~new_n3899_) & (new_n7992_ | new_n3899_ | (new_n7991_ & (new_n7919_ | ~new_n6308_)));
  assign new_n7991_ = ~new_n4074_ & (~\i[2707]  | (~\i[2704]  & ~\i[2705]  & ~\i[2706] ));
  assign new_n7992_ = new_n4074_ & (new_n7993_ | \i[1407]  | (new_n5559_ & (~\i[916]  | ~\i[917] )));
  assign new_n7993_ = \i[2727]  & (\i[2726]  | \i[2725] );
  assign new_n7994_ = (new_n7998_ | ~new_n7999_ | new_n7541_) & (new_n7995_ | new_n7996_ | ~new_n7541_);
  assign new_n7995_ = ~new_n3242_ & ~new_n4288_ & ~\i[2167]  & (~\i[2166]  | ~\i[2165] );
  assign new_n7996_ = new_n3242_ & (\i[1145]  | \i[1146]  | \i[1147]  | ~new_n7997_);
  assign new_n7997_ = ~\i[715]  & ~\i[714]  & ~\i[712]  & ~\i[713] ;
  assign new_n7998_ = (new_n5031_ | ~new_n4019_) & (~\i[2867]  | new_n4019_ | (~\i[2866]  & (~\i[2864]  | ~\i[2865] )));
  assign new_n7999_ = ~\i[2875]  & ~\i[2873]  & ~\i[2874] ;
  assign new_n8000_ = new_n3494_ ? new_n8001_ : ((new_n8011_ | ~new_n8009_) & (~new_n8007_ | new_n8010_));
  assign new_n8001_ = new_n3233_ ? (~new_n8005_ & (new_n3413_ | new_n4206_ | ~new_n4275_)) : new_n8002_;
  assign new_n8002_ = ~new_n8004_ & (~new_n8003_ | (~new_n5770_ & (\i[1151]  | (\i[1149]  & \i[1150] ))));
  assign new_n8003_ = (\i[1363]  | \i[1361]  | \i[1362] ) & (~new_n5770_ | ~\i[1366]  | ~\i[1367] );
  assign new_n8004_ = ~\i[1361]  & ~\i[1362]  & ~\i[1363]  & (new_n3373_ ? new_n3754_ : new_n3898_);
  assign new_n8005_ = new_n3413_ & ~new_n8006_ & new_n4134_;
  assign new_n8006_ = ~\i[1707]  & ~\i[1705]  & ~\i[1706] ;
  assign new_n8007_ = ~new_n8008_ & new_n6885_ & new_n4985_ & (\i[829]  | \i[828] );
  assign new_n8008_ = new_n4803_ & (\i[2749]  | \i[2748] );
  assign new_n8009_ = ~new_n4985_ & ~\i[2515]  & \i[590]  & \i[591]  & (~\i[2514]  | new_n3776_);
  assign new_n8010_ = \i[727]  & (\i[725]  | \i[726]  | \i[724] );
  assign new_n8011_ = \i[923]  & (\i[922]  | (\i[921]  & \i[920] ));
  assign \o[50]  = new_n8013_ ^ new_n8115_;
  assign new_n8013_ = new_n8014_ ? (~new_n8113_ ^ new_n8114_) : (new_n8113_ ^ new_n8114_);
  assign new_n8014_ = new_n8015_ ? (~new_n8093_ ^ new_n8094_) : (new_n8093_ ^ new_n8094_);
  assign new_n8015_ = new_n8016_ ? (~new_n8066_ ^ new_n8067_) : (new_n8066_ ^ new_n8067_);
  assign new_n8016_ = new_n8017_ ? (~new_n8053_ ^ new_n8065_) : (new_n8053_ ^ new_n8065_);
  assign new_n8017_ = new_n8018_ ? (~new_n8037_ ^ new_n8038_) : (new_n8037_ ^ new_n8038_);
  assign new_n8018_ = new_n8019_ ? (new_n8027_ ^ new_n8031_) : (~new_n8027_ ^ new_n8031_);
  assign new_n8019_ = new_n3549_ ? (new_n4206_ ? ~new_n8026_ : ~new_n8024_) : new_n8020_;
  assign new_n8020_ = new_n7965_ ? new_n8021_ : new_n8023_;
  assign new_n8021_ = (new_n8022_ | ~new_n4078_ | (~\i[1956]  & ~\i[1957] )) & (\i[1623]  | new_n4865_ | (new_n4078_ & (\i[1956]  | \i[1957] )));
  assign new_n8022_ = (~new_n4985_ | new_n4119_) & (~\i[1046]  | ~\i[1047]  | ~new_n4119_);
  assign new_n8023_ = new_n7964_ ? ~new_n4661_ : ((\i[1846]  & \i[1847] ) ? ~new_n5102_ : ~new_n3258_);
  assign new_n8024_ = (new_n6001_ | new_n3451_ | new_n6899_) & (new_n8025_ | \i[2711]  | ~new_n3555_ | ~new_n6899_);
  assign new_n8025_ = \i[2710]  & (\i[2709]  | \i[2708] );
  assign new_n8026_ = (new_n7960_ | new_n4768_) & (new_n3988_ | ~new_n5513_ | ~new_n4768_);
  assign new_n8027_ = (new_n8030_ | ~new_n4074_ | new_n3899_) & (~new_n3899_ | (~new_n8029_ & (~new_n7541_ | new_n8028_)));
  assign new_n8028_ = ~new_n7995_ & (~new_n7996_ | (~new_n6956_ & (\i[1145]  | ~new_n5810_)));
  assign new_n8029_ = ~new_n7541_ & ~new_n7999_ & (new_n4206_ ? ~\i[2071]  : ~new_n3513_);
  assign new_n8030_ = (~new_n4723_ | ~new_n7993_ | \i[1407] ) & (~\i[1407]  | (new_n3549_ ? ~new_n3996_ : ~new_n5398_));
  assign new_n8031_ = (new_n8033_ | new_n8032_ | new_n6354_) & (~new_n6354_ | (new_n5625_ ? new_n8034_ : new_n8035_));
  assign new_n8032_ = new_n4074_ & (~new_n4704_ | new_n4965_ | ~new_n4309_) & (new_n6361_ | ~new_n7541_ | new_n4309_);
  assign new_n8033_ = ~new_n4074_ & (new_n7919_ | (~new_n5262_ & (~\i[599]  | ~\i[598] )));
  assign new_n8034_ = (new_n4111_ | ~new_n4162_ | (~\i[2719]  & ~\i[2718] )) & (new_n7080_ | new_n3985_ | new_n4162_);
  assign new_n8035_ = (new_n8036_ | ~new_n5648_ | ~\i[2955]  | new_n3594_) & (~new_n3492_ | ~new_n4437_ | ~new_n3594_);
  assign new_n8036_ = ~\i[2954]  & (~\i[2953]  | ~\i[2952] );
  assign new_n8037_ = (~new_n7921_ & ~new_n7934_) | (~new_n7912_ & (~new_n7921_ | ~new_n7934_));
  assign new_n8038_ = new_n8039_ ? (~new_n8043_ ^ new_n8048_) : (new_n8043_ ^ new_n8048_);
  assign new_n8039_ = new_n7933_ ? new_n8042_ : new_n8040_;
  assign new_n8040_ = new_n5625_ ? ((new_n4131_ & new_n4109_) | (~new_n7931_ & ~new_n7932_ & ~new_n4109_)) : new_n8041_;
  assign new_n8041_ = (\i[926]  | \i[927]  | new_n7929_) & (new_n4065_ | ~new_n4463_ | ~new_n7929_);
  assign new_n8042_ = new_n4317_ & ((~new_n7925_ & new_n5316_ & new_n5571_) | (new_n3548_ & new_n7924_ & ~new_n5571_));
  assign new_n8043_ = (new_n8044_ & new_n3494_) | (~new_n8046_ & ~new_n3494_ & (~new_n8011_ | ~new_n8047_));
  assign new_n8044_ = new_n3233_ ? new_n8045_ : (new_n5770_ | (~\i[1361]  & ~\i[1362]  & ~\i[1363] ));
  assign new_n8045_ = (~new_n8006_ | ~new_n6254_ | ~new_n3413_) & (\i[2170]  | \i[2171]  | ~new_n4206_ | new_n3413_);
  assign new_n8046_ = new_n4985_ & ((new_n3284_ & new_n7098_ & new_n8010_) | (new_n8008_ & new_n6232_ & ~new_n8010_));
  assign new_n8047_ = ~new_n4985_ & ~\i[2319]  & new_n4335_ & (~\i[2318]  | (~\i[2316]  & ~\i[2317] ));
  assign new_n8048_ = new_n3299_ ? ((new_n8050_ | ~new_n5625_) & (new_n7939_ | new_n8052_ | new_n5625_)) : ~new_n8049_;
  assign new_n8049_ = new_n7890_ & ~\i[623]  & ~\i[622]  & ~new_n4985_ & ~\i[621] ;
  assign new_n8050_ = (~new_n5176_ | new_n5684_ | new_n6519_) & (~new_n6519_ | (new_n8051_ & (\i[2270]  | \i[2271] )));
  assign new_n8051_ = ~\i[2987]  & ~\i[2985]  & ~\i[2986] ;
  assign new_n8052_ = new_n3221_ & (~new_n4373_ | ~new_n4379_ | ~\i[1073] );
  assign new_n8053_ = new_n8054_ ? (new_n8055_ ^ new_n8064_) : (~new_n8055_ ^ new_n8064_);
  assign new_n8054_ = (~new_n7880_ & new_n7891_) | (~new_n7868_ & (~new_n7880_ | new_n7891_));
  assign new_n8055_ = new_n8056_ ? (~new_n8061_ ^ new_n8063_) : (new_n8061_ ^ new_n8063_);
  assign new_n8056_ = (~new_n8059_ & ~new_n7774_ & ~new_n7775_) | (new_n7775_ & (new_n5032_ ? new_n8058_ : new_n8057_));
  assign new_n8057_ = (~new_n3445_ | ~new_n4050_ | new_n7769_) & (~new_n7769_ | (new_n5316_ ? ~new_n4430_ : ~new_n7213_));
  assign new_n8058_ = new_n7731_ ? (new_n7766_ ? ~new_n4167_ : ~new_n7767_) : ~new_n7765_;
  assign new_n8059_ = new_n5440_ & ((new_n7772_ & ~new_n7773_) | (new_n4087_ & new_n8060_ & new_n7773_));
  assign new_n8060_ = ~\i[2306]  & ~\i[2307]  & (~\i[2305]  | ~\i[2304] );
  assign new_n8061_ = new_n7785_ & (new_n7786_ ? (new_n7780_ ? new_n7778_ : ~new_n8062_) : new_n7782_);
  assign new_n8062_ = new_n4019_ ? ~new_n7423_ : new_n3395_;
  assign new_n8063_ = new_n4063_ & new_n3473_ & new_n6839_ & ~new_n7235_ & ~new_n7968_;
  assign new_n8064_ = (new_n7957_ & new_n7966_) | (~new_n7944_ & (new_n7957_ | new_n7966_));
  assign new_n8065_ = (~new_n7943_ & ~new_n7906_) | (~new_n7911_ & (~new_n7943_ | ~new_n7906_));
  assign new_n8066_ = (~new_n7910_ & new_n7972_) | (~new_n7866_ & (~new_n7910_ | new_n7972_));
  assign new_n8067_ = new_n8068_ ? (new_n8069_ ^ new_n8092_) : (~new_n8069_ ^ new_n8092_);
  assign new_n8068_ = (~new_n7815_ & new_n7735_) | (~new_n7790_ & (~new_n7815_ | new_n7735_));
  assign new_n8069_ = new_n8070_ ? (new_n8071_ ^ new_n8084_) : (~new_n8071_ ^ new_n8084_);
  assign new_n8070_ = (new_n7825_ & new_n7834_) | (~new_n7816_ & (new_n7825_ | new_n7834_));
  assign new_n8071_ = new_n8072_ ? (new_n8077_ ^ new_n8082_) : (~new_n8077_ ^ new_n8082_);
  assign new_n8072_ = new_n5436_ ? ((~new_n6473_ | ~new_n8076_) & (~new_n7953_ | ~new_n8075_)) : new_n8073_;
  assign new_n8073_ = (~new_n7947_ | ~new_n8074_ | ~new_n5626_) & (new_n7770_ | new_n3326_ | new_n7950_ | new_n5626_);
  assign new_n8074_ = ~\i[2659]  & ~\i[2658]  & ~new_n4664_ & ~\i[2657] ;
  assign new_n8075_ = ~new_n7954_ & new_n4819_;
  assign new_n8076_ = \i[827]  & \i[826]  & ~new_n4819_ & new_n3365_;
  assign new_n8077_ = (new_n7762_ & (~new_n6446_ | new_n8078_)) | (~new_n8081_ & ~new_n8080_ & ~new_n7762_);
  assign new_n8078_ = ~new_n8079_ & (new_n7770_ | new_n4735_ | \i[1879]  | (\i[1878]  & new_n5396_));
  assign new_n8079_ = new_n4735_ & new_n3229_ & (\i[2963]  | (\i[2962]  & (\i[2961]  | \i[2960] )));
  assign new_n8080_ = new_n7989_ & new_n6906_ & ~new_n4369_ & new_n4195_;
  assign new_n8081_ = new_n7985_ & ~new_n7986_ & ~new_n4195_ & ~new_n6252_;
  assign new_n8082_ = ~new_n8083_ & (new_n5051_ | \i[723]  | ~new_n7775_ | ~new_n7878_ | ~new_n4781_);
  assign new_n8083_ = \i[1959]  & \i[1958]  & \i[1957]  & new_n6074_ & ~new_n4234_ & ~new_n7775_;
  assign new_n8084_ = new_n8085_ ? (~new_n8088_ ^ new_n8090_) : (new_n8088_ ^ new_n8090_);
  assign new_n8085_ = ~new_n7850_ & (~new_n7851_ | (~new_n8086_ & new_n7823_) | (new_n4070_ & new_n8087_ & ~new_n7823_));
  assign new_n8086_ = (~new_n7847_ | new_n7824_) & (new_n4062_ | ~new_n7386_ | ~new_n7824_);
  assign new_n8087_ = ~new_n4719_ & ~new_n7849_;
  assign new_n8088_ = ~new_n3652_ & (new_n8089_ | (~new_n7714_ & new_n6110_ & new_n7744_ & new_n7743_));
  assign new_n8089_ = new_n7360_ & new_n5316_ & new_n7714_ & ~\i[2630]  & ~\i[2631] ;
  assign new_n8090_ = ~new_n8091_ & new_n7785_;
  assign new_n8091_ = (new_n7893_ | ~new_n5845_ | ~new_n3432_ | new_n5896_) & (~\i[1939]  | ~new_n7895_ | ~new_n5896_);
  assign new_n8092_ = (~new_n7906_ & new_n7896_) | (~new_n7867_ & (~new_n7906_ | new_n7896_));
  assign new_n8093_ = (~new_n7865_ & ~new_n7977_) | (~new_n7788_ & (~new_n7865_ | ~new_n7977_));
  assign new_n8094_ = new_n8095_ ? (new_n8096_ ^ new_n8112_) : (~new_n8096_ ^ new_n8112_);
  assign new_n8095_ = (~new_n7747_ & new_n7738_) | (~new_n7697_ & (~new_n7747_ | new_n7738_));
  assign new_n8096_ = new_n8097_ ? (new_n8098_ ^ new_n8109_) : (~new_n8098_ ^ new_n8109_);
  assign new_n8097_ = (new_n7723_ & new_n7735_) | (~new_n7698_ & (new_n7723_ | new_n7735_));
  assign new_n8098_ = new_n8099_ ? (new_n8100_ ^ new_n8101_) : (~new_n8100_ ^ new_n8101_);
  assign new_n8099_ = (~new_n7798_ & new_n7807_) | (~new_n7791_ & (~new_n7798_ | new_n7807_));
  assign new_n8100_ = (~new_n7706_ & new_n7715_) | (~new_n7699_ & (~new_n7706_ | new_n7715_));
  assign new_n8101_ = new_n8102_ ? (new_n8105_ ^ new_n8107_) : (~new_n8105_ ^ new_n8107_);
  assign new_n8102_ = new_n4020_ ? new_n8103_ : (\i[2323]  ? new_n7821_ : ~new_n7822_);
  assign new_n8103_ = new_n5256_ ? (new_n7818_ | (~new_n7819_ & new_n5497_)) : new_n8104_;
  assign new_n8104_ = new_n3741_ ? new_n7820_ : (new_n4724_ ? new_n6773_ : new_n3548_);
  assign new_n8105_ = (~new_n8106_ | ~new_n7864_) & (~new_n7862_ | ~new_n7783_ | new_n7864_);
  assign new_n8106_ = \i[2307]  & ~\i[2975]  & ~\i[2974]  & ~new_n6306_ & ~new_n7464_;
  assign new_n8107_ = new_n8108_ & new_n6848_ & ~new_n7258_ & new_n5422_;
  assign new_n8108_ = new_n3940_ & \i[1167]  & ~\i[1843]  & \i[1166] ;
  assign new_n8109_ = ~new_n8110_ & new_n7905_;
  assign new_n8110_ = new_n6278_ ? new_n8111_ : ((~new_n7900_ | new_n3524_) & (new_n4132_ | ~new_n5778_ | ~new_n3524_));
  assign new_n8111_ = new_n7849_ ? ~new_n7902_ : ((\i[2974]  | \i[2975]  | ~new_n4521_) & (~new_n3275_ | new_n4521_));
  assign new_n8112_ = (~new_n7844_ & ~new_n7852_) | (~new_n7789_ & (~new_n7844_ | ~new_n7852_));
  assign new_n8113_ = (~new_n7787_ & ~new_n7990_) | (~new_n7695_ & (~new_n7787_ | ~new_n7990_));
  assign new_n8114_ = (new_n7763_ & new_n7776_) | (~new_n7696_ & (new_n7763_ | new_n7776_));
  assign new_n8115_ = ~new_n7694_ & ~new_n8000_;
  assign \o[51]  = ~new_n8117_ ^ new_n8118_;
  assign new_n8117_ = new_n8013_ & new_n8115_;
  assign new_n8118_ = new_n8119_ ^ new_n8120_;
  assign new_n8119_ = (new_n8113_ & new_n8114_) | (new_n8014_ & (new_n8113_ | new_n8114_));
  assign new_n8120_ = new_n8121_ ? (~new_n8122_ ^ new_n8156_) : (new_n8122_ ^ new_n8156_);
  assign new_n8121_ = (new_n8093_ & new_n8094_) | (new_n8015_ & (new_n8093_ | new_n8094_));
  assign new_n8122_ = new_n8123_ ? (new_n8124_ ^ new_n8148_) : (~new_n8124_ ^ new_n8148_);
  assign new_n8123_ = (new_n8066_ & new_n8067_) | (new_n8016_ & (new_n8066_ | new_n8067_));
  assign new_n8124_ = new_n8125_ ? (new_n8126_ ^ new_n8144_) : (~new_n8126_ ^ new_n8144_);
  assign new_n8125_ = (new_n8053_ & new_n8065_) | (new_n8017_ & (new_n8053_ | new_n8065_));
  assign new_n8126_ = new_n8127_ ? (new_n8130_ ^ new_n8131_) : (~new_n8130_ ^ new_n8131_);
  assign new_n8127_ = ~new_n8128_ ^ new_n8129_;
  assign new_n8128_ = (~new_n8027_ & ~new_n8031_) | (~new_n8019_ & (~new_n8027_ | ~new_n8031_));
  assign new_n8129_ = (new_n8061_ & new_n8063_) | (~new_n8056_ & (new_n8061_ | new_n8063_));
  assign new_n8130_ = (new_n8037_ & new_n8038_) | (new_n8018_ & (new_n8037_ | new_n8038_));
  assign new_n8131_ = new_n8132_ ? (~new_n8142_ ^ new_n8143_) : (new_n8142_ ^ new_n8143_);
  assign new_n8132_ = new_n8133_ ? (new_n8140_ ^ new_n8141_) : (~new_n8140_ ^ new_n8141_);
  assign new_n8133_ = ~new_n8134_ & (~new_n7933_ | (new_n8136_ & ~new_n5571_) | (new_n8138_ & new_n5571_));
  assign new_n8134_ = ~new_n7933_ & (new_n8135_ | ~new_n5625_) & (new_n3696_ | ~new_n4065_ | ~new_n7929_ | new_n5625_);
  assign new_n8135_ = (new_n7931_ | ~new_n7932_ | new_n4109_) & (~new_n4109_ | (new_n4131_ ? ~new_n4134_ : ~new_n3650_));
  assign new_n8136_ = new_n4317_ ? (new_n7924_ ? new_n3548_ : new_n4275_) : new_n8137_;
  assign new_n8137_ = new_n4890_ & ~\i[1387]  & ~\i[1385]  & ~\i[1386] ;
  assign new_n8138_ = (new_n5316_ & (new_n7925_ ? ~new_n5896_ : new_n4317_)) | (~new_n8139_ & new_n5896_ & new_n7925_) | (~new_n6740_ & ~new_n5316_ & ~new_n7925_);
  assign new_n8139_ = ~\i[1135]  & ~\i[1134]  & ~\i[1132]  & ~\i[1133] ;
  assign new_n8140_ = new_n6473_ & new_n8076_ & new_n5436_;
  assign new_n8141_ = new_n8139_ & new_n3299_ & new_n6519_ & ~new_n8051_ & new_n5625_;
  assign new_n8142_ = (~new_n8043_ & ~new_n8048_) | (new_n8039_ & (~new_n8043_ | ~new_n8048_));
  assign new_n8143_ = ~new_n7762_ & new_n8080_;
  assign new_n8144_ = new_n8145_ ? (new_n8146_ ^ new_n8147_) : (~new_n8146_ ^ new_n8147_);
  assign new_n8145_ = (~new_n8055_ & new_n8064_) | (new_n8054_ & (~new_n8055_ | new_n8064_));
  assign new_n8146_ = (new_n8071_ & new_n8084_) | (new_n8070_ & (new_n8071_ | new_n8084_));
  assign new_n8147_ = (~new_n8082_ & new_n8077_) | (new_n8072_ & (~new_n8082_ | new_n8077_));
  assign new_n8148_ = new_n8149_ ? (~new_n8150_ ^ new_n8155_) : (new_n8150_ ^ new_n8155_);
  assign new_n8149_ = (new_n8098_ & new_n8109_) | (new_n8097_ & (new_n8098_ | new_n8109_));
  assign new_n8150_ = new_n8151_ ^ new_n8152_;
  assign new_n8151_ = (~new_n8101_ & new_n8100_) | (new_n8099_ & (~new_n8101_ | new_n8100_));
  assign new_n8152_ = ~new_n8153_ ^ new_n8154_;
  assign new_n8153_ = (~new_n8105_ & new_n8107_) | (~new_n8102_ & (~new_n8105_ | new_n8107_));
  assign new_n8154_ = (new_n8088_ & new_n8090_) | (new_n8085_ & (new_n8088_ | new_n8090_));
  assign new_n8155_ = (~new_n8069_ & new_n8092_) | (new_n8068_ & (~new_n8069_ | new_n8092_));
  assign new_n8156_ = (~new_n8096_ & new_n8112_) | (new_n8095_ & (~new_n8096_ | new_n8112_));
  assign \o[52]  = ((new_n8158_ | new_n8159_) & (~new_n8160_ ^ ~new_n8161_)) | (~new_n8158_ & ~new_n8159_ & (~new_n8160_ ^ new_n8161_));
  assign new_n8158_ = ~new_n8118_ & new_n8117_;
  assign new_n8159_ = ~new_n8120_ & new_n8119_;
  assign new_n8160_ = (~new_n8122_ & new_n8156_) | (new_n8121_ & (~new_n8122_ | new_n8156_));
  assign new_n8161_ = new_n8162_ ? (~new_n8163_ ^ new_n8175_) : (new_n8163_ ^ new_n8175_);
  assign new_n8162_ = (~new_n8124_ & ~new_n8148_) | (new_n8123_ & (~new_n8124_ | ~new_n8148_));
  assign new_n8163_ = new_n8164_ ? (new_n8165_ ^ new_n8171_) : (~new_n8165_ ^ new_n8171_);
  assign new_n8164_ = (~new_n8126_ & ~new_n8144_) | (new_n8125_ & (~new_n8126_ | ~new_n8144_));
  assign new_n8165_ = new_n8166_ ? (~new_n8167_ ^ new_n8168_) : (new_n8167_ ^ new_n8168_);
  assign new_n8166_ = (~new_n8131_ & new_n8130_) | (~new_n8127_ & (~new_n8131_ | new_n8130_));
  assign new_n8167_ = new_n8128_ & new_n8129_;
  assign new_n8168_ = new_n8169_ ^ new_n8170_;
  assign new_n8169_ = (~new_n8142_ & ~new_n8143_) | (new_n8132_ & (~new_n8142_ | ~new_n8143_));
  assign new_n8170_ = (new_n8140_ & new_n8141_) | (new_n8133_ & (new_n8140_ | new_n8141_));
  assign new_n8171_ = new_n8172_ ? (new_n8173_ ^ new_n8174_) : (~new_n8173_ ^ new_n8174_);
  assign new_n8172_ = (new_n8146_ & new_n8147_) | (new_n8145_ & (new_n8146_ | new_n8147_));
  assign new_n8173_ = ~new_n8152_ & new_n8151_;
  assign new_n8174_ = new_n8153_ & new_n8154_;
  assign new_n8175_ = (~new_n8150_ & new_n8155_) | (new_n8149_ & (~new_n8150_ | new_n8155_));
  assign \o[53]  = ~new_n8177_ ^ new_n8178_;
  assign new_n8177_ = (new_n8160_ | (~new_n8161_ & (new_n8159_ | new_n8158_))) & (new_n8159_ | new_n8158_ | ~new_n8161_);
  assign new_n8178_ = new_n8179_ ^ new_n8180_;
  assign new_n8179_ = (~new_n8163_ & new_n8175_) | (new_n8162_ & (~new_n8163_ | new_n8175_));
  assign new_n8180_ = new_n8181_ ? (~new_n8182_ ^ new_n8185_) : (new_n8182_ ^ new_n8185_);
  assign new_n8181_ = (~new_n8165_ & ~new_n8171_) | (new_n8164_ & (~new_n8165_ | ~new_n8171_));
  assign new_n8182_ = ~new_n8183_ ^ new_n8184_;
  assign new_n8183_ = (~new_n8168_ & new_n8167_) | (new_n8166_ & (~new_n8168_ | new_n8167_));
  assign new_n8184_ = ~new_n8169_ & new_n8170_;
  assign new_n8185_ = (new_n8173_ & new_n8174_) | (new_n8172_ & (new_n8173_ | new_n8174_));
  assign \o[54]  = ((new_n8187_ | new_n8188_) & (~new_n8189_ ^ new_n8190_)) | (~new_n8187_ & ~new_n8188_ & (~new_n8189_ ^ ~new_n8190_));
  assign new_n8187_ = ~new_n8178_ & new_n8177_;
  assign new_n8188_ = ~new_n8180_ & new_n8179_;
  assign new_n8189_ = (~new_n8182_ & new_n8185_) | (new_n8181_ & (~new_n8182_ | new_n8185_));
  assign new_n8190_ = new_n8183_ & new_n8184_;
  assign \o[55]  = (new_n8190_ | new_n8187_ | new_n8188_) & (new_n8189_ | (new_n8190_ & (new_n8187_ | new_n8188_)));
  assign \o[56]  = new_n8193_ ^ new_n8551_;
  assign new_n8193_ = new_n8194_ ? (~new_n8483_ ^ new_n8537_) : (new_n8483_ ^ new_n8537_);
  assign new_n8194_ = new_n8195_ ? (~new_n8307_ ^ new_n8471_) : (new_n8307_ ^ new_n8471_);
  assign new_n8195_ = new_n8196_ ? (~new_n8284_ ^ new_n8295_) : (new_n8284_ ^ new_n8295_);
  assign new_n8196_ = new_n8197_ ? (~new_n8241_ ^ new_n8272_) : (new_n8241_ ^ new_n8272_);
  assign new_n8197_ = new_n8198_ ? (~new_n8213_ ^ new_n8227_) : (new_n8213_ ^ new_n8227_);
  assign new_n8198_ = new_n3342_ ? (~new_n8209_ & (new_n8210_ | new_n8212_ | ~new_n6683_)) : new_n8199_;
  assign new_n8199_ = new_n8208_ ? new_n8200_ : (new_n8203_ | (~\i[743]  & new_n3744_ & new_n8206_));
  assign new_n8200_ = new_n3756_ ? ((~\i[1721]  & new_n4521_) ? new_n7785_ : new_n8202_) : new_n8201_;
  assign new_n8201_ = new_n3395_ ? new_n4470_ : (\i[1967]  & (\i[1964]  | \i[1965]  | \i[1966] ));
  assign new_n8202_ = ~\i[2623]  & (~\i[2622]  | (~\i[2621]  & ~\i[2620] ));
  assign new_n8203_ = ~new_n3744_ & (new_n8204_ ? (\i[1439]  | (\i[1437]  & \i[1438] )) : new_n8205_);
  assign new_n8204_ = ~\i[1199]  & (~\i[1197]  | ~\i[1198]  | ~\i[1196] );
  assign new_n8205_ = ~\i[2747]  & (~\i[2745]  | ~\i[2746]  | ~\i[2744] );
  assign new_n8206_ = (\i[743]  | ~new_n8207_ | ~\i[742] ) & (\i[2723]  | (\i[2722]  & \i[2721] ));
  assign new_n8207_ = \i[740]  & \i[741] ;
  assign new_n8208_ = \i[1087]  & \i[1086]  & \i[1084]  & \i[1085] ;
  assign new_n8209_ = ~new_n6683_ & ((~new_n3373_ & ~new_n4315_) | (new_n6839_ & new_n4315_ & (\i[2389]  | ~new_n3264_)));
  assign new_n8210_ = new_n8211_ & new_n4781_ & (\i[1083]  | (\i[1081]  & \i[1082] ));
  assign new_n8211_ = ~\i[1395]  & (~\i[1393]  | ~\i[1394]  | ~\i[1392] );
  assign new_n8212_ = ~\i[1083]  & (~\i[1081]  | ~\i[1082] ) & (~\i[1367]  | (~\i[1365]  & ~\i[1366] ));
  assign new_n8213_ = (new_n8214_ & (\i[2286]  | \i[2287] )) | (~\i[2286]  & ~\i[2287]  & (new_n3263_ ? ~new_n8224_ : ~new_n8220_));
  assign new_n8214_ = new_n8219_ ? (new_n8218_ | (~\i[1167]  & new_n4880_ & new_n5703_)) : new_n8215_;
  assign new_n8215_ = (\i[1950]  & \i[1951] ) ? new_n8216_ : (new_n8217_ | (~new_n4764_ & \i[2507] ));
  assign new_n8216_ = new_n5589_ ? new_n4353_ : new_n6470_;
  assign new_n8217_ = \i[2279]  & \i[2278]  & new_n4764_ & \i[2277] ;
  assign new_n8218_ = new_n6219_ & \i[1167]  & (~new_n3287_ | (~\i[2056]  & ~\i[2057] ));
  assign new_n8219_ = \i[2743]  & (\i[2741]  | \i[2742]  | \i[2740] );
  assign new_n8220_ = (~new_n8223_ | (new_n8221_ ? new_n8222_ : ~new_n3233_)) & (new_n5063_ | ~new_n3324_ | new_n8223_);
  assign new_n8221_ = ~\i[2047]  & (~\i[2046]  | (~\i[2045]  & ~\i[2044] ));
  assign new_n8222_ = \i[2054]  & \i[2055]  & (\i[2053]  | \i[2052] );
  assign new_n8223_ = \i[2515]  & \i[2514]  & \i[2512]  & \i[2513] ;
  assign new_n8224_ = (new_n8225_ | (\i[818]  & \i[819] )) & (new_n3574_ | new_n8226_ | \i[1375]  | ~\i[818]  | ~\i[819] );
  assign new_n8225_ = ~new_n3634_ & (\i[2271]  | (\i[2268]  & \i[2269]  & \i[2270] ));
  assign new_n8226_ = \i[1372]  & \i[1374]  & ~\i[1375]  & \i[1373] ;
  assign new_n8227_ = (new_n8235_ | new_n8232_ | ~new_n4821_) & (new_n4821_ | (~new_n8228_ & (new_n8239_ | new_n4199_)));
  assign new_n8228_ = new_n4199_ & (new_n8231_ ? new_n8229_ : (~new_n5651_ | ~new_n4779_));
  assign new_n8229_ = (\i[2527]  | new_n8230_ | ~new_n4990_) & (~\i[2399]  | new_n4990_ | (~\i[2398]  & ~\i[2397] ));
  assign new_n8230_ = \i[2526]  & (\i[2525]  | \i[2524] );
  assign new_n8231_ = ~\i[2643]  & (~\i[2642]  | ~\i[2641] );
  assign new_n8232_ = new_n4880_ & (new_n3421_ ? (~\i[2391]  | ~\i[2390] ) : new_n8233_);
  assign new_n8233_ = (\i[2075]  | ~new_n8234_) & (~\i[2742]  | ~\i[2743]  | new_n8234_ | (~\i[2741]  & ~\i[2740] ));
  assign new_n8234_ = \i[1947]  & (\i[1946]  | (\i[1945]  & \i[1944] ));
  assign new_n8235_ = new_n8236_ & ((~new_n8238_ & ~\i[1857]  & ~\i[1858]  & ~\i[1859] ) | (~new_n8237_ & (\i[1857]  | \i[1858]  | \i[1859] )));
  assign new_n8236_ = ~new_n4880_ & ~\i[1851]  & (~\i[1850]  | ~\i[1849] );
  assign new_n8237_ = ~\i[2299]  & ~\i[2297]  & ~\i[2298] ;
  assign new_n8238_ = \i[1527]  & \i[1526]  & \i[1524]  & \i[1525] ;
  assign new_n8239_ = new_n3288_ ? ((\i[2494]  | \i[2495] ) & (\i[2395]  | \i[2394] )) : new_n8240_;
  assign new_n8240_ = ~new_n3339_ & (~\i[2615]  | (~\i[2612]  & ~\i[2613]  & ~\i[2614] ));
  assign new_n8241_ = new_n8242_ ? (~new_n8254_ ^ new_n8264_) : (new_n8254_ ^ new_n8264_);
  assign new_n8242_ = new_n3618_ ? new_n8243_ : ((~new_n8251_ & ~new_n8253_ & new_n4048_) | (~new_n8248_ & ~new_n4048_));
  assign new_n8243_ = ~new_n8244_ & (~new_n8246_ | (new_n7464_ & (new_n4362_ ? ~\i[1271]  : new_n3376_)));
  assign new_n8244_ = ~new_n8245_ & ~new_n3682_ & new_n6770_ & (~\i[2075]  | ~\i[2074]  | ~\i[2073] );
  assign new_n8245_ = new_n7464_ & (\i[1837]  | \i[1836] );
  assign new_n8246_ = ~new_n6770_ & (~new_n8247_ | (\i[1930]  & \i[1931]  & (\i[1929]  | \i[1928] )));
  assign new_n8247_ = ~new_n7464_ & ~\i[1851]  & (~\i[1850]  | (~\i[1848]  & ~\i[1849] ));
  assign new_n8248_ = (new_n8249_ | ~new_n8250_) & (~new_n3683_ | ~new_n5052_ | new_n8250_);
  assign new_n8249_ = (\i[617]  | \i[618]  | \i[619]  | ~new_n3777_) & (~new_n3234_ | new_n3777_);
  assign new_n8250_ = \i[1067]  & (\i[1065]  | \i[1066]  | \i[1064] );
  assign new_n8251_ = ~\i[1731]  & new_n8252_ & (~\i[1730]  | ~\i[1729] );
  assign new_n8252_ = \i[1627]  & \i[2631]  & (\i[2630]  | (\i[2628]  & \i[2629] ));
  assign new_n8253_ = ~new_n4057_ & ~\i[2110]  & ~\i[2111]  & (\i[1731]  | (\i[1729]  & \i[1730] ));
  assign new_n8254_ = new_n4821_ ? (new_n3528_ ? ~new_n8263_ : ~new_n8262_) : new_n8255_;
  assign new_n8255_ = ~new_n8256_ & ((~\i[1954]  & ~\i[1955] ) | (~new_n8261_ & (new_n3322_ | new_n8259_)));
  assign new_n8256_ = ~new_n8257_ & ~\i[1954]  & ~\i[1955]  & (~new_n6770_ | new_n6729_ | ~new_n8245_);
  assign new_n8257_ = ~new_n6770_ & (new_n8258_ ? (~\i[1947]  | (~\i[1945]  & ~\i[1946] )) : new_n3372_);
  assign new_n8258_ = ~\i[819]  & (~\i[818]  | (~\i[817]  & ~\i[816] ));
  assign new_n8259_ = (\i[1431]  & (\i[1429]  | \i[1430] )) ? new_n8260_ : ~\i[987] ;
  assign new_n8260_ = \i[1606]  & \i[1607]  & (\i[1605]  | \i[1604] );
  assign new_n8261_ = new_n3322_ & (new_n4136_ ? (~new_n4396_ | (~\i[952]  & ~\i[953] )) : new_n5094_);
  assign new_n8262_ = (new_n7032_ | ~new_n5586_) & (new_n4220_ | ~new_n4171_ | new_n5586_);
  assign new_n8263_ = new_n3230_ ? ((new_n6168_ | ~new_n6172_) & (~\i[1294]  | ~\i[1295]  | new_n6172_)) : ~new_n4039_;
  assign new_n8264_ = (new_n8270_ & ~new_n7071_) | (~new_n8267_ & ~new_n8265_ & new_n7071_);
  assign new_n8265_ = new_n8266_ & (new_n3502_ | ~new_n3365_ | (\i[2539]  & (\i[2537]  | \i[2538] )));
  assign new_n8266_ = ~new_n3299_ & (~new_n3502_ | (\i[1735]  & (\i[1965]  | \i[1966]  | \i[1967] )));
  assign new_n8267_ = new_n3299_ & ((~\i[2283]  & (~\i[2281]  | ~\i[2282] )) ? ~new_n8269_ : ~new_n8268_);
  assign new_n8268_ = (~\i[2407]  & (~\i[2406]  | (~\i[2404]  & ~\i[2405] ))) ? new_n5048_ : ~new_n4069_;
  assign new_n8269_ = new_n4331_ ? (~\i[647]  & (~\i[644]  | ~\i[645]  | ~\i[646] )) : ~new_n3395_;
  assign new_n8270_ = (new_n4804_ | new_n8271_ | new_n3791_) & (new_n3898_ | ~new_n3608_ | ~new_n3791_);
  assign new_n8271_ = \i[1491]  & \i[1490]  & \i[1488]  & \i[1489] ;
  assign new_n8272_ = (new_n8273_ | new_n8276_ | ~new_n5543_) & (new_n5543_ | (~new_n8280_ & (new_n8281_ | ~new_n8283_)));
  assign new_n8273_ = new_n4667_ & ~new_n8274_ & ~\i[1283] ;
  assign new_n8274_ = (~new_n8275_ & ~new_n4850_) | (\i[1071]  & new_n4850_ & (\i[1070]  | \i[1069] ));
  assign new_n8275_ = \i[1274]  & \i[1275]  & (\i[1273]  | \i[1272] );
  assign new_n8276_ = ~new_n4667_ & (new_n8279_ ? (new_n3993_ ? new_n7307_ : new_n4071_) : ~new_n8277_);
  assign new_n8277_ = new_n3619_ ? ~new_n8278_ : ~new_n5422_;
  assign new_n8278_ = ~\i[1103]  & ~\i[1101]  & ~\i[1102] ;
  assign new_n8279_ = \i[615]  & (\i[614]  | \i[613] );
  assign new_n8280_ = new_n4080_ & ((~new_n3233_ & ~new_n3544_) | (new_n4066_ & new_n4950_ & new_n3544_));
  assign new_n8281_ = ~new_n8282_ & ~\i[2279]  & new_n3363_ & (~\i[2278]  | ~\i[2277]  | ~\i[2276] );
  assign new_n8282_ = \i[1282]  & \i[1283]  & (\i[1281]  | \i[1280] );
  assign new_n8283_ = ~new_n4080_ & ((~new_n4407_ & \i[2731] ) | ~new_n8282_ | ~new_n4100_);
  assign new_n8284_ = new_n6742_ ? (new_n3369_ ? new_n8289_ : new_n8291_) : new_n8285_;
  assign new_n8285_ = (new_n4939_ | new_n7227_ | ~new_n8288_) & (new_n8288_ | (new_n4424_ ? new_n8286_ : new_n8287_));
  assign new_n8286_ = (new_n6062_ | ~new_n7016_) & (\i[2596]  | \i[2597]  | \i[2598]  | \i[2599]  | new_n7016_);
  assign new_n8287_ = (new_n3258_ & ~new_n5567_) | (~\i[1959]  & new_n5567_ & (~\i[1958]  | ~\i[1957] ));
  assign new_n8288_ = \i[1139]  & (\i[1138]  | \i[1137] );
  assign new_n8289_ = (new_n3556_ & ~\i[1297] ) ? new_n8290_ : (new_n5725_ | (~\i[1837]  & new_n3994_));
  assign new_n8290_ = (new_n3448_ | (new_n6101_ & (~\i[724]  | ~\i[725] ))) & (~\i[607]  | ~\i[606]  | ~new_n6101_ | (\i[724]  & \i[725] ));
  assign new_n8291_ = (~new_n5077_ & new_n8294_ & new_n6336_) | (~new_n6336_ & (new_n8293_ | new_n8292_));
  assign new_n8292_ = ~\i[1275]  & (new_n3720_ | \i[1183] ) & (~\i[1274]  | (~\i[1272]  & ~\i[1273] ));
  assign new_n8293_ = ~new_n3720_ & ~\i[1183]  & ~\i[1498]  & ~\i[1499]  & (~\i[1497]  | ~\i[1496] );
  assign new_n8294_ = ~\i[1103]  & (~\i[1101]  | ~\i[1102]  | ~\i[1100] );
  assign new_n8295_ = (new_n8302_ | new_n8305_ | new_n5516_) & (~new_n5516_ | (~new_n8296_ & (~new_n8301_ | new_n8300_)));
  assign new_n8296_ = ~\i[2263]  & ~\i[2262]  & ~\i[2261]  & ~\i[2260]  & ~new_n8297_ & ~new_n8299_;
  assign new_n8297_ = new_n8298_ & ((~\i[2433]  & ~\i[2432] ) | \i[2435]  | ~\i[2434] );
  assign new_n8298_ = \i[1831]  & \i[1830]  & ~\i[2435]  & ~\i[2267]  & ~\i[2265]  & ~\i[2266] ;
  assign new_n8299_ = (~\i[1831]  | ~\i[1830] ) & (~new_n7464_ | ~\i[1836]  | ~\i[1837] );
  assign new_n8300_ = new_n4355_ & \i[1995]  & (\i[1994]  | \i[1993]  | \i[1992] );
  assign new_n8301_ = new_n5842_ & (\i[2260]  | \i[2261]  | \i[2262]  | \i[2263] );
  assign new_n8302_ = new_n4968_ & ((~new_n4662_ & ~new_n8303_ & new_n8304_) | (~new_n3985_ & new_n4520_ & ~new_n8304_));
  assign new_n8303_ = \i[2739]  & (\i[2738]  | (\i[2737]  & \i[2736] ));
  assign new_n8304_ = ~\i[2158]  & ~\i[2159]  & (~\i[2157]  | ~\i[2156] );
  assign new_n8305_ = ~new_n4968_ & new_n8306_ & (\i[1954]  | \i[1953]  | \i[1952] );
  assign new_n8306_ = \i[2179]  & \i[2178]  & \i[1955]  & \i[1262]  & \i[1263] ;
  assign new_n8307_ = new_n8308_ ? (~new_n8374_ ^ new_n8459_) : (new_n8374_ ^ new_n8459_);
  assign new_n8308_ = new_n8309_ ? (~new_n8351_ ^ new_n8364_) : (new_n8351_ ^ new_n8364_);
  assign new_n8309_ = new_n8310_ ? (~new_n8326_ ^ new_n8337_) : (new_n8326_ ^ new_n8337_);
  assign new_n8310_ = (new_n8314_ | new_n8311_ | new_n3795_) & (new_n8321_ | ~new_n3795_ | (new_n8325_ & ~new_n8317_));
  assign new_n8311_ = ~new_n8313_ & ((~new_n8312_ & new_n7442_) | (~new_n6956_ & \i[2291]  & ~new_n7442_));
  assign new_n8312_ = (\i[2521]  | \i[2522]  | \i[2523]  | ~new_n5148_) & (~new_n4109_ | new_n5148_);
  assign new_n8313_ = \i[2519]  & \i[2518]  & \i[2516]  & \i[2517] ;
  assign new_n8314_ = new_n8313_ & ((~new_n4980_ & new_n3704_ & ~new_n3314_) | (new_n3314_ & (new_n8316_ | new_n8315_)));
  assign new_n8315_ = ~new_n4414_ & (~\i[1747]  | (~\i[1746]  & (~\i[1745]  | ~\i[1744] )));
  assign new_n8316_ = new_n4414_ & \i[2411]  & (\i[2410]  | (\i[2408]  & \i[2409] ));
  assign new_n8317_ = (~new_n6956_ | new_n6726_ | new_n8320_) & (~new_n8320_ | (new_n8318_ ? new_n8319_ : ~new_n7483_));
  assign new_n8318_ = ~\i[2295]  & (~\i[2293]  | ~\i[2294]  | ~\i[2292] );
  assign new_n8319_ = \i[2654]  & \i[2655] ;
  assign new_n8320_ = ~\i[2615]  & (~\i[2614]  | (~\i[2613]  & ~\i[2612] ));
  assign new_n8321_ = ~new_n8325_ & ((~\i[2409]  & new_n4674_) ? new_n8322_ : new_n8323_);
  assign new_n8322_ = (~new_n3469_ & \i[2426]  & \i[2427]  & (\i[2424]  | \i[2425] )) | (~new_n4186_ & (~\i[2426]  | ~\i[2427]  | (~\i[2424]  & ~\i[2425] )));
  assign new_n8323_ = (~new_n5102_ & ~new_n8324_) | (\i[2325]  & \i[2326]  & \i[2327]  & new_n8324_);
  assign new_n8324_ = ~\i[1651]  & ~\i[1649]  & ~\i[1650] ;
  assign new_n8325_ = ~\i[2538]  & ~\i[2539]  & (~\i[2537]  | ~\i[2536] );
  assign new_n8326_ = (new_n8334_ | new_n8327_ | ~\i[1159] ) & (\i[1159]  | (new_n8336_ ? ~new_n8331_ : ~new_n8333_));
  assign new_n8327_ = ~\i[1395]  & (new_n8328_ | (~new_n8329_ & ~new_n8330_));
  assign new_n8328_ = ~new_n3366_ & new_n8329_ & \i[2415]  & (\i[2414]  | \i[2413]  | \i[2412] );
  assign new_n8329_ = new_n3269_ & ~\i[1608]  & ~\i[1609] ;
  assign new_n8330_ = ~\i[1958]  & ~\i[1959]  & (~\i[1957]  | ~\i[1956] );
  assign new_n8331_ = (~new_n8332_ | (~\i[1499]  & (~\i[1497]  | ~\i[1498] ))) & (new_n4094_ | new_n7744_ | \i[1499]  | (\i[1497]  & \i[1498] ));
  assign new_n8332_ = (~\i[1993]  | ~\i[1994]  | ~\i[1995] ) & (~new_n5810_ | (\i[1145]  & \i[1144] ));
  assign new_n8333_ = (new_n5612_ | new_n8211_ | new_n6791_) & (new_n3795_ | new_n7762_ | ~new_n6791_);
  assign new_n8334_ = \i[1395]  & (new_n5744_ ? new_n8335_ : (~new_n7806_ | (~\i[2626]  & ~\i[2627] )));
  assign new_n8335_ = \i[1623]  & (~\i[1055]  | (~\i[1054]  & ~\i[1053] ));
  assign new_n8336_ = \i[1391]  & \i[1389]  & \i[1390] ;
  assign new_n8337_ = (new_n8344_ | new_n8348_ | new_n4440_) & (~new_n4440_ | (new_n8350_ ? new_n8341_ : new_n8338_));
  assign new_n8338_ = (~\i[2506]  & ~\i[2507]  & (new_n8340_ | new_n8339_)) | (~new_n4434_ & new_n3993_ & (\i[2506]  | \i[2507] ));
  assign new_n8339_ = (~\i[2515]  | ~\i[2514] ) & (~\i[2615]  | (~\i[2614]  & ~\i[2613] ));
  assign new_n8340_ = \i[2615]  & (\i[2382]  | \i[2383]  | \i[2381] ) & (\i[2613]  | \i[2614] );
  assign new_n8341_ = ~new_n8342_ & (new_n7320_ | ~new_n5156_ | ~\i[767]  | (~\i[766]  & ~\i[765] ));
  assign new_n8342_ = ~new_n5156_ & (new_n8343_ ? (\i[1263]  | \i[1262] ) : new_n6287_);
  assign new_n8343_ = ~\i[2415]  & (~\i[2414]  | (~\i[2413]  & ~\i[2412] ));
  assign new_n8344_ = new_n3376_ & (new_n3905_ ? new_n8345_ : (new_n5494_ ? new_n3644_ : ~new_n8347_));
  assign new_n8345_ = (new_n8346_ | new_n4426_) & (~\i[2494]  | ~\i[2495]  | ~new_n4426_);
  assign new_n8346_ = \i[1047]  & (\i[1045]  | \i[1046]  | \i[1044] );
  assign new_n8347_ = ~\i[527]  & (~\i[525]  | ~\i[526]  | ~\i[524] );
  assign new_n8348_ = ~new_n3376_ & ~new_n8349_ & (\i[1755]  | \i[1754] );
  assign new_n8349_ = (~new_n6138_ & new_n3451_) | (~\i[1972]  & ~\i[1973]  & ~\i[1974]  & ~\i[1975]  & ~new_n3451_);
  assign new_n8350_ = \i[1303]  & \i[1302]  & \i[1300]  & \i[1301] ;
  assign new_n8351_ = (new_n8352_ | ~new_n8362_) & (new_n8361_ | ~new_n8363_ | new_n8362_);
  assign new_n8352_ = (new_n8353_ & ~new_n8360_) | (~new_n8357_ & new_n8360_ & (~new_n8359_ | ~new_n8355_));
  assign new_n8353_ = (new_n4168_ | new_n3376_ | new_n3775_) & (~new_n3775_ | (new_n4727_ ? new_n5263_ : new_n8354_));
  assign new_n8354_ = ~\i[843]  & (~\i[842]  | ~\i[841] );
  assign new_n8355_ = ~new_n8356_ & (~\i[2866]  | (~\i[2864]  & ~\i[2865] ));
  assign new_n8356_ = \i[2639]  & \i[2637]  & \i[2638] ;
  assign new_n8357_ = new_n8356_ & (new_n3442_ | new_n8358_) & (~\i[1069]  | ~\i[1070]  | ~\i[1071]  | ~new_n8358_);
  assign new_n8358_ = \i[2187]  & (\i[2185]  | \i[2186]  | \i[2184] );
  assign new_n8359_ = ~\i[2867]  & (~\i[2505]  | ~\i[2506]  | ~\i[2507]  | ~\i[2504] );
  assign new_n8360_ = \i[2643]  & (\i[2641]  | \i[2642]  | \i[2640] );
  assign new_n8361_ = (new_n3828_ & ~new_n7429_) | (~new_n5529_ & new_n6237_ & new_n7429_);
  assign new_n8362_ = ~\i[1211]  & (~\i[1210]  | (~\i[1209]  & ~\i[1208] ));
  assign new_n8363_ = ~\i[2823]  & ~\i[2821]  & ~\i[2822] ;
  assign new_n8364_ = ~new_n8365_ & (~new_n8372_ | (~new_n8369_ & ~new_n4491_));
  assign new_n8365_ = ~new_n4194_ & (new_n8366_ | ~new_n7381_) & (\i[1407]  | ~new_n6232_ | ~new_n4087_ | new_n7381_);
  assign new_n8366_ = (new_n8367_ | ~new_n5019_) & (~new_n8368_ | new_n5019_ | (\i[1043]  & (\i[1042]  | ~new_n3225_)));
  assign new_n8367_ = new_n5387_ ? ~new_n5738_ : (\i[2267]  | (\i[2265]  & \i[2266] ));
  assign new_n8368_ = ~\i[1075]  & ~\i[1073]  & ~\i[1074] ;
  assign new_n8369_ = (~new_n8370_ | new_n8371_) & (new_n5063_ | ~new_n3534_ | ~new_n8371_);
  assign new_n8370_ = new_n7893_ & (~\i[2396]  | ~\i[2397]  | ~\i[2398]  | ~\i[2399] );
  assign new_n8371_ = ~\i[1639]  & (~\i[1637]  | ~\i[1638]  | ~\i[1636] );
  assign new_n8372_ = new_n4194_ & (~new_n8373_ | ((~new_n4930_ | new_n8211_) & (~\i[2422]  | ~\i[2423]  | ~new_n8211_)));
  assign new_n8373_ = new_n4491_ & (~\i[507]  | (~\i[505]  & ~\i[506] ));
  assign new_n8374_ = new_n8375_ ? (~new_n8420_ ^ new_n8429_) : (new_n8420_ ^ new_n8429_);
  assign new_n8375_ = new_n8376_ ? (~new_n8391_ ^ new_n8407_) : (new_n8391_ ^ new_n8407_);
  assign new_n8376_ = new_n6673_ ? (new_n8384_ | (~new_n8389_ & new_n3889_ & new_n6306_)) : new_n8377_;
  assign new_n8377_ = (new_n8378_ | new_n4049_) & (new_n8380_ | new_n8383_ | ~new_n4049_);
  assign new_n8378_ = new_n3760_ ? new_n8379_ : (new_n5957_ | (\i[1597]  & \i[1598]  & \i[1599] ));
  assign new_n8379_ = (\i[2083]  | (\i[2082]  & \i[2081] )) & (\i[1867]  | \i[1866] );
  assign new_n8380_ = new_n3564_ & (new_n4067_ ? new_n8382_ : (~\i[1267]  | new_n8381_));
  assign new_n8381_ = ~\i[1266]  & (~\i[1265]  | ~\i[1264] );
  assign new_n8382_ = \i[2531]  & \i[2529]  & \i[2530] ;
  assign new_n8383_ = \i[1603]  & \i[1602]  & \i[1601]  & ~new_n6065_ & ~new_n3564_;
  assign new_n8384_ = ~new_n3889_ & (new_n7781_ ? ~new_n8388_ : new_n8385_);
  assign new_n8385_ = (~new_n8387_ & new_n8386_) | (\i[2406]  & \i[2407]  & ~new_n8386_);
  assign new_n8386_ = ~\i[2179]  & (~\i[2177]  | ~\i[2178]  | ~\i[2176] );
  assign new_n8387_ = \i[1834]  & \i[1835]  & (\i[1833]  | \i[1832] );
  assign new_n8388_ = new_n4759_ & \i[2623]  & (\i[2622]  | (\i[2620]  & \i[2621] ));
  assign new_n8389_ = (~new_n3454_ | new_n8390_) & (~\i[2181]  | ~\i[2182]  | ~\i[2183]  | ~new_n8390_);
  assign new_n8390_ = \i[1515]  & (\i[1514]  | (\i[1513]  & \i[1512] ));
  assign new_n8391_ = new_n7071_ ? new_n8392_ : ((~new_n8403_ & ~new_n8406_ & new_n5913_) | (new_n8399_ & ~new_n5913_));
  assign new_n8392_ = (new_n8395_ | new_n8397_ | new_n4132_) & (new_n8393_ | new_n8394_ | ~new_n4132_);
  assign new_n8393_ = new_n5636_ & (new_n6724_ ? ~new_n5704_ : new_n6762_);
  assign new_n8394_ = ~new_n5636_ & (new_n7722_ | new_n3587_) & (~\i[2489]  | ~\i[2490]  | ~\i[2491]  | ~new_n3587_);
  assign new_n8395_ = new_n8396_ & new_n4757_ & new_n4961_;
  assign new_n8396_ = \i[843]  & \i[841]  & \i[842] ;
  assign new_n8397_ = ~new_n8396_ & new_n4235_ & new_n8398_ & (~\i[1285]  | ~\i[1284] );
  assign new_n8398_ = ~\i[1503]  & (~\i[1501]  | ~\i[1502]  | ~\i[1500] );
  assign new_n8399_ = (new_n8400_ | new_n8401_ | new_n4277_) & (new_n8402_ | ~\i[1635]  | ~new_n4277_);
  assign new_n8400_ = ~new_n6289_ & ((~\i[1521]  & ~\i[1520] ) | ~\i[1523]  | ~\i[1522] );
  assign new_n8401_ = new_n6289_ & (~\i[833]  | ~\i[834]  | ~\i[835] );
  assign new_n8402_ = ~\i[2527]  & (~\i[2526]  | ~\i[2525] );
  assign new_n8403_ = ~new_n8405_ & (new_n4109_ ? new_n5606_ : (~\i[2599]  | new_n8404_));
  assign new_n8404_ = ~\i[2598]  & (~\i[2597]  | ~\i[2596] );
  assign new_n8405_ = ~\i[2271]  & (~\i[2270]  | ~\i[2269] );
  assign new_n8406_ = new_n8405_ & (new_n4209_ ? new_n3281_ : (~\i[1607]  | ~\i[1606] ));
  assign new_n8407_ = new_n4673_ ? (~new_n8415_ & (new_n6429_ | new_n8417_ | ~new_n8418_)) : new_n8408_;
  assign new_n8408_ = new_n8413_ ? new_n8409_ : ((new_n8412_ | new_n5617_) & (new_n8414_ | ~\i[1291]  | ~new_n5617_));
  assign new_n8409_ = new_n3663_ ? new_n8410_ : (new_n4382_ | (~\i[730]  & ~\i[731] ));
  assign new_n8410_ = (new_n4998_ | ~new_n8411_) & (~\i[1329]  | ~\i[1330]  | ~\i[1331]  | new_n8411_);
  assign new_n8411_ = \i[615]  & (\i[613]  | \i[614]  | \i[612] );
  assign new_n8412_ = ~new_n6902_ & (~\i[1533]  | ~\i[1534]  | ~\i[1535] );
  assign new_n8413_ = \i[2087]  & (\i[2086]  | \i[2085] );
  assign new_n8414_ = \i[1439]  & (\i[1437]  | \i[1438]  | \i[1436] );
  assign new_n8415_ = new_n8417_ & (new_n7751_ ? new_n8416_ : (~new_n4968_ | ~new_n4693_));
  assign new_n8416_ = \i[1211]  & (~\i[1731]  | ~\i[1730] );
  assign new_n8417_ = ~\i[1154]  & ~\i[1155]  & (~\i[1153]  | ~\i[1152] );
  assign new_n8418_ = new_n8419_ ? (\i[2503]  & (\i[2500]  | \i[2501]  | \i[2502] )) : ~new_n3240_;
  assign new_n8419_ = ~\i[1607]  & (~\i[1606]  | (~\i[1605]  & ~\i[1604] ));
  assign new_n8420_ = (new_n8421_ & ~new_n3376_) | (~new_n8425_ & new_n3376_ & (new_n5077_ | new_n8427_));
  assign new_n8421_ = new_n6973_ ? ((new_n8424_ | new_n5237_) & (new_n7442_ | ~new_n8303_ | ~new_n5237_)) : new_n8422_;
  assign new_n8422_ = (new_n8423_ & ~new_n5460_) | (~new_n5957_ & new_n5460_ & (~\i[2531]  | ~\i[2530] ));
  assign new_n8423_ = new_n7756_ ? new_n3756_ : new_n7336_;
  assign new_n8424_ = ~new_n3497_ & (~new_n4330_ | ~\i[1496]  | ~\i[1497] );
  assign new_n8425_ = new_n8426_ & (new_n7309_ | \i[931]  | ~new_n7001_ | (\i[930]  & \i[929] ));
  assign new_n8426_ = new_n5077_ & (new_n7001_ | (~new_n3383_ & ~\i[2417]  & ~\i[2418]  & ~\i[2419] ));
  assign new_n8427_ = ~new_n8428_ & (~new_n7743_ | ~\i[2424]  | ~\i[2425]  | ~\i[2426]  | ~\i[2427] );
  assign new_n8428_ = ~new_n7743_ & (new_n4657_ ? (~new_n4286_ | (\i[2520]  & \i[2521] )) : ~new_n3363_);
  assign new_n8429_ = new_n8430_ ? (~new_n8441_ ^ new_n8451_) : (new_n8441_ ^ new_n8451_);
  assign new_n8430_ = (new_n3219_ | (~new_n8438_ & (new_n8440_ | new_n8431_))) & (new_n8434_ | new_n8436_ | ~new_n3219_);
  assign new_n8431_ = (new_n6931_ | ~new_n8433_ | new_n6885_) & (new_n8432_ | ~new_n6885_ | (new_n7071_ & new_n3762_));
  assign new_n8432_ = ~new_n7071_ & ~\i[1599]  & (~\i[1598]  | ~\i[1597]  | ~\i[1596] );
  assign new_n8433_ = \i[883]  & \i[881]  & \i[882] ;
  assign new_n8434_ = new_n3233_ & ((new_n5083_ & ~new_n7756_) | (~new_n7437_ & ~new_n8435_ & new_n7756_));
  assign new_n8435_ = \i[1723]  & (\i[1722]  | (\i[1721]  & \i[1720] ));
  assign new_n8436_ = ~new_n3233_ & (new_n6670_ ? (new_n4162_ ? ~new_n6072_ : ~new_n3781_) : ~new_n8437_);
  assign new_n8437_ = \i[1195]  & new_n3988_ & \i[1194] ;
  assign new_n8438_ = new_n8440_ & (new_n8439_ | ~new_n3672_ | new_n7755_) & (new_n3242_ | new_n6519_ | ~new_n7755_);
  assign new_n8439_ = ~\i[2631]  & (~\i[2630]  | (~\i[2629]  & ~\i[2628] ));
  assign new_n8440_ = ~\i[2087]  & ~\i[2085]  & ~\i[2086] ;
  assign new_n8441_ = new_n3462_ ? ((new_n8442_ | new_n8450_ | ~new_n7401_) & (new_n8444_ | new_n7401_)) : new_n8445_;
  assign new_n8442_ = new_n4891_ ? ~new_n8443_ : (\i[1631]  | (\i[1629]  & \i[1630] ));
  assign new_n8443_ = \i[2515]  & ~new_n3776_ & \i[2514] ;
  assign new_n8444_ = (new_n3587_ | ~new_n4084_ | ~new_n7516_) & (new_n7293_ | ~new_n5383_ | new_n7516_);
  assign new_n8445_ = (new_n8447_ | new_n4336_) & (new_n8446_ | new_n4693_ | ~new_n4336_);
  assign new_n8446_ = (~new_n3645_ | new_n4804_) & (~\i[1717]  | ~\i[1718]  | ~\i[1719]  | ~new_n4804_);
  assign new_n8447_ = (new_n3893_ | new_n8449_ | ~new_n8448_) & (~new_n3730_ | ~new_n3890_ | new_n8448_);
  assign new_n8448_ = ~\i[1947]  & (~\i[1946]  | (~\i[1945]  & ~\i[1944] ));
  assign new_n8449_ = ~\i[2278]  & ~\i[2279]  & (~\i[2277]  | ~\i[2276] );
  assign new_n8450_ = ~\i[2387]  & (~\i[2385]  | ~\i[2386]  | ~\i[2384] );
  assign new_n8451_ = (~new_n8456_ & ~new_n8457_ & new_n8458_) | (~new_n8458_ & (new_n5316_ ? new_n8452_ : new_n8453_));
  assign new_n8452_ = (new_n3323_ | ~new_n8435_ | new_n4247_) & (new_n5067_ | ~new_n4247_ | (~\i[1955]  & ~\i[1954] ));
  assign new_n8453_ = new_n3715_ ? new_n8454_ : ((new_n8455_ & new_n4389_) | (\i[2402]  & \i[2403]  & ~new_n4389_));
  assign new_n8454_ = new_n6863_ ? (~\i[2735]  & (~\i[2732]  | ~\i[2733]  | ~\i[2734] )) : new_n3257_;
  assign new_n8455_ = new_n3491_ & (~\i[2641]  | ~\i[2640] );
  assign new_n8456_ = new_n3467_ & ((~new_n4209_ & new_n4725_ & new_n5435_) | (~new_n5847_ & new_n3716_ & ~new_n5435_));
  assign new_n8457_ = ~new_n3467_ & (~new_n6708_ | ~new_n6833_ | ~new_n3997_) & (new_n5383_ | new_n4659_ | new_n3997_);
  assign new_n8458_ = \i[1622]  & \i[1623]  & (\i[1621]  | \i[1620] );
  assign new_n8459_ = new_n3448_ ? new_n8460_ : ((new_n8465_ | ~new_n8245_) & (new_n8468_ | new_n8470_ | new_n8245_));
  assign new_n8460_ = new_n4804_ ? new_n8461_ : (new_n8463_ | (~new_n3264_ & ~new_n4785_ & \i[2175] ));
  assign new_n8461_ = new_n3405_ ? (new_n5455_ ? ~new_n5428_ : new_n5616_) : new_n8462_;
  assign new_n8462_ = (new_n7783_ | ~new_n4074_) & (~\i[1951]  | new_n4074_ | (~\i[1950]  & (~\i[1948]  | ~\i[1949] )));
  assign new_n8463_ = new_n8464_ & (\i[1499]  | (\i[1498]  & (\i[1497]  | \i[1496] )));
  assign new_n8464_ = ~\i[2439]  & new_n3264_ & (~\i[2438]  | (~\i[2436]  & ~\i[2437] ));
  assign new_n8465_ = new_n3834_ ? (new_n8467_ ? ~new_n5589_ : ~new_n5196_) : new_n8466_;
  assign new_n8466_ = (~new_n5704_ & \i[630]  & \i[631]  & (\i[628]  | \i[629] )) | (new_n5025_ & (~\i[630]  | ~\i[631]  | (~\i[628]  & ~\i[629] )));
  assign new_n8467_ = ~\i[2270]  & ~\i[2271]  & (~\i[2269]  | ~\i[2268] );
  assign new_n8468_ = new_n8469_ & ((new_n4424_ & new_n5586_) | (~\i[2635]  & ~new_n5586_ & (~\i[2634]  | ~\i[2633] )));
  assign new_n8469_ = \i[1307]  & \i[1305]  & \i[1306] ;
  assign new_n8470_ = \i[2327]  & \i[2326]  & \i[2325]  & \i[2324]  & ~new_n4389_ & ~new_n8469_;
  assign new_n8471_ = new_n8482_ ? ((new_n8480_ | ~new_n8481_) & (~new_n8479_ | new_n8477_)) : new_n8472_;
  assign new_n8472_ = (new_n8474_ | new_n8473_ | new_n3306_) & (~new_n3306_ | (new_n8476_ ? new_n8475_ : ~new_n5036_));
  assign new_n8473_ = ~\i[1107]  & ~\i[1106]  & ~new_n4440_ & ~new_n7737_;
  assign new_n8474_ = ~new_n5148_ & ~\i[2391]  & new_n4440_ & (~\i[2390]  | (~\i[2388]  & ~\i[2389] ));
  assign new_n8475_ = (~\i[1088]  | ~\i[1089]  | ~\i[1090]  | ~\i[1091]  | new_n4093_) & (new_n4697_ | ~new_n4093_);
  assign new_n8476_ = ~\i[1615]  & (~\i[1614]  | (~\i[1613]  & ~\i[1612] ));
  assign new_n8477_ = new_n4190_ & (new_n8478_ ? ~new_n5584_ : ~new_n6539_);
  assign new_n8478_ = ~\i[927]  & (~\i[925]  | ~\i[926]  | ~\i[924] );
  assign new_n8479_ = ~new_n5577_ & (new_n3491_ | new_n4190_);
  assign new_n8480_ = new_n4428_ & \i[2607]  & (\i[2736]  | \i[2737]  | \i[2738]  | \i[2739] );
  assign new_n8481_ = new_n5577_ & (new_n4428_ | new_n6068_ | \i[2626]  | \i[2627] );
  assign new_n8482_ = ~\i[1767]  & ~\i[1766]  & ~\i[1764]  & ~\i[1765] ;
  assign new_n8483_ = new_n8484_ ? (~new_n8518_ ^ new_n8527_) : (new_n8518_ ^ new_n8527_);
  assign new_n8484_ = new_n8485_ ? (~new_n8495_ ^ new_n8507_) : (new_n8495_ ^ new_n8507_);
  assign new_n8485_ = new_n4141_ ? new_n8486_ : (new_n8382_ ? new_n8491_ : new_n8493_);
  assign new_n8486_ = (new_n4199_ | new_n4382_ | new_n4724_ | ~new_n8490_) & (new_n8487_ | new_n8490_);
  assign new_n8487_ = new_n6238_ ? (new_n4806_ ? new_n8489_ : new_n3775_) : new_n8488_;
  assign new_n8488_ = (~\i[1415]  & new_n4705_ & \i[2408]  & \i[2409] ) | (new_n4726_ & (~new_n4705_ | ~\i[2408]  | ~\i[2409] ));
  assign new_n8489_ = ~\i[2310]  & ~\i[2311]  & (~\i[2309]  | ~\i[2308] );
  assign new_n8490_ = \i[1749]  & new_n5679_ & \i[1748] ;
  assign new_n8491_ = new_n4103_ ? (new_n4437_ | (\i[946]  & \i[947] )) : new_n8492_;
  assign new_n8492_ = (~new_n4232_ | new_n4750_) & (~\i[1047]  | ~new_n4750_ | (~\i[1046]  & (~\i[1044]  | ~\i[1045] )));
  assign new_n8493_ = (\i[719]  & (\i[718]  | (\i[716]  & \i[717] ))) ? new_n8494_ : new_n4136_;
  assign new_n8494_ = \i[2531]  ? (~new_n5530_ | (~\i[1624]  & ~\i[1625] )) : new_n6257_;
  assign new_n8495_ = new_n3624_ ? ((new_n8498_ | ~new_n4979_) & (new_n8496_ | new_n8506_ | new_n4979_)) : new_n8501_;
  assign new_n8496_ = ~new_n8497_ & ~\i[2291]  & (~\i[2290]  | ~\i[2289] );
  assign new_n8497_ = (~new_n4919_ | new_n5262_) & (~\i[2325]  | ~\i[2326]  | ~\i[2327]  | ~new_n5262_);
  assign new_n8498_ = new_n4010_ ? new_n8499_ : (new_n6073_ ? new_n8500_ : new_n4985_);
  assign new_n8499_ = (~\i[2611]  | ~new_n3263_ | (~\i[2610]  & (~\i[2608]  | ~\i[2609] ))) & (new_n3423_ | new_n3263_);
  assign new_n8500_ = ~\i[1819]  & ~\i[1817]  & ~\i[1818] ;
  assign new_n8501_ = new_n3254_ ? new_n8502_ : ((~new_n8505_ & ~new_n5048_) | (~new_n4257_ & new_n7920_ & new_n5048_));
  assign new_n8502_ = new_n3711_ ? new_n8503_ : new_n8504_;
  assign new_n8503_ = (~\i[2183]  & (~\i[2182]  | (~\i[2180]  & ~\i[2181] ))) ? new_n8449_ : ~new_n7405_;
  assign new_n8504_ = (~new_n4337_ & (\i[514]  | \i[515] )) | (~\i[737]  & ~\i[738]  & ~\i[739]  & ~\i[514]  & ~\i[515] );
  assign new_n8505_ = (~new_n5025_ | new_n5108_) & (\i[1094]  | \i[1095]  | ~new_n5108_);
  assign new_n8506_ = (~\i[1287]  | ~\i[1285]  | ~\i[1286] ) & (\i[2291]  | (\i[2290]  & \i[2289] ));
  assign new_n8507_ = ~new_n8508_ & (~new_n5156_ | ((new_n8513_ | ~new_n7751_) & (new_n8516_ | new_n8517_ | new_n7751_)));
  assign new_n8508_ = new_n8511_ & (~\i[941]  | ~\i[942]  | ~\i[943]  | (~new_n8510_ & ~new_n8509_));
  assign new_n8509_ = new_n3504_ & (new_n5442_ | ~\i[1507] ) & (~\i[2645]  | ~\i[2646]  | ~\i[2647]  | \i[1507] );
  assign new_n8510_ = new_n3302_ & ~new_n3504_ & ~new_n7374_;
  assign new_n8511_ = ~new_n5156_ & (~new_n7269_ | ~new_n8512_ | ~\i[2417]  | ~\i[2418]  | ~\i[2419] );
  assign new_n8512_ = (~\i[943]  | ~\i[941]  | ~\i[942] ) & (~\i[1279]  | (~\i[1278]  & ~\i[1277] ));
  assign new_n8513_ = (~\i[2615]  & (~\i[2612]  | ~\i[2613]  | ~\i[2614] )) ? new_n8515_ : new_n8514_;
  assign new_n8514_ = ~\i[1603]  & (new_n4808_ | ~\i[1602] ) & (~\i[1843]  | new_n3940_);
  assign new_n8515_ = ~\i[1159]  & new_n3409_ & (~\i[1158]  | ~\i[1157]  | ~\i[1156] );
  assign new_n8516_ = new_n6662_ & ((~new_n5822_ & ~new_n8303_) | (~\i[631]  & new_n8303_ & (~\i[630]  | ~\i[629] )));
  assign new_n8517_ = ~new_n6662_ & new_n6724_ & \i[2182]  & \i[2183]  & (\i[2181]  | \i[2180] );
  assign new_n8518_ = new_n3373_ ? (new_n4653_ ? ~new_n8523_ : ~new_n8526_) : new_n8519_;
  assign new_n8519_ = new_n4007_ ? (new_n8522_ | (new_n8520_ & new_n7307_)) : new_n8521_;
  assign new_n8520_ = \i[1299]  & new_n6357_ & \i[1298] ;
  assign new_n8521_ = ~new_n7287_ & ~new_n4013_ & (\i[2179]  | (\i[2178]  & (\i[2177]  | \i[2176] )));
  assign new_n8522_ = ~new_n7307_ & (\i[2635]  | \i[2634]  | ~new_n4881_) & (~\i[1391]  | ~\i[1390]  | new_n4881_);
  assign new_n8523_ = (~new_n8524_ | new_n4310_) & (~new_n4194_ | ~\i[1967]  | ~new_n4310_ | (~\i[1966]  & ~\i[1965] ));
  assign new_n8524_ = ~\i[1059]  & new_n8525_ & (~\i[1058]  | ~\i[1057] );
  assign new_n8525_ = \i[2282]  & \i[2283]  & (\i[2281]  | \i[2280] );
  assign new_n8526_ = (new_n6757_ | \i[1643]  | new_n3221_) & (~new_n3221_ | (new_n5678_ ? new_n6263_ : ~new_n4985_));
  assign new_n8527_ = new_n8536_ ? (new_n8530_ | (~new_n8528_ & ~new_n8534_ & new_n4285_)) : new_n8531_;
  assign new_n8528_ = new_n8529_ & ((new_n4936_ & ~new_n8450_) | (\i[2301]  & \i[2302]  & \i[2303]  & new_n8450_));
  assign new_n8529_ = ~\i[2742]  & ~\i[2743]  & (~\i[2741]  | ~\i[2740] );
  assign new_n8530_ = ~new_n5720_ & ~new_n5513_ & ~new_n4285_ & ~new_n3634_;
  assign new_n8531_ = (~new_n7006_ & ~\i[847]  & new_n7351_ & new_n4134_) | (~new_n4134_ & (new_n8533_ | new_n8532_));
  assign new_n8532_ = ~new_n4794_ & new_n3691_ & (~\i[1715]  | ~\i[1714]  | ~\i[1713] );
  assign new_n8533_ = new_n5742_ & new_n4794_ & (~\i[1407]  | (~\i[1404]  & ~\i[1405]  & ~\i[1406] ));
  assign new_n8534_ = ~new_n8529_ & ~new_n8535_ & (\i[1943]  | ~\i[1610]  | ~\i[1611]  | ~\i[1609] );
  assign new_n8535_ = \i[1943]  & (\i[2279]  | (\i[2277]  & \i[2278] ));
  assign new_n8536_ = ~\i[995]  & ~\i[994]  & ~\i[992]  & ~\i[993] ;
  assign new_n8537_ = new_n8550_ ? new_n8538_ : (new_n8546_ ? new_n8547_ : new_n8545_);
  assign new_n8538_ = ~new_n8539_ & (new_n7032_ | (new_n8543_ & new_n8544_) | (~new_n8541_ & ~new_n8544_));
  assign new_n8539_ = new_n7032_ & (new_n7370_ ? (new_n5717_ ? ~new_n5810_ : ~new_n4428_) : ~new_n8540_);
  assign new_n8540_ = new_n5494_ & new_n3459_ & ~\i[2176]  & ~\i[2177] ;
  assign new_n8541_ = ~new_n8542_ & (new_n5837_ | (\i[2746]  & \i[2747] ));
  assign new_n8542_ = new_n5837_ & ~\i[2831]  & ~\i[2829]  & ~\i[2830] ;
  assign new_n8543_ = ~new_n5685_ & ~\i[2526]  & ~\i[2527]  & (~\i[2525]  | ~\i[2524] );
  assign new_n8544_ = \i[1199]  & (\i[1198]  | (\i[1197]  & \i[1196] ));
  assign new_n8545_ = (new_n4973_ | ~new_n5070_ | ~new_n7364_) & (new_n8411_ | ~\i[967]  | new_n7364_);
  assign new_n8546_ = new_n7473_ & ~\i[2436]  & ~\i[2437] ;
  assign new_n8547_ = (~new_n8549_ | new_n8548_) & (new_n4330_ | new_n3618_ | ~new_n8548_);
  assign new_n8548_ = \i[1331]  & (\i[1330]  | \i[1329] );
  assign new_n8549_ = ~\i[1767]  & ~\i[1978]  & ~\i[1979]  & (~\i[1766]  | (~\i[1765]  & ~\i[1764] ));
  assign new_n8550_ = ~\i[1762]  & ~\i[1763]  & (~\i[1761]  | ~\i[1760] );
  assign new_n8551_ = new_n4249_ ? ((new_n8560_ | new_n8562_ | ~new_n3564_) & (new_n8557_ | new_n3564_)) : new_n8552_;
  assign new_n8552_ = (new_n8553_ | new_n6656_) & (new_n8556_ | ~new_n6656_ | (new_n4056_ & (~new_n3719_ | ~\i[1287] )));
  assign new_n8553_ = new_n3995_ ? new_n8554_ : (new_n8555_ ? new_n8294_ : ~new_n4779_);
  assign new_n8554_ = new_n5101_ ? (~\i[2651]  & (~\i[2648]  | ~\i[2649]  | ~\i[2650] )) : new_n5508_;
  assign new_n8555_ = ~\i[2651]  & (~\i[2650]  | ~\i[2649] );
  assign new_n8556_ = ~new_n4056_ & (new_n4336_ ? (\i[1947]  | \i[1946] ) : ~new_n3602_);
  assign new_n8557_ = ~new_n8558_ & (~new_n4937_ | (~new_n8278_ & ~new_n8411_) | (~new_n8559_ & new_n8411_));
  assign new_n8558_ = ~new_n8336_ & ~new_n4937_ & \i[1291]  & (\i[1290]  | (\i[1288]  & \i[1289] ));
  assign new_n8559_ = ~\i[1047]  & (~\i[1046]  | (~\i[1045]  & ~\i[1044] ));
  assign new_n8560_ = ~\i[1735]  & ((~\i[1608]  & ~\i[1609] ) | ~new_n8561_ | ~new_n7353_);
  assign new_n8561_ = ~\i[1671]  & (~\i[1670]  | (~\i[1669]  & ~\i[1668] ));
  assign new_n8562_ = ~new_n3680_ & \i[1735]  & (~\i[1951]  | (~\i[1948]  & ~\i[1949]  & ~\i[1950] ));
  assign \o[57]  = new_n8564_ ^ new_n8565_;
  assign new_n8564_ = ~new_n8193_ & ~new_n8551_;
  assign new_n8565_ = new_n8566_ ? (~new_n8567_ ^ new_n8649_) : (new_n8567_ ^ new_n8649_);
  assign new_n8566_ = (~new_n8483_ & ~new_n8537_) | (~new_n8194_ & (~new_n8483_ | ~new_n8537_));
  assign new_n8567_ = new_n8568_ ? (~new_n8569_ ^ new_n8641_) : (new_n8569_ ^ new_n8641_);
  assign new_n8568_ = (~new_n8307_ & ~new_n8471_) | (~new_n8195_ & (~new_n8307_ | ~new_n8471_));
  assign new_n8569_ = new_n8570_ ? (~new_n8592_ ^ new_n8593_) : (new_n8592_ ^ new_n8593_);
  assign new_n8570_ = new_n8571_ ? (new_n8572_ ^ new_n8591_) : (~new_n8572_ ^ new_n8591_);
  assign new_n8571_ = (~new_n8241_ & ~new_n8272_) | (~new_n8197_ & (~new_n8241_ | ~new_n8272_));
  assign new_n8572_ = new_n8573_ ? (new_n8574_ ^ new_n8585_) : (~new_n8574_ ^ new_n8585_);
  assign new_n8573_ = (~new_n8213_ & ~new_n8227_) | (~new_n8198_ & (~new_n8213_ | ~new_n8227_));
  assign new_n8574_ = new_n8575_ ? (new_n8579_ ^ new_n8584_) : (~new_n8579_ ^ new_n8584_);
  assign new_n8575_ = (new_n8576_ | new_n6673_) & (new_n8578_ | new_n3889_ | ~new_n6673_);
  assign new_n8576_ = (~new_n3564_ | ~new_n4067_ | ~new_n8382_ | ~new_n4049_) & (~new_n8577_ | new_n3760_ | new_n4049_);
  assign new_n8577_ = new_n5957_ & ((~\i[2717]  & ~\i[2716] ) | ~\i[2719]  | ~\i[2718] );
  assign new_n8578_ = (~new_n8385_ | new_n7781_) & (new_n4759_ | ~new_n7781_ | (~\i[1647]  & (~\i[1645]  | ~\i[1646] )));
  assign new_n8579_ = ~new_n8581_ & (~new_n8482_ | new_n8481_ | (~new_n8477_ & ~new_n5577_ & ~new_n8580_));
  assign new_n8580_ = ~new_n4190_ & ~new_n3491_ & ~\i[2378]  & ~\i[2379]  & (~\i[2377]  | ~\i[2376] );
  assign new_n8581_ = ~new_n8482_ & new_n3306_ & ((new_n8582_ & ~new_n8476_) | (new_n4093_ & new_n4697_ & new_n8476_));
  assign new_n8582_ = ~new_n5036_ & new_n8583_;
  assign new_n8583_ = ~\i[2082]  & ~\i[2083]  & (~\i[2081]  | ~\i[2080] );
  assign new_n8584_ = (new_n8529_ | ~new_n4285_ | ~new_n8535_ | ~new_n8536_) & (~new_n8532_ | new_n4134_ | new_n8536_);
  assign new_n8585_ = new_n8586_ ? (~new_n8588_ ^ new_n8590_) : (new_n8588_ ^ new_n8590_);
  assign new_n8586_ = \i[1159]  ? new_n8587_ : (new_n8336_ ? new_n8331_ : new_n8333_);
  assign new_n8587_ = ~new_n8334_ & (new_n8329_ | new_n8330_ | \i[1395]  | (\i[599]  & \i[598] ));
  assign new_n8588_ = (new_n3369_ | new_n6336_ | ~new_n8292_ | ~new_n6742_) & (~new_n8589_ | new_n4939_ | new_n6742_);
  assign new_n8589_ = new_n7227_ & new_n8288_;
  assign new_n8590_ = new_n4440_ & new_n8340_ & ~\i[2507]  & ~new_n8350_ & ~\i[2506] ;
  assign new_n8591_ = (~new_n8351_ & ~new_n8364_) | (~new_n8309_ & (~new_n8351_ | ~new_n8364_));
  assign new_n8592_ = (~new_n8374_ & ~new_n8459_) | (~new_n8308_ & (~new_n8374_ | ~new_n8459_));
  assign new_n8593_ = new_n8594_ ? (~new_n8595_ ^ new_n8629_) : (new_n8595_ ^ new_n8629_);
  assign new_n8594_ = (~new_n8420_ & ~new_n8429_) | (~new_n8375_ & (~new_n8420_ | ~new_n8429_));
  assign new_n8595_ = new_n8596_ ? (~new_n8608_ ^ new_n8628_) : (new_n8608_ ^ new_n8628_);
  assign new_n8596_ = ~new_n8597_ ^ new_n8601_;
  assign new_n8597_ = new_n3219_ ? new_n8598_ : ((new_n8600_ | ~new_n8440_) & (~new_n8432_ | ~new_n6885_ | new_n8440_));
  assign new_n8598_ = ~new_n8436_ & (~new_n3233_ | (~new_n8599_ & (new_n4368_ | ~new_n7437_ | ~new_n7756_)));
  assign new_n8599_ = ~new_n7756_ & (~new_n5857_ | ~new_n5083_) & (~new_n3898_ | ~\i[1180]  | ~\i[1181]  | new_n5083_);
  assign new_n8600_ = (new_n6519_ | new_n3242_ | ~new_n7755_) & (new_n7755_ | (new_n3672_ ? new_n8439_ : new_n7887_));
  assign new_n8601_ = new_n8458_ ? new_n8604_ : (new_n5316_ ? new_n8602_ : new_n8607_);
  assign new_n8602_ = (new_n8603_ | ~new_n4247_) & (~new_n3323_ | ~\i[1623]  | new_n4247_ | (~\i[1622]  & ~\i[1621] ));
  assign new_n8603_ = (~\i[646]  | ~\i[647]  | ~\i[645]  | ~new_n5067_) & (new_n5067_ | (~\i[1955]  & ~\i[1954] ));
  assign new_n8604_ = (new_n3997_ | new_n4659_ | new_n3467_) & (new_n8606_ | ~new_n3467_ | (new_n4209_ & new_n8605_));
  assign new_n8605_ = new_n4725_ & new_n5435_;
  assign new_n8606_ = ~new_n5435_ & (new_n3716_ ? new_n5847_ : ~new_n3293_);
  assign new_n8607_ = (new_n6863_ | new_n3257_ | ~new_n3715_) & (new_n4389_ | ~\i[2402]  | ~\i[2403]  | new_n3715_);
  assign new_n8608_ = new_n8609_ ? (~new_n8613_ ^ new_n8623_) : (new_n8613_ ^ new_n8623_);
  assign new_n8609_ = (new_n8610_ | new_n8550_) & (new_n7032_ | new_n8544_ | ~new_n8542_ | ~new_n8550_);
  assign new_n8610_ = (new_n8611_ | new_n8546_) & (new_n3618_ | ~new_n4330_ | ~new_n8548_ | ~new_n8546_);
  assign new_n8611_ = ~new_n8612_ & (\i[1822]  | \i[1823]  | ~new_n4973_ | ~new_n7364_);
  assign new_n8612_ = ~new_n7364_ & ~\i[519]  & new_n8411_ & (~\i[518]  | ~\i[517]  | ~\i[516] );
  assign new_n8613_ = new_n3462_ ? (new_n7401_ ? new_n8619_ : new_n8622_) : new_n8614_;
  assign new_n8614_ = new_n4336_ ? new_n8616_ : ((new_n8615_ | ~new_n8448_) & (new_n3890_ | ~new_n6324_ | new_n8448_));
  assign new_n8615_ = new_n3893_ ? new_n4470_ : ~new_n8449_;
  assign new_n8616_ = (new_n3645_ | new_n4804_ | new_n4693_) & (new_n8617_ | new_n8618_ | ~new_n4693_);
  assign new_n8617_ = ~\i[1403]  & new_n3287_ & (~\i[1402]  | (~\i[1400]  & ~\i[1401] ));
  assign new_n8618_ = ~new_n3287_ & (~\i[2181]  | ~\i[2182]  | ~\i[2183] );
  assign new_n8619_ = (new_n8620_ | ~new_n8450_) & (new_n4891_ | new_n8450_ | (~\i[1631]  & (~\i[1629]  | ~\i[1630] )));
  assign new_n8620_ = (new_n8621_ | ~\i[2546]  | ~\i[2547] ) & (~\i[2858]  | ~\i[2859]  | (\i[2546]  & \i[2547] ));
  assign new_n8621_ = ~\i[2527]  & ~\i[2525]  & ~\i[2526] ;
  assign new_n8622_ = (new_n4084_ | ~new_n3737_ | ~new_n7516_) & (new_n5383_ | ~new_n5073_ | new_n7516_);
  assign new_n8623_ = ~new_n8624_ & (new_n4249_ | (~new_n8627_ & (new_n8626_ | new_n8556_ | ~new_n6656_)));
  assign new_n8624_ = new_n8625_ & (~new_n3564_ | ((new_n8561_ | \i[1735] ) & (~new_n3680_ | ~new_n5231_ | ~\i[1735] )));
  assign new_n8625_ = new_n4249_ & (new_n3564_ | ~new_n4937_ | (new_n8411_ ? new_n8559_ : new_n8278_));
  assign new_n8626_ = new_n4056_ & (\i[1287]  ? ~new_n3719_ : (\i[1495]  | (\i[1493]  & \i[1494] )));
  assign new_n8627_ = ~new_n6656_ & (~new_n5508_ | new_n5101_ | ~new_n3995_) & (new_n4779_ | new_n8555_ | new_n3995_);
  assign new_n8628_ = (~new_n8441_ & ~new_n8451_) | (~new_n8430_ & (~new_n8441_ | ~new_n8451_));
  assign new_n8629_ = new_n8630_ ? (new_n8631_ ^ new_n8632_) : (~new_n8631_ ^ new_n8632_);
  assign new_n8630_ = (~new_n8326_ & ~new_n8337_) | (~new_n8310_ & (~new_n8326_ | ~new_n8337_));
  assign new_n8631_ = (~new_n8391_ & ~new_n8407_) | (~new_n8376_ & (~new_n8391_ | ~new_n8407_));
  assign new_n8632_ = new_n8633_ ? (~new_n8637_ ^ new_n8639_) : (new_n8637_ ^ new_n8639_);
  assign new_n8633_ = (new_n8635_ | new_n8413_ | new_n4673_) & (~new_n4673_ | (new_n8417_ ? ~new_n8636_ : ~new_n8634_));
  assign new_n8634_ = new_n6429_ ? (new_n3347_ ? new_n3539_ : ~new_n8330_) : ~new_n8418_;
  assign new_n8635_ = (~new_n8412_ | new_n5617_) & (~new_n6855_ | ~new_n8414_ | ~new_n5617_);
  assign new_n8636_ = new_n7751_ & \i[1730]  & \i[1731]  & (\i[1159]  | \i[1158]  | \i[1157] );
  assign new_n8637_ = ~new_n8638_ & (new_n5636_ | new_n3587_ | ~new_n4132_ | ~new_n7071_ | ~new_n7722_);
  assign new_n8638_ = ~new_n5913_ & ~new_n7071_ & ((new_n8401_ & ~new_n4277_) | (new_n4245_ & new_n8402_ & new_n4277_));
  assign new_n8639_ = (new_n3373_ | (new_n4007_ ? ~new_n8522_ : ~new_n8521_)) & (new_n8640_ | new_n4653_ | ~new_n3373_);
  assign new_n8640_ = (new_n6757_ | \i[1643]  | new_n3221_) & (new_n5678_ | ~new_n4985_ | ~new_n3221_);
  assign new_n8641_ = new_n8642_ ? (new_n8643_ ^ new_n8648_) : (~new_n8643_ ^ new_n8648_);
  assign new_n8642_ = (~new_n8284_ & ~new_n8295_) | (~new_n8196_ & (~new_n8284_ | ~new_n8295_));
  assign new_n8643_ = (~new_n8646_ & (~new_n8644_ ^ ~new_n8645_)) | (new_n8647_ & (~new_n8644_ ^ new_n8645_));
  assign new_n8644_ = (~new_n8254_ & ~new_n8264_) | (~new_n8242_ & (~new_n8254_ | ~new_n8264_));
  assign new_n8645_ = (~new_n8305_ | new_n5516_) & (~new_n8301_ | ~new_n8300_ | ~new_n5516_);
  assign new_n8646_ = new_n5616_ & new_n4804_ & new_n3448_ & ~new_n5455_ & new_n3405_;
  assign new_n8647_ = new_n5616_ & new_n4804_ & new_n3448_ & ~new_n5455_ & new_n3405_;
  assign new_n8648_ = (~new_n8495_ & ~new_n8507_) | (~new_n8485_ & (~new_n8495_ | ~new_n8507_));
  assign new_n8649_ = (~new_n8518_ & ~new_n8527_) | (~new_n8484_ & (~new_n8518_ | ~new_n8527_));
  assign \o[58]  = ~new_n8651_ ^ new_n8652_;
  assign new_n8651_ = new_n8564_ & new_n8565_;
  assign new_n8652_ = new_n8653_ ^ new_n8654_;
  assign new_n8653_ = (new_n8567_ & new_n8649_) | (new_n8566_ & (new_n8567_ | new_n8649_));
  assign new_n8654_ = new_n8655_ ? (~new_n8656_ ^ new_n8681_) : (new_n8656_ ^ new_n8681_);
  assign new_n8655_ = (new_n8569_ & new_n8641_) | (new_n8568_ & (new_n8569_ | new_n8641_));
  assign new_n8656_ = new_n8657_ ? (new_n8661_ ^ new_n8662_) : (~new_n8661_ ^ new_n8662_);
  assign new_n8657_ = new_n8658_ ? (~new_n8659_ ^ new_n8660_) : (new_n8659_ ^ new_n8660_);
  assign new_n8658_ = (~new_n8572_ & new_n8591_) | (new_n8571_ & (~new_n8572_ | new_n8591_));
  assign new_n8659_ = (~new_n8647_ & new_n8645_) | (~new_n8644_ & (~new_n8647_ | new_n8645_));
  assign new_n8660_ = (~new_n8588_ & new_n8590_) | (~new_n8586_ & (~new_n8588_ | new_n8590_));
  assign new_n8661_ = (new_n8592_ & new_n8593_) | (new_n8570_ & (new_n8592_ | new_n8593_));
  assign new_n8662_ = new_n8663_ ? (new_n8667_ ^ new_n8668_) : (~new_n8667_ ^ new_n8668_);
  assign new_n8663_ = new_n8664_ ? (new_n8665_ ^ new_n8666_) : (~new_n8665_ ^ new_n8666_);
  assign new_n8664_ = (new_n8574_ & new_n8585_) | (new_n8573_ & (new_n8574_ | new_n8585_));
  assign new_n8665_ = (~new_n8632_ & new_n8631_) | (new_n8630_ & (~new_n8632_ | new_n8631_));
  assign new_n8666_ = (~new_n8579_ & ~new_n8584_) | (~new_n8575_ & (~new_n8579_ | ~new_n8584_));
  assign new_n8667_ = (new_n8595_ & new_n8629_) | (new_n8594_ & (new_n8595_ | new_n8629_));
  assign new_n8668_ = new_n8669_ ? (new_n8672_ ^ new_n8673_) : (~new_n8672_ ^ new_n8673_);
  assign new_n8669_ = ~new_n8670_ ^ new_n8671_;
  assign new_n8670_ = (~new_n8613_ & new_n8623_) | (~new_n8609_ & (~new_n8613_ | new_n8623_));
  assign new_n8671_ = (~new_n8637_ & ~new_n8639_) | (~new_n8633_ & (~new_n8637_ | ~new_n8639_));
  assign new_n8672_ = (new_n8608_ & new_n8628_) | (new_n8596_ & (new_n8608_ | new_n8628_));
  assign new_n8673_ = ~new_n8674_ ^ new_n8675_;
  assign new_n8674_ = new_n8597_ & new_n8601_;
  assign new_n8675_ = (new_n8676_ & (new_n4245_ | new_n5913_ | new_n7071_ | ~new_n4277_ | ~new_n8402_)) | (~new_n4245_ & ~new_n5913_ & ~new_n7071_ & new_n4277_ & new_n8402_ & ~new_n8676_);
  assign new_n8676_ = (new_n8677_ | ~new_n8458_) & (new_n5316_ | new_n4389_ | ~new_n8680_ | new_n8458_);
  assign new_n8677_ = (new_n8678_ | new_n3467_) & (new_n3442_ | new_n4725_ | ~new_n5435_ | ~new_n3467_);
  assign new_n8678_ = (new_n6708_ | new_n8679_ | ~new_n3997_) & (new_n3997_ | (new_n4659_ ? new_n4160_ : new_n5383_));
  assign new_n8679_ = ~\i[2623]  & ~\i[2621]  & ~\i[2622] ;
  assign new_n8680_ = ~new_n3715_ & (~\i[2403]  | ~\i[2402] );
  assign new_n8681_ = (~new_n8643_ & new_n8648_) | (new_n8642_ & (~new_n8643_ | new_n8648_));
  assign \o[59]  = ((new_n8683_ | new_n8684_) & (~new_n8685_ ^ new_n8686_)) | (~new_n8683_ & ~new_n8684_ & (~new_n8685_ ^ ~new_n8686_));
  assign new_n8683_ = ~new_n8652_ & new_n8651_;
  assign new_n8684_ = ~new_n8654_ & new_n8653_;
  assign new_n8685_ = (~new_n8656_ & new_n8681_) | (new_n8655_ & (~new_n8656_ | new_n8681_));
  assign new_n8686_ = new_n8687_ ? (new_n8688_ ^ new_n8697_) : (~new_n8688_ ^ new_n8697_);
  assign new_n8687_ = (~new_n8662_ & new_n8661_) | (~new_n8657_ & (~new_n8662_ | new_n8661_));
  assign new_n8688_ = new_n8689_ ? (~new_n8690_ ^ new_n8696_) : (new_n8690_ ^ new_n8696_);
  assign new_n8689_ = (~new_n8668_ & new_n8667_) | (~new_n8663_ & (~new_n8668_ | new_n8667_));
  assign new_n8690_ = new_n8691_ ? (~new_n8692_ ^ new_n8695_) : (new_n8692_ ^ new_n8695_);
  assign new_n8691_ = (~new_n8673_ & new_n8672_) | (~new_n8669_ & (~new_n8673_ | new_n8672_));
  assign new_n8692_ = new_n8693_ ^ new_n8694_;
  assign new_n8693_ = ~new_n8674_ & ~new_n8675_;
  assign new_n8694_ = new_n8402_ & new_n4277_ & ~new_n7071_ & ~new_n5913_ & ~new_n8676_ & ~new_n4245_;
  assign new_n8695_ = new_n8670_ & new_n8671_;
  assign new_n8696_ = (new_n8665_ & new_n8666_) | (new_n8664_ & (new_n8665_ | new_n8666_));
  assign new_n8697_ = (~new_n8659_ & new_n8660_) | (new_n8658_ & (~new_n8659_ | new_n8660_));
  assign \o[60]  = ~new_n8699_ ^ new_n8700_;
  assign new_n8699_ = (new_n8686_ | new_n8683_ | new_n8684_) & (new_n8685_ | (new_n8686_ & (new_n8683_ | new_n8684_)));
  assign new_n8700_ = new_n8701_ ^ new_n8702_;
  assign new_n8701_ = (~new_n8688_ & new_n8697_) | (new_n8687_ & (~new_n8688_ | new_n8697_));
  assign new_n8702_ = ~new_n8703_ ^ new_n8704_;
  assign new_n8703_ = (~new_n8690_ & new_n8696_) | (new_n8689_ & (~new_n8690_ | new_n8696_));
  assign new_n8704_ = ~new_n8705_ ^ new_n8706_;
  assign new_n8705_ = (~new_n8692_ & new_n8695_) | (new_n8691_ & (~new_n8692_ | new_n8695_));
  assign new_n8706_ = ~new_n8693_ & ~new_n8694_;
  assign \o[61]  = ((new_n8708_ | new_n8709_) & (~new_n8710_ ^ new_n8711_)) | (~new_n8708_ & ~new_n8709_ & (~new_n8710_ ^ ~new_n8711_));
  assign new_n8708_ = ~new_n8700_ & new_n8699_;
  assign new_n8709_ = ~new_n8702_ & new_n8701_;
  assign new_n8710_ = new_n8703_ & new_n8704_;
  assign new_n8711_ = ~new_n8706_ & new_n8705_;
  assign \o[62]  = (new_n8711_ | new_n8708_ | new_n8709_) & (new_n8710_ | (new_n8711_ & (new_n8708_ | new_n8709_)));
  assign \o[63]  = new_n8714_ ? (new_n9007_ ^ new_n9016_) : (~new_n9007_ ^ new_n9016_);
  assign new_n8714_ = new_n8715_ ? (~new_n8987_ ^ new_n8997_) : (new_n8987_ ^ new_n8997_);
  assign new_n8715_ = new_n8716_ ? (~new_n8912_ ^ new_n8985_) : (new_n8912_ ^ new_n8985_);
  assign new_n8716_ = new_n8717_ ? (~new_n8796_ ^ new_n8901_) : (new_n8796_ ^ new_n8901_);
  assign new_n8717_ = new_n8718_ ? (~new_n8782_ ^ new_n8790_) : (new_n8782_ ^ new_n8790_);
  assign new_n8718_ = new_n8719_ ? (~new_n8745_ ^ new_n8772_) : (new_n8745_ ^ new_n8772_);
  assign new_n8719_ = new_n8720_ ? (~new_n8728_ ^ new_n8739_) : (new_n8728_ ^ new_n8739_);
  assign new_n8720_ = new_n7454_ ? ((~new_n3305_ & new_n8727_) | (~new_n5550_ & new_n8726_ & ~new_n8727_)) : new_n8721_;
  assign new_n8721_ = new_n5532_ ? new_n8722_ : new_n8724_;
  assign new_n8722_ = new_n3452_ ? (new_n4317_ ? new_n4412_ : ~new_n4192_) : new_n8723_;
  assign new_n8723_ = new_n5138_ ? new_n6429_ : new_n3538_;
  assign new_n8724_ = (~new_n4891_ & (~\i[1757]  | ~\i[1758]  | ~\i[1759] )) | (new_n8725_ & \i[1757]  & \i[1758]  & \i[1759] );
  assign new_n8725_ = new_n5730_ & (~\i[613]  | ~\i[614]  | ~\i[615] );
  assign new_n8726_ = new_n3392_ & ~\i[2491]  & ~\i[2489]  & ~\i[2490] ;
  assign new_n8727_ = \i[1538]  & \i[1539]  & (\i[1537]  | \i[1536] );
  assign new_n8728_ = new_n7925_ ? new_n8729_ : (~new_n8735_ & (new_n4697_ | ~new_n8737_ | ~new_n8738_));
  assign new_n8729_ = new_n8734_ ? (new_n5479_ ? ~new_n8733_ : ~new_n8732_) : new_n8730_;
  assign new_n8730_ = new_n4895_ ? new_n4520_ : ((new_n7751_ | ~new_n5665_) & (new_n8731_ | \i[1183]  | new_n5665_));
  assign new_n8731_ = \i[1182]  & (\i[1181]  | \i[1180] );
  assign new_n8732_ = (new_n3562_ & \i[1536]  & \i[1537]  & \i[1538]  & \i[1539] ) | (\i[1639]  & (~\i[1536]  | ~\i[1537]  | ~\i[1538]  | ~\i[1539] ));
  assign new_n8733_ = ~new_n4050_ & ((~\i[2401]  & ~\i[2400] ) | ~\i[2403]  | ~\i[2402] );
  assign new_n8734_ = ~\i[2959]  & ~\i[2957]  & ~\i[2958] ;
  assign new_n8735_ = ~new_n8737_ & ((~\i[825]  & new_n4120_ & (~new_n5742_ | ~new_n5316_)) | (new_n8736_ & (\i[825]  | ~new_n4120_)));
  assign new_n8736_ = new_n5673_ & (~\i[1977]  | ~\i[1978]  | ~\i[1979] );
  assign new_n8737_ = ~\i[2307]  & (~\i[2305]  | ~\i[2306]  | ~\i[2304] );
  assign new_n8738_ = \i[847]  & (\i[846]  | (\i[845]  & \i[844] ));
  assign new_n8739_ = new_n4179_ ? new_n8740_ : ~\i[1655] ;
  assign new_n8740_ = (~new_n8743_ & ~new_n8744_ & new_n8742_) | (~new_n8742_ & (~new_n7785_ | new_n8741_));
  assign new_n8741_ = new_n6127_ & ~\i[731]  & ~\i[729]  & ~\i[730] ;
  assign new_n8742_ = \i[609]  & new_n4690_ & \i[608] ;
  assign new_n8743_ = ~new_n3759_ & (~new_n8222_ | new_n3615_) & (~\i[613]  | ~\i[614]  | ~\i[615]  | ~new_n3615_);
  assign new_n8744_ = new_n6762_ & new_n3759_ & (\i[1263]  | (\i[1260]  & \i[1261]  & \i[1262] ));
  assign new_n8745_ = new_n8746_ ? (new_n8756_ ^ new_n8763_) : (~new_n8756_ ^ new_n8763_);
  assign new_n8746_ = (new_n8747_ & ~new_n8734_) | (~new_n8752_ & new_n8734_ & (new_n8754_ | ~new_n8749_));
  assign new_n8747_ = (~new_n8748_ | ~new_n5930_) & (~\i[935]  | new_n5930_ | (\i[847]  & (\i[845]  | \i[846] )));
  assign new_n8748_ = \i[2739]  & \i[2738]  & \i[2737]  & new_n4168_ & \i[2736] ;
  assign new_n8749_ = ~new_n5387_ & ((~new_n8751_ & new_n4833_) | new_n7031_ | new_n8750_);
  assign new_n8750_ = \i[2843]  & ~new_n4833_ & \i[2842] ;
  assign new_n8751_ = \i[1759]  & \i[1758]  & \i[1756]  & \i[1757] ;
  assign new_n8752_ = ~new_n8753_ & ~new_n4950_ & ~\i[1643]  & new_n5387_ & (~\i[1642]  | ~\i[1641] );
  assign new_n8753_ = ~\i[2731]  & (~\i[2730]  | (~\i[2729]  & ~\i[2728] ));
  assign new_n8754_ = new_n7031_ & (new_n8755_ ? (~\i[2063]  | (~\i[2061]  & ~\i[2062] )) : ~new_n4950_);
  assign new_n8755_ = ~\i[1643]  & (~\i[1642]  | (~\i[1641]  & ~\i[1640] ));
  assign new_n8756_ = (new_n8762_ | ~\i[1475] ) & (new_n8761_ | new_n8757_ | \i[1475] );
  assign new_n8757_ = (~\i[2983]  | (~\i[2981]  & ~\i[2982] )) & (new_n3290_ ? new_n8758_ : new_n8759_);
  assign new_n8758_ = (~new_n3227_ | new_n3350_) & (~\i[2838]  | ~\i[2839]  | ~new_n3350_ | (~\i[2837]  & ~\i[2836] ));
  assign new_n8759_ = (\i[1541]  | \i[1542]  | \i[1543]  | ~new_n8760_) & (new_n5654_ | new_n8760_);
  assign new_n8760_ = ~\i[1986]  & ~\i[1987]  & (~\i[1985]  | ~\i[1984] );
  assign new_n8761_ = ~new_n3539_ & new_n3993_ & \i[2983]  & (\i[2982]  | \i[2981] );
  assign new_n8762_ = (new_n7812_ & new_n5522_ & new_n5558_) | (~new_n5558_ & (~\i[1059]  | ~\i[1058] ));
  assign new_n8763_ = (~\i[599]  & (~\i[598]  | (~\i[596]  & ~\i[597] ))) ? new_n8768_ : new_n8764_;
  assign new_n8764_ = (new_n8765_ | new_n8767_) & (~new_n4342_ | ~\i[840]  | ~\i[841]  | ~new_n8767_);
  assign new_n8765_ = new_n8766_ & (~\i[2732]  | ~\i[2733]  | ~\i[2734]  | ~\i[2735] );
  assign new_n8766_ = ~\i[511]  & (~\i[509]  | ~\i[510]  | ~\i[508] );
  assign new_n8767_ = \i[2663]  & (\i[2662]  | (\i[2661]  & \i[2660] ));
  assign new_n8768_ = (new_n8771_ | ~\i[2274]  | ~\i[2275] ) & (new_n8770_ | new_n8769_ | (\i[2274]  & \i[2275] ));
  assign new_n8769_ = \i[955]  & new_n3249_ & ~new_n7920_ & new_n3631_;
  assign new_n8770_ = new_n7920_ & (\i[747]  ? ~new_n6406_ : (\i[2299]  | (\i[2297]  & \i[2298] )));
  assign new_n8771_ = (~new_n7348_ | ~new_n3348_) & (~new_n6519_ | ~\i[1493]  | ~\i[1494]  | ~\i[1495]  | new_n3348_);
  assign new_n8772_ = new_n5098_ ? new_n8773_ : (new_n8781_ ? ~new_n8780_ : new_n8778_);
  assign new_n8773_ = new_n6119_ ? new_n8774_ : (~new_n8777_ & (new_n4094_ | ~new_n5654_ | ~new_n6417_));
  assign new_n8774_ = (~new_n8775_ | new_n5408_) & (\i[2533]  | \i[2534]  | \i[2535]  | ~new_n8776_ | ~new_n5408_);
  assign new_n8775_ = new_n4245_ & ~\i[1615]  & ~\i[1613]  & ~\i[1614] ;
  assign new_n8776_ = \i[1163]  & (\i[1161]  | \i[1162]  | \i[1160] );
  assign new_n8777_ = new_n4190_ & ~new_n6417_ & new_n3564_;
  assign new_n8778_ = (new_n8779_ | new_n3236_) & (~new_n3777_ | ~new_n4954_ | ~new_n3236_);
  assign new_n8779_ = (new_n5605_ & \i[2763]  & (\i[2761]  | \i[2762] )) | (\i[1854]  & \i[1855]  & (~\i[2763]  | (~\i[2761]  & ~\i[2762] )));
  assign new_n8780_ = new_n4915_ ? ((~new_n3289_ | new_n4471_) & (~\i[1254]  | ~\i[1255]  | ~new_n4471_)) : \i[2567] ;
  assign new_n8781_ = \i[1755]  & (\i[1753]  | \i[1754]  | \i[1752] );
  assign new_n8782_ = (~new_n8753_ | new_n8783_ | ~new_n8789_) & (new_n8784_ | new_n8789_ | (~new_n8788_ & new_n8787_));
  assign new_n8783_ = ~\i[1715]  & new_n5148_ & (~\i[1659]  | (~\i[1656]  & ~\i[1657]  & ~\i[1658] ));
  assign new_n8784_ = new_n8786_ & (new_n4430_ ? (new_n5684_ ? new_n5646_ : ~\i[723] ) : new_n8785_);
  assign new_n8785_ = \i[2057]  & \i[2056]  & ~new_n3609_ & new_n3287_;
  assign new_n8786_ = \i[1378]  & \i[1379]  & (\i[1377]  | \i[1376] );
  assign new_n8787_ = ~new_n8786_ & (\i[2095]  | (\i[2093]  & \i[2094] ));
  assign new_n8788_ = (~new_n7993_ | ~new_n4792_) & (new_n4153_ | \i[2430]  | \i[2431]  | new_n4792_);
  assign new_n8789_ = \i[1479]  & \i[1477]  & \i[1478] ;
  assign new_n8790_ = ~new_n8791_ & (~new_n4179_ | (~new_n8795_ & (new_n4865_ | ~new_n8793_ | ~new_n5134_)));
  assign new_n8791_ = \i[2079]  & \i[2078]  & \i[2077]  & \i[2076]  & ~new_n4179_ & new_n8792_;
  assign new_n8792_ = \i[2643]  & \i[2642]  & \i[2640]  & \i[2641] ;
  assign new_n8793_ = ~new_n8794_ & (~\i[2556]  | ~\i[2557]  | ~\i[2558]  | ~\i[2559] );
  assign new_n8794_ = ~\i[1999]  & ~\i[1997]  & ~\i[1998] ;
  assign new_n8795_ = new_n8794_ & new_n4007_ & new_n3238_ & ~\i[1619]  & ~\i[1617]  & ~\i[1618] ;
  assign new_n8796_ = new_n8797_ ? (~new_n8866_ ^ new_n8790_) : (new_n8866_ ^ new_n8790_);
  assign new_n8797_ = new_n8798_ ? (new_n8824_ ^ new_n8865_) : (~new_n8824_ ^ new_n8865_);
  assign new_n8798_ = ~new_n8799_ ^ new_n8813_;
  assign new_n8799_ = new_n8812_ ? new_n8800_ : new_n8807_;
  assign new_n8800_ = new_n5896_ ? ((~new_n8804_ & new_n8805_) | (new_n3994_ & new_n8806_ & ~new_n8805_)) : new_n8801_;
  assign new_n8801_ = (~new_n8802_ | new_n8803_) & (~new_n4520_ | (new_n8398_ ? new_n6856_ : new_n5626_));
  assign new_n8802_ = ~new_n4520_ & (~new_n6085_ | (\i[959]  & (\i[956]  | \i[957]  | \i[958] )));
  assign new_n8803_ = ~new_n6085_ & ~\i[822]  & ~\i[823]  & (~\i[821]  | ~\i[820] );
  assign new_n8804_ = (~new_n3710_ & ~\i[2880]  & ~\i[2881]  & ~\i[2882]  & ~\i[2883] ) | (new_n4361_ & (\i[2880]  | \i[2881]  | \i[2882]  | \i[2883] ));
  assign new_n8805_ = ~\i[2843]  & ~\i[2842]  & ~\i[2840]  & ~\i[2841] ;
  assign new_n8806_ = ~\i[1623]  & ~\i[1621]  & ~\i[1622] ;
  assign new_n8807_ = new_n4215_ ? (new_n7212_ ? new_n5802_ : ~new_n8811_) : new_n8808_;
  assign new_n8808_ = (~new_n6093_ | ~new_n6296_ | ~new_n7287_) & (new_n8809_ | ~new_n8810_ | new_n7287_);
  assign new_n8809_ = ~\i[926]  & ~\i[927]  & (~\i[925]  | ~\i[924] );
  assign new_n8810_ = \i[1875]  & \i[1873]  & \i[1874] ;
  assign new_n8811_ = ~\i[1042]  & ~\i[1043]  & new_n6101_ & (~\i[1041]  | ~\i[1040] );
  assign new_n8812_ = ~\i[2871]  & ~\i[2870]  & ~\i[2868]  & ~\i[2869] ;
  assign new_n8813_ = (new_n8818_ & ~new_n5079_) | (~new_n8814_ & new_n5079_ & (new_n8823_ | ~new_n8817_));
  assign new_n8814_ = new_n5763_ & (new_n8815_ | (~new_n8816_ & (new_n4331_ ? ~new_n6155_ : ~new_n3778_)));
  assign new_n8815_ = new_n8816_ & (~new_n5397_ | ~new_n3488_) & (~\i[1473]  | ~\i[1474]  | ~\i[1475]  | new_n3488_);
  assign new_n8816_ = new_n4323_ & (~\i[1385]  | ~\i[1384] );
  assign new_n8817_ = ~new_n5763_ & (new_n6375_ | (~new_n6127_ & new_n4214_) | (~new_n4371_ & ~new_n4214_));
  assign new_n8818_ = ~new_n8819_ & (~new_n7842_ | (~new_n8822_ & new_n4134_) | (new_n8821_ & ~new_n4134_));
  assign new_n8819_ = ~new_n7842_ & new_n3414_ & (new_n4273_ ? new_n4036_ : (\i[2715]  | new_n8820_));
  assign new_n8820_ = \i[2714]  & \i[2712]  & \i[2713] ;
  assign new_n8821_ = new_n3490_ & new_n5624_ & (~\i[2849]  | ~\i[2848] );
  assign new_n8822_ = ~\i[1419]  & (~\i[1417]  | ~\i[1418]  | ~\i[1416] );
  assign new_n8823_ = new_n6375_ & ((new_n4343_ & new_n6143_) | (\i[1075]  & ~new_n6143_ & (\i[1074]  | \i[1073] )));
  assign new_n8824_ = new_n8825_ ? (~new_n8838_ ^ new_n8854_) : (new_n8838_ ^ new_n8854_);
  assign new_n8825_ = ~new_n8826_ & (new_n8832_ | (~new_n8837_ & ~\i[1831]  & new_n7442_) | (~new_n8833_ & ~new_n7442_));
  assign new_n8826_ = new_n8832_ & (new_n3509_ ? ~new_n8827_ : (new_n8828_ | (~new_n8829_ & ~\i[727] )));
  assign new_n8827_ = (~new_n7204_ | ~\i[931]  | ~new_n3593_) & (new_n3540_ | ~new_n7709_ | new_n3593_);
  assign new_n8828_ = ~new_n3584_ & ~\i[2291]  & \i[727]  & (~\i[2290]  | (~\i[2288]  & ~\i[2289] ));
  assign new_n8829_ = (~new_n8831_ & new_n8830_) | (~\i[2986]  & ~\i[2987]  & ~new_n8830_);
  assign new_n8830_ = \i[2055]  & (\i[2054]  | (\i[2053]  & \i[2052] ));
  assign new_n8831_ = ~\i[827]  & (~\i[826]  | (~\i[825]  & ~\i[824] ));
  assign new_n8832_ = ~\i[2974]  & ~\i[2975]  & (~\i[2973]  | ~\i[2972] );
  assign new_n8833_ = (new_n8834_ | ~new_n8835_) & (~new_n3445_ | ~new_n8836_ | new_n8835_);
  assign new_n8834_ = (\i[2199]  & (\i[2198]  | (\i[2196]  & \i[2197] ))) ? ~new_n3544_ : ~new_n3646_;
  assign new_n8835_ = \i[1175]  & \i[1173]  & \i[1174] ;
  assign new_n8836_ = ~\i[1290]  & ~\i[1291]  & (~\i[1289]  | ~\i[1288] );
  assign new_n8837_ = \i[1387]  & (\i[1385]  | \i[1386]  | \i[1384] );
  assign new_n8838_ = (new_n6437_ & (new_n8853_ ? ~new_n8839_ : ~new_n8843_)) | (~new_n8847_ & ~new_n8850_ & ~new_n6437_);
  assign new_n8839_ = (~new_n8840_ | ~new_n6316_) & (new_n8841_ | new_n8842_ | new_n6316_);
  assign new_n8840_ = new_n6971_ & (\i[751]  | (\i[750]  & (\i[749]  | \i[748] )));
  assign new_n8841_ = \i[1647]  & (\i[1645]  | \i[1646]  | \i[1644] ) & (\i[861]  | ~new_n3504_);
  assign new_n8842_ = new_n8396_ & ~\i[863]  & ~\i[861]  & ~\i[862] ;
  assign new_n8843_ = new_n8844_ ? new_n8845_ : ((new_n6539_ | ~new_n8846_) & (~\i[2754]  | ~\i[2755]  | new_n8846_));
  assign new_n8844_ = \i[1146]  & \i[1147]  & (\i[1145]  | \i[1144] );
  assign new_n8845_ = (~\i[714]  | ~\i[715] ) & (\i[2883]  | (\i[2881]  & \i[2882]  & \i[2880] ));
  assign new_n8846_ = ~\i[2879]  & ~\i[2878]  & ~\i[2876]  & ~\i[2877] ;
  assign new_n8847_ = new_n3754_ & ~new_n8849_ & new_n8848_;
  assign new_n8848_ = \i[1267]  & \i[1266]  & \i[1264]  & \i[1265] ;
  assign new_n8849_ = \i[1871]  & \i[1870]  & \i[1868]  & \i[1869] ;
  assign new_n8850_ = ~new_n8848_ & (new_n8851_ | (new_n8852_ & (\i[1054]  | (\i[1052]  & \i[1053] ))));
  assign new_n8851_ = \i[995]  & (\i[993]  | \i[994]  | \i[992] );
  assign new_n8852_ = \i[499]  & \i[1055]  & (\i[498]  | \i[497] );
  assign new_n8853_ = ~\i[703]  & ~\i[702]  & ~\i[700]  & ~\i[701] ;
  assign new_n8854_ = ~new_n8863_ & (~new_n4179_ | (~new_n8855_ & (new_n3290_ | new_n8860_)));
  assign new_n8855_ = new_n3290_ & (new_n3220_ ? new_n8856_ : (new_n8859_ ? new_n3535_ : new_n5238_));
  assign new_n8856_ = (~new_n8858_ | ~new_n8857_) & (\i[1514]  | \i[1515]  | new_n8857_);
  assign new_n8857_ = ~\i[1643]  & (~\i[1641]  | ~\i[1642]  | ~\i[1640] );
  assign new_n8858_ = ~\i[1763]  & (~\i[1762]  | (~\i[1761]  & ~\i[1760] ));
  assign new_n8859_ = ~\i[2666]  & ~\i[2667]  & (~\i[2665]  | ~\i[2664] );
  assign new_n8860_ = new_n4077_ ? (new_n5913_ ? new_n3583_ : ~new_n5742_) : new_n8861_;
  assign new_n8861_ = (new_n8862_ | ~new_n8467_) & (~\i[1266]  | ~\i[1267]  | new_n8467_);
  assign new_n8862_ = \i[711]  & (\i[710]  | (\i[709]  & \i[708] ));
  assign new_n8863_ = ~new_n4179_ & new_n3506_ & new_n8864_ & (\i[1986]  | \i[1985]  | \i[1984] );
  assign new_n8864_ = \i[2647]  & \i[2646]  & \i[2645]  & \i[1987]  & \i[2644] ;
  assign new_n8865_ = new_n4412_ & new_n5532_ & new_n4317_ & ~new_n7454_ & new_n3452_;
  assign new_n8866_ = new_n8867_ ? (new_n8894_ ^ new_n8865_) : (~new_n8894_ ^ new_n8865_);
  assign new_n8867_ = new_n8868_ ? (new_n8877_ ^ new_n8889_) : (~new_n8877_ ^ new_n8889_);
  assign new_n8868_ = new_n8789_ ? (new_n3793_ | (~new_n8876_ & ~new_n8875_)) : new_n8869_;
  assign new_n8869_ = (new_n8874_ | new_n5080_ | \i[987]  | (\i[985]  & \i[986] )) & (new_n8870_ | (~\i[987]  & (~\i[985]  | ~\i[986] )));
  assign new_n8870_ = ~new_n8872_ & (~new_n8871_ | (\i[1655]  & (\i[1654]  | (\i[1652]  & \i[1653] ))));
  assign new_n8871_ = ~new_n6132_ & \i[838]  & \i[839]  & (\i[837]  | \i[836] );
  assign new_n8872_ = (new_n8873_ | ~\i[995]  | (\i[758]  & \i[759] )) & new_n6132_ & (~new_n3726_ | ~\i[758]  | ~\i[759] );
  assign new_n8873_ = ~\i[994]  & (~\i[993]  | ~\i[992] );
  assign new_n8874_ = ~\i[2835]  & ~\i[2834]  & ~new_n3744_ & ~\i[2833] ;
  assign new_n8875_ = new_n3400_ & new_n6798_ & (\i[1920]  | \i[1921]  | \i[1922]  | \i[1923] );
  assign new_n8876_ = ~new_n6798_ & ~\i[2882]  & ~\i[2883]  & (~\i[2555]  | (~\i[2553]  & ~\i[2554] ));
  assign new_n8877_ = ~new_n8878_ & (new_n3843_ | (~new_n8886_ & (new_n8888_ | (\i[1258]  & \i[1259] ))));
  assign new_n8878_ = new_n3843_ & (new_n4377_ ? (new_n8884_ ? ~new_n8885_ : ~new_n8883_) : new_n8879_);
  assign new_n8879_ = ~new_n8880_ & ((~\i[1665]  & ~\i[1666]  & ~\i[1667] ) | new_n7239_ | ~new_n4424_);
  assign new_n8880_ = ~\i[1667]  & ~\i[1666]  & ~\i[1665]  & ~new_n8881_ & ~new_n8882_;
  assign new_n8881_ = ~\i[2775]  & (~\i[2774]  | (~\i[2773]  & ~\i[2772] ));
  assign new_n8882_ = \i[1031]  & (\i[1029]  | \i[1030]  | \i[1028] );
  assign new_n8883_ = new_n6266_ ? new_n3351_ : ~new_n7421_;
  assign new_n8884_ = ~\i[2731]  & (~\i[2730]  | ~\i[2729] );
  assign new_n8885_ = \i[2719]  & \i[2718]  & \i[2717]  & \i[1319]  & \i[2716] ;
  assign new_n8886_ = \i[1258]  & \i[1259]  & (new_n6828_ ? new_n8884_ : (new_n8887_ | ~new_n4160_));
  assign new_n8887_ = \i[1603]  & (\i[1602]  | \i[1601] );
  assign new_n8888_ = new_n3366_ & \i[2866]  & \i[2867]  & (\i[2865]  | \i[2864] );
  assign new_n8889_ = (new_n8792_ | new_n8893_ | new_n4179_) & (new_n8890_ | ~new_n4179_ | (new_n8794_ & ~new_n8891_));
  assign new_n8890_ = new_n8793_ & (~new_n4865_ | (~\i[2447]  & (~\i[2446]  | ~\i[2445] )));
  assign new_n8891_ = (~new_n4186_ | ~new_n4323_ | new_n3238_) & (~new_n3238_ | (new_n8892_ ? ~new_n4007_ : \i[1375] ));
  assign new_n8892_ = ~\i[1619]  & ~\i[1617]  & ~\i[1618] ;
  assign new_n8893_ = ~\i[1435]  & (~\i[1433]  | ~\i[1434]  | ~\i[1432] );
  assign new_n8894_ = (new_n8895_ | ~new_n8794_) & (~\i[1429]  | ~\i[1430]  | ~\i[1431]  | new_n8794_);
  assign new_n8895_ = new_n4338_ ? (new_n7565_ ? new_n8899_ : new_n8900_) : new_n8896_;
  assign new_n8896_ = (new_n8897_ & \i[1422]  & \i[1423]  & (\i[1420]  | \i[1421] )) | (~new_n8898_ & (~\i[1422]  | ~\i[1423]  | (~\i[1420]  & ~\i[1421] )));
  assign new_n8897_ = (new_n6132_ | ~new_n6713_) & (\i[1541]  | \i[1542]  | \i[1543]  | new_n6713_);
  assign new_n8898_ = ~new_n5408_ & (~\i[1077]  | ~\i[1078]  | ~\i[1079] );
  assign new_n8899_ = (~\i[963]  & ~\i[962]  & new_n4186_) | (~new_n4186_ & (~\i[2723]  | ~\i[2722] ));
  assign new_n8900_ = (\i[2743]  | new_n5796_) & (~\i[2860]  | ~\i[2861]  | ~\i[2862]  | ~\i[2863]  | ~new_n5796_);
  assign new_n8901_ = new_n7925_ ? ((~new_n8911_ & ~new_n7933_) | (~new_n8908_ & \i[2987]  & new_n7933_)) : new_n8902_;
  assign new_n8902_ = new_n8907_ ? new_n8903_ : ((~new_n8906_ & new_n8738_) | (~new_n7421_ & ~new_n6332_ & ~new_n8738_));
  assign new_n8903_ = (new_n8904_ & ~new_n8905_) | (~new_n3368_ & new_n8905_ & (~\i[2749]  | ~new_n4803_));
  assign new_n8904_ = new_n3445_ ? new_n5773_ : new_n4356_;
  assign new_n8905_ = ~\i[967]  & (~\i[966]  | (~\i[965]  & ~\i[964] ));
  assign new_n8906_ = (~new_n3557_ & new_n4080_) | (new_n4049_ & ~new_n4080_ & (\i[1081]  | \i[1080] ));
  assign new_n8907_ = \i[2307]  & (\i[2306]  | (\i[2305]  & \i[2304] ));
  assign new_n8908_ = ~new_n8909_ & (~new_n8910_ | (\i[1751]  & (\i[1750]  | (\i[1748]  & \i[1749] ))));
  assign new_n8909_ = ~new_n8910_ & ~\i[843]  & (~\i[842]  | (~\i[840]  & ~\i[841] ));
  assign new_n8910_ = \i[1271]  & \i[1270]  & \i[1268]  & \i[1269] ;
  assign new_n8911_ = (new_n7810_ | new_n8275_ | new_n8621_) & (new_n4244_ | new_n4790_ | ~new_n8621_);
  assign new_n8912_ = new_n8913_ ? (~new_n8959_ ^ new_n8973_) : (new_n8959_ ^ new_n8973_);
  assign new_n8913_ = new_n8914_ ? (~new_n8944_ ^ new_n8953_) : (new_n8944_ ^ new_n8953_);
  assign new_n8914_ = new_n8915_ ? (~new_n8772_ ^ new_n8935_) : (new_n8772_ ^ new_n8935_);
  assign new_n8915_ = new_n8916_ ? (~new_n8922_ ^ new_n8930_) : (new_n8922_ ^ new_n8930_);
  assign new_n8916_ = ~\i[807]  & ~\i[806]  & ~new_n8917_ & ~\i[805] ;
  assign new_n8917_ = (new_n8918_ | new_n8919_ | ~\i[1371] ) & (\i[1371]  | (~new_n8920_ & (new_n8921_ | ~new_n5080_)));
  assign new_n8918_ = new_n3670_ & (~\i[1940]  | ~\i[1941] ) & (new_n5151_ ? new_n6194_ : new_n6429_);
  assign new_n8919_ = ~new_n5668_ & new_n3321_ & (~new_n3670_ | (\i[1940]  & \i[1941] ));
  assign new_n8920_ = ~new_n5080_ & new_n4919_ & ((\i[976]  & \i[977] ) | \i[979]  | \i[978] );
  assign new_n8921_ = new_n3368_ ? ~new_n6297_ : new_n5749_;
  assign new_n8922_ = (new_n8928_ | ~\i[1483]  | new_n4865_) & (new_n8923_ | ~new_n4865_ | (~new_n4694_ & ~new_n8925_));
  assign new_n8923_ = new_n4694_ & (new_n3364_ ? new_n8924_ : (new_n6357_ ? ~new_n7961_ : ~\i[2055] ));
  assign new_n8924_ = new_n6691_ ? ~new_n4379_ : ~new_n3544_;
  assign new_n8925_ = new_n8927_ ? new_n8926_ : (~new_n4028_ | (~\i[2882]  & ~\i[2883] ));
  assign new_n8926_ = (~new_n3528_ | ~new_n4949_) & (~\i[1375]  | new_n4949_ | (~\i[1374]  & (~\i[1372]  | ~\i[1373] )));
  assign new_n8927_ = \i[1299]  & \i[1297]  & \i[1298] ;
  assign new_n8928_ = (~new_n8929_ & ~new_n3637_) | (\i[1715]  & new_n3637_ & (\i[1714]  | \i[1713] ));
  assign new_n8929_ = \i[1927]  & (\i[1926]  | \i[1925] );
  assign new_n8930_ = ~new_n8931_ & (\i[598]  | \i[599]  | (~new_n8933_ & (new_n8932_ | ~new_n8467_)));
  assign new_n8931_ = new_n3521_ & (\i[598]  | \i[599] ) & (~new_n5810_ | (\i[1144]  & \i[1145] ));
  assign new_n8932_ = (~new_n3257_ | ~new_n4461_ | ~new_n3278_) & (new_n3278_ | (new_n7840_ & (~\i[2842]  | ~\i[2843] )));
  assign new_n8933_ = ~new_n8467_ & (new_n3348_ | new_n8934_) & (~\i[837]  | ~\i[838]  | ~\i[839]  | ~new_n8934_);
  assign new_n8934_ = \i[2527]  & \i[2525]  & \i[2526] ;
  assign new_n8935_ = new_n5408_ ? new_n8936_ : ((~\i[1294]  & ~\i[1295] ) ? ~new_n8940_ : ~new_n8942_);
  assign new_n8936_ = (~new_n6475_ & \i[2061]  & \i[2062]  & \i[2063] ) | (new_n8937_ & (~\i[2061]  | ~\i[2062]  | ~\i[2063] ));
  assign new_n8937_ = new_n4757_ ? (new_n5054_ ? ~new_n8223_ : new_n8939_) : new_n8938_;
  assign new_n8938_ = ~new_n6252_ & (\i[933]  | \i[934]  | \i[935] );
  assign new_n8939_ = \i[1086]  & \i[1087]  & (\i[1085]  | \i[1084] );
  assign new_n8940_ = (~new_n6289_ | ~new_n4381_ | new_n6280_) & (new_n8941_ | ~new_n4291_ | ~new_n6280_);
  assign new_n8941_ = \i[1735]  & (\i[1734]  | \i[1733] );
  assign new_n8942_ = (new_n8060_ | new_n7423_ | ~new_n4705_) & (new_n8943_ | \i[1063]  | ~new_n4361_ | new_n4705_);
  assign new_n8943_ = \i[1062]  & (\i[1061]  | \i[1060] );
  assign new_n8944_ = new_n8952_ ? ((~new_n8950_ & new_n3628_) | (new_n8951_ & new_n4372_ & ~new_n3628_)) : new_n8945_;
  assign new_n8945_ = new_n3550_ ? new_n8946_ : ((~new_n8949_ & new_n5408_) | (~new_n8583_ & new_n4013_ & ~new_n5408_));
  assign new_n8946_ = new_n3269_ ? (new_n5128_ ? new_n3797_ : ~new_n8948_) : new_n8947_;
  assign new_n8947_ = new_n4850_ ? (~\i[1487]  | (~\i[1485]  & ~\i[1486] )) : new_n4071_;
  assign new_n8948_ = ~\i[2863]  & (~\i[2861]  | ~\i[2862]  | ~\i[2860] );
  assign new_n8949_ = (~new_n5035_ | ~new_n5530_) & (\i[2627]  | new_n5530_ | (\i[2626]  & (\i[2624]  | \i[2625] )));
  assign new_n8950_ = new_n8411_ ? new_n7405_ : (new_n6875_ | (new_n4861_ & \i[864]  & \i[865] ));
  assign new_n8951_ = ~new_n3997_ & (~new_n6525_ | new_n3225_);
  assign new_n8952_ = \i[1423]  & (\i[1421]  | \i[1422]  | \i[1420] );
  assign new_n8953_ = new_n5098_ ? new_n8954_ : (new_n8781_ ? new_n8780_ : new_n8957_);
  assign new_n8954_ = (new_n8956_ | new_n8777_ | new_n6119_) & (~new_n6119_ | (~new_n8955_ & (new_n8775_ | new_n5408_)));
  assign new_n8955_ = new_n5408_ & (~new_n4412_ | new_n8776_) & (\i[2533]  | \i[2534]  | \i[2535]  | ~new_n8776_);
  assign new_n8956_ = new_n6417_ & ((new_n5654_ & ~new_n4094_) | (\i[2867]  & new_n4094_ & (\i[2866]  | \i[2865] )));
  assign new_n8957_ = new_n3236_ ? (new_n4954_ ? new_n3777_ : new_n3680_) : new_n8958_;
  assign new_n8958_ = (~new_n5605_ | ~\i[2763]  | (~\i[2761]  & ~\i[2762] )) & (~\i[1854]  | ~\i[1855]  | (\i[2763]  & (\i[2761]  | \i[2762] )));
  assign new_n8959_ = (new_n8960_ & ~\i[2962]  & ~\i[2963] ) | (~new_n8971_ & (new_n8969_ | new_n7751_) & (\i[2962]  | \i[2963] ));
  assign new_n8960_ = (new_n8964_ | new_n8961_ | ~new_n8968_) & (new_n8968_ | (~new_n8962_ & (new_n8967_ | new_n3437_)));
  assign new_n8961_ = (new_n4395_ | \i[847] ) & (\i[2870]  | \i[2871] ) & (~new_n3383_ | ~\i[847] );
  assign new_n8962_ = ~new_n8963_ & new_n3437_ & (\i[1847]  | \i[1846]  | ~new_n7090_);
  assign new_n8963_ = ~new_n7090_ & (\i[1627]  | \i[1626] );
  assign new_n8964_ = new_n8966_ & ~\i[2871]  & ~new_n8965_ & ~\i[2870] ;
  assign new_n8965_ = ~\i[2303]  & (~\i[2302]  | (~\i[2301]  & ~\i[2300] ));
  assign new_n8966_ = \i[2835]  & (\i[2834]  | \i[2833] );
  assign new_n8967_ = ~new_n7442_ & (~\i[1039]  | ~\i[1038] );
  assign new_n8968_ = ~\i[2978]  & ~\i[2979]  & (~\i[2977]  | ~\i[2976] );
  assign new_n8969_ = (~new_n4433_ & ~\i[1045]  & ~\i[1046]  & ~\i[1047] ) | (new_n8970_ & (\i[1045]  | \i[1046]  | \i[1047] ));
  assign new_n8970_ = new_n4016_ & (\i[2953]  | \i[2954]  | \i[2955] );
  assign new_n8971_ = new_n7751_ & new_n8972_ & (~\i[2407]  | new_n5394_);
  assign new_n8972_ = ~new_n5896_ & ((~\i[1394]  & ~\i[1393] ) | \i[2407]  | ~\i[1395] );
  assign new_n8973_ = (new_n8974_ & new_n8467_) | (~new_n8983_ & ~new_n8467_ & (~new_n5837_ | new_n8980_));
  assign new_n8974_ = (new_n8976_ | new_n8977_ | ~new_n8979_) & (new_n8979_ | (new_n3572_ ? new_n8978_ : new_n8975_));
  assign new_n8975_ = (~\i[1943]  & (~\i[1940]  | ~\i[1941]  | ~\i[1942] )) ? new_n3548_ : ~new_n4300_;
  assign new_n8976_ = new_n4393_ & (\i[2291]  | new_n4977_);
  assign new_n8977_ = new_n5394_ & ~new_n4393_ & new_n3782_;
  assign new_n8978_ = new_n3313_ ? new_n4061_ : (~\i[2307]  | (~\i[2305]  & ~\i[2306] ));
  assign new_n8979_ = ~\i[2639]  & (~\i[2637]  | ~\i[2638]  | ~\i[2636] );
  assign new_n8980_ = ~new_n8981_ & (~new_n3511_ | ~new_n8411_ | ~\i[2419]  | (~\i[2418]  & ~\i[2417] ));
  assign new_n8981_ = ~new_n8411_ & ((~new_n8982_ & ~new_n6475_) | (new_n4987_ & \i[1528]  & \i[1529]  & new_n6475_));
  assign new_n8982_ = ~\i[1802]  & ~\i[1803]  & (~\i[1801]  | ~\i[1800] );
  assign new_n8983_ = ~new_n5837_ & ~\i[2315]  & new_n8984_ & (~\i[2314]  | ~\i[2313]  | ~\i[2312] );
  assign new_n8984_ = ~new_n6406_ & new_n4842_;
  assign new_n8985_ = new_n8986_ & (\i[2674]  | \i[2675]  | \i[2673]  | (\i[2755]  & new_n5491_));
  assign new_n8986_ = new_n6799_ & (\i[1776]  | \i[1777]  | \i[1778]  | \i[1779] );
  assign new_n8987_ = new_n3258_ ? new_n8988_ : (~new_n8993_ & (new_n8995_ | new_n8996_ | new_n4186_));
  assign new_n8988_ = new_n7750_ ? ((new_n8992_ | ~new_n4494_) & (new_n7358_ | new_n8966_ | new_n4494_)) : new_n8989_;
  assign new_n8989_ = new_n4317_ ? ~new_n5456_ : (new_n8990_ ? ~new_n3326_ : new_n8991_);
  assign new_n8990_ = \i[1267]  & (\i[1265]  | \i[1266]  | \i[1264] );
  assign new_n8991_ = ~\i[2963]  & ~\i[2961]  & ~\i[2962] ;
  assign new_n8992_ = (new_n5526_ & ~new_n6252_) | (~\i[1723]  & new_n6252_ & (~\i[1722]  | ~\i[1721] ));
  assign new_n8993_ = ~new_n8994_ & new_n4186_ & (~new_n3347_ | (new_n3510_ & ~new_n3777_) | (~new_n5837_ & new_n3777_));
  assign new_n8994_ = ~new_n3347_ & ~\i[1167]  & new_n6287_ & (~\i[1166]  | new_n4932_);
  assign new_n8995_ = new_n7295_ & ((\i[743]  & new_n3536_) | (~\i[1418]  & ~\i[1419]  & ~new_n3536_));
  assign new_n8996_ = ~new_n7295_ & (new_n4657_ | ~new_n4915_) & (~\i[1481]  | ~\i[1482]  | ~\i[1483]  | new_n4915_);
  assign new_n8997_ = (new_n8998_ & ~new_n7746_) | (~new_n9001_ & new_n7746_ & (new_n9002_ | (~new_n9003_ & ~new_n9006_)));
  assign new_n8998_ = new_n5156_ ? ~new_n8999_ : (new_n5665_ ? ~new_n3855_ : new_n9000_);
  assign new_n8999_ = new_n3661_ & new_n4166_ & (\i[509]  | \i[508] );
  assign new_n9000_ = (~\i[1539]  | ~\i[2083] ) & (\i[2424]  | \i[2425]  | \i[2426]  | \i[2427]  | \i[2083] );
  assign new_n9001_ = new_n9002_ & (~new_n3731_ | ~new_n4062_ | new_n7386_) & (~new_n7969_ | ~new_n6690_ | ~new_n7386_);
  assign new_n9002_ = ~\i[2383]  & (~\i[2382]  | ~\i[2381] );
  assign new_n9003_ = ~new_n9005_ & (new_n4694_ | ~new_n9004_) & (\i[2817]  | \i[2818]  | \i[2819]  | new_n9004_);
  assign new_n9004_ = \i[823]  & (\i[822]  | \i[821] );
  assign new_n9005_ = \i[1431]  & \i[1430]  & \i[1428]  & \i[1429] ;
  assign new_n9006_ = \i[1323]  & \i[1322]  & new_n5609_ & new_n9005_;
  assign new_n9007_ = new_n3223_ ? new_n9008_ : (~new_n9012_ & (new_n6289_ | new_n9014_ | ~new_n9015_));
  assign new_n9008_ = new_n7028_ ? (~new_n9010_ & (new_n9011_ | ~new_n5584_ | ~new_n4449_)) : new_n9009_;
  assign new_n9009_ = (~new_n6469_ | ~new_n5041_ | new_n6240_) & (new_n7496_ | ~\i[2958]  | ~\i[2959]  | ~new_n6240_);
  assign new_n9010_ = new_n4843_ & new_n9011_ & ((\i[2876]  & \i[2877] ) | \i[2879]  | \i[2878] );
  assign new_n9011_ = ~\i[1527]  & ~\i[1525]  & ~\i[1526] ;
  assign new_n9012_ = new_n9014_ & (\i[2767]  ? (~new_n3687_ | new_n3229_) : new_n9013_);
  assign new_n9013_ = new_n8363_ ? (\i[2759]  | (\i[2757]  & \i[2758] )) : ~new_n5231_;
  assign new_n9014_ = ~\i[2830]  & ~\i[2831] ;
  assign new_n9015_ = ~\i[1507]  & (~\i[1506]  | ~\i[1505] );
  assign new_n9016_ = new_n6437_ ? new_n9017_ : (new_n9023_ | (~new_n9022_ & ~\i[995] ));
  assign new_n9017_ = (new_n9021_ | new_n9018_ | ~new_n3478_) & (new_n3478_ | (new_n5684_ ? new_n9020_ : new_n9019_));
  assign new_n9018_ = ~new_n6459_ & (~\i[1479]  | (~\i[1476]  & ~\i[1477]  & ~\i[1478] ));
  assign new_n9019_ = (~\i[1491]  | ~new_n5238_ | (~\i[1490]  & (~\i[1488]  | ~\i[1489] ))) & (new_n3497_ | new_n5238_);
  assign new_n9020_ = new_n6873_ & (\i[760]  | \i[761]  | \i[762]  | \i[763] );
  assign new_n9021_ = \i[1846]  & \i[1847]  & (\i[1845]  | \i[1844] );
  assign new_n9022_ = \i[829]  & \i[828]  & new_n6885_ & ~\i[839]  & ~\i[837]  & ~\i[838] ;
  assign new_n9023_ = \i[1039]  & \i[1038]  & \i[1036]  & \i[1037] ;
  assign \o[64]  = new_n9025_ ? (new_n9026_ ^ new_n9027_) : (~new_n9026_ ^ new_n9027_);
  assign new_n9025_ = (~new_n9007_ & ~new_n9016_) | (~new_n8714_ & (~new_n9007_ | ~new_n9016_));
  assign new_n9026_ = (~new_n8987_ & ~new_n8997_) | (~new_n8715_ & (~new_n8987_ | ~new_n8997_));
  assign new_n9027_ = new_n9028_ ? (~new_n9029_ ^ new_n9122_) : (new_n9029_ ^ new_n9122_);
  assign new_n9028_ = (~new_n8912_ & ~new_n8985_) | (~new_n8716_ & (~new_n8912_ | ~new_n8985_));
  assign new_n9029_ = new_n9030_ ? (new_n9050_ ^ new_n9051_) : (~new_n9050_ ^ new_n9051_);
  assign new_n9030_ = new_n9031_ ? (~new_n9032_ ^ new_n9049_) : (new_n9032_ ^ new_n9049_);
  assign new_n9031_ = (~new_n8782_ & ~new_n8790_) | (~new_n8718_ & (~new_n8782_ | ~new_n8790_));
  assign new_n9032_ = new_n9033_ ? (~new_n9044_ ^ new_n9045_) : (new_n9044_ ^ new_n9045_);
  assign new_n9033_ = new_n9034_ ? (~new_n9035_ ^ new_n9036_) : (new_n9035_ ^ new_n9036_);
  assign new_n9034_ = (~new_n8728_ & ~new_n8739_) | (~new_n8720_ & (~new_n8728_ | ~new_n8739_));
  assign new_n9035_ = (~new_n8930_ & new_n8922_) | (new_n8916_ & (~new_n8930_ | new_n8922_));
  assign new_n9036_ = new_n9037_ ? (~new_n9041_ ^ new_n9043_) : (new_n9041_ ^ new_n9043_);
  assign new_n9037_ = new_n7925_ ? new_n9038_ : (new_n8907_ ? new_n9040_ : ~new_n9039_);
  assign new_n9038_ = (~new_n8909_ | ~\i[2987]  | ~new_n7933_) & (new_n4244_ | ~new_n8621_ | new_n7933_);
  assign new_n9039_ = ~new_n4080_ & new_n8738_ & (~new_n4049_ | (~\i[1080]  & ~\i[1081] ));
  assign new_n9040_ = (new_n3445_ | ~new_n4356_ | new_n8905_) & (new_n3368_ | ~new_n8905_ | (\i[2749]  & new_n4803_));
  assign new_n9041_ = (new_n7031_ | new_n5387_ | ~new_n8750_ | ~new_n8734_) & (~new_n9042_ | new_n5930_ | new_n8734_);
  assign new_n9042_ = ~\i[1631]  & ~\i[935]  & ~\i[1630]  & \i[2623]  & (\i[2622]  | \i[2621] );
  assign new_n9043_ = (new_n8753_ | ~new_n8789_) & (~new_n4792_ | ~new_n7993_ | ~new_n8787_ | new_n8789_);
  assign new_n9044_ = (~new_n8772_ & ~new_n8935_) | (~new_n8915_ & (~new_n8772_ | ~new_n8935_));
  assign new_n9045_ = new_n7925_ & ((~new_n5479_ & new_n9046_ & new_n8734_) | (~new_n9047_ & new_n9048_ & ~new_n8734_));
  assign new_n9046_ = \i[1539]  & \i[1538]  & \i[1537]  & ~new_n3562_ & \i[1536] ;
  assign new_n9047_ = ~new_n8731_ & ~\i[1183] ;
  assign new_n9048_ = ~new_n4895_ & ~new_n5665_;
  assign new_n9049_ = (~new_n8944_ & ~new_n8953_) | (~new_n8914_ & (~new_n8944_ | ~new_n8953_));
  assign new_n9050_ = (~new_n8796_ & ~new_n8901_) | (~new_n8717_ & (~new_n8796_ | ~new_n8901_));
  assign new_n9051_ = new_n9052_ ? (new_n9077_ ^ new_n9078_) : (~new_n9077_ ^ new_n9078_);
  assign new_n9052_ = new_n9053_ ? (~new_n9054_ ^ new_n9055_) : (new_n9054_ ^ new_n9055_);
  assign new_n9053_ = (~new_n8745_ & ~new_n8772_) | (~new_n8719_ & (~new_n8745_ | ~new_n8772_));
  assign new_n9054_ = (~new_n8894_ & new_n8865_) | (~new_n8867_ & (~new_n8894_ | new_n8865_));
  assign new_n9055_ = new_n9056_ ? (new_n9065_ ^ new_n9076_) : (~new_n9065_ ^ new_n9076_);
  assign new_n9056_ = new_n9057_ ? (new_n9060_ ^ new_n9064_) : (~new_n9060_ ^ new_n9064_);
  assign new_n9057_ = ~new_n8826_ & (new_n8832_ | (~\i[1831]  & new_n7442_) | (~new_n9059_ & ~new_n9058_ & ~new_n7442_));
  assign new_n9058_ = ~new_n8835_ & (new_n8836_ ? ~new_n3445_ : ~new_n4238_);
  assign new_n9059_ = ~new_n3544_ & new_n8835_ & \i[2199]  & (\i[2198]  | (\i[2196]  & \i[2197] ));
  assign new_n9060_ = new_n3843_ ? (new_n4377_ ? new_n9063_ : ~new_n8880_) : new_n9061_;
  assign new_n9061_ = (~new_n8888_ & (~\i[1258]  | ~\i[1259] )) | (~new_n9062_ & \i[1258]  & \i[1259]  & (new_n8884_ | ~new_n6828_));
  assign new_n9062_ = ~new_n6828_ & (new_n8887_ ? ~new_n6887_ : new_n4160_);
  assign new_n9063_ = new_n8884_ ? ~new_n8885_ : (new_n6266_ ? ~new_n3351_ : new_n7421_);
  assign new_n9064_ = new_n8986_ & (\i[2673]  | \i[2674]  | \i[2675] );
  assign new_n9065_ = new_n9066_ ? (~new_n9070_ ^ new_n9073_) : (new_n9070_ ^ new_n9073_);
  assign new_n9066_ = (~\i[2962]  & ~\i[2963] ) ? (new_n9069_ | new_n8968_) : new_n9067_;
  assign new_n9067_ = (new_n8972_ | ~new_n7751_) & (new_n9068_ | \i[1045]  | \i[1046]  | \i[1047]  | new_n7751_);
  assign new_n9068_ = new_n4433_ & \i[1415]  & (\i[1414]  | (\i[1412]  & \i[1413] ));
  assign new_n9069_ = new_n3437_ ? ~new_n8963_ : ~new_n8967_;
  assign new_n9070_ = (new_n5837_ | new_n9072_ | ~new_n8984_ | new_n8467_) & (~new_n8979_ | new_n9071_ | ~new_n8467_);
  assign new_n9071_ = ~new_n8977_ & (~new_n4393_ | ~\i[743]  | ~\i[2291]  | (~\i[742]  & ~new_n8207_));
  assign new_n9072_ = ~\i[2315]  & (~\i[2313]  | ~\i[2314]  | ~\i[2312] );
  assign new_n9073_ = (new_n7338_ | new_n8753_ | ~new_n3793_ | ~new_n8789_) & (~new_n9074_ | new_n9075_ | new_n8789_);
  assign new_n9074_ = ~new_n5080_ & ~\i[987]  & (~\i[986]  | ~\i[985] );
  assign new_n9075_ = ~\i[2833]  & new_n5480_;
  assign new_n9076_ = (~new_n8756_ & ~new_n8763_) | (new_n8746_ & (~new_n8756_ | ~new_n8763_));
  assign new_n9077_ = (~new_n8866_ & ~new_n8790_) | (~new_n8797_ & (~new_n8866_ | ~new_n8790_));
  assign new_n9078_ = new_n9079_ ? (new_n9091_ ^ new_n9092_) : (~new_n9091_ ^ new_n9092_);
  assign new_n9079_ = new_n9080_ ? (~new_n9081_ ^ new_n9082_) : (new_n9081_ ^ new_n9082_);
  assign new_n9080_ = (~new_n8877_ & ~new_n8889_) | (new_n8868_ & (~new_n8877_ | ~new_n8889_));
  assign new_n9081_ = (~new_n8854_ & new_n8838_) | (new_n8825_ & (~new_n8854_ | new_n8838_));
  assign new_n9082_ = new_n9083_ ? (~new_n9086_ ^ new_n9089_) : (new_n9086_ ^ new_n9089_);
  assign new_n9083_ = (new_n9084_ | ~new_n3258_) & (~new_n4657_ | ~new_n4915_ | new_n3258_ | new_n4186_ | new_n7295_);
  assign new_n9084_ = (~new_n9085_ | new_n7750_) & (new_n6132_ | new_n4494_ | ~new_n8966_ | ~new_n7750_);
  assign new_n9085_ = ~new_n5456_ & new_n4317_ & ((\i[1588]  & \i[1589] ) | \i[1591]  | \i[1590] );
  assign new_n9086_ = ~new_n9087_ & (~new_n9005_ | ~new_n9088_ | ~new_n7746_ | (\i[1323]  & \i[1322] ));
  assign new_n9087_ = new_n3855_ & new_n5804_ & new_n5665_ & ~new_n5156_ & ~new_n7746_;
  assign new_n9088_ = ~new_n9002_ & (\i[1643]  | (\i[1641]  & \i[1642] ));
  assign new_n9089_ = (~new_n9090_ | new_n4179_) & (new_n3220_ | new_n5238_ | new_n8859_ | ~new_n3290_ | ~new_n4179_);
  assign new_n9090_ = \i[2427]  & \i[2426]  & \i[2425]  & ~new_n3506_ & \i[2424] ;
  assign new_n9091_ = (~new_n8824_ & new_n8865_) | (~new_n8798_ & (~new_n8824_ | new_n8865_));
  assign new_n9092_ = new_n9093_ ? (~new_n9094_ ^ new_n9109_) : (new_n9094_ ^ new_n9109_);
  assign new_n9093_ = ~new_n8813_ & new_n8799_;
  assign new_n9094_ = new_n9095_ ? (~new_n9100_ ^ new_n9105_) : (new_n9100_ ^ new_n9105_);
  assign new_n9095_ = (new_n9096_ & new_n6437_) | (~new_n8850_ & ~new_n9099_ & ~new_n6437_);
  assign new_n9096_ = new_n8853_ ? (new_n6316_ ? new_n8840_ : ~new_n8841_) : new_n9097_;
  assign new_n9097_ = (new_n9098_ | ~new_n8844_) & (~new_n6539_ | ~new_n8846_ | new_n8844_);
  assign new_n9098_ = ~new_n8845_ & (~new_n3254_ | ~\i[714]  | ~\i[715] );
  assign new_n9099_ = new_n8848_ & ((new_n3754_ & ~new_n8849_) | (new_n3647_ & new_n5777_ & new_n8849_));
  assign new_n9100_ = new_n5079_ ? new_n9101_ : ((new_n7842_ | new_n9104_) & (~new_n8822_ | ~new_n9103_));
  assign new_n9101_ = ~new_n9102_ & (~new_n8817_ | (new_n6375_ & (~new_n6143_ | new_n4343_)));
  assign new_n9102_ = new_n5763_ & ((~new_n3488_ & new_n8816_) | (~new_n6155_ & new_n4331_ & ~new_n8816_));
  assign new_n9103_ = new_n7842_ & new_n4134_ & \i[2711]  & (\i[2710]  | \i[2709]  | \i[2708] );
  assign new_n9104_ = (~new_n4273_ | ~new_n4036_ | ~new_n3414_) & (~new_n4806_ | new_n3414_ | (~\i[867]  & ~\i[866] ));
  assign new_n9105_ = (~new_n9023_ | ~new_n8849_ | new_n6437_) & (new_n9106_ | ~new_n3478_ | ~new_n9021_ | ~new_n6437_);
  assign new_n9106_ = (new_n9108_ & new_n9107_) | (~\i[2890]  & ~\i[2891]  & ~new_n9107_ & (~\i[2889]  | ~\i[2888] ));
  assign new_n9107_ = \i[1647]  & (\i[1646]  | (\i[1645]  & \i[1644] ));
  assign new_n9108_ = ~\i[1379]  & (~\i[1377]  | ~\i[1378]  | ~\i[1376] );
  assign new_n9109_ = ~new_n9110_ ^ new_n9117_;
  assign new_n9110_ = new_n3223_ ? (new_n7028_ ? ~new_n9113_ : ~new_n9111_) : new_n9114_;
  assign new_n9111_ = (new_n9112_ | ~new_n7496_ | ~new_n6240_) & (new_n6240_ | (new_n5041_ ? new_n6469_ : ~new_n5094_));
  assign new_n9112_ = ~\i[955]  & (~\i[952]  | ~new_n3249_);
  assign new_n9113_ = (new_n4843_ | new_n3592_ | ~new_n9011_) & (new_n4449_ | new_n7032_ | new_n9011_);
  assign new_n9114_ = (new_n9115_ & ~new_n9014_) | (~new_n3687_ & \i[2094]  & \i[2095]  & \i[2767]  & new_n9014_);
  assign new_n9115_ = (new_n6948_ | ~new_n6289_ | ~new_n9015_) & (new_n9116_ | ~new_n6926_ | new_n9015_);
  assign new_n9116_ = \i[2178]  & \i[2179]  & (\i[2177]  | \i[2176] );
  assign new_n9117_ = new_n8812_ ? ((new_n9118_ | ~new_n5896_) & (new_n9121_ | ~new_n8802_ | new_n5896_)) : new_n9120_;
  assign new_n9118_ = (new_n9119_ | ~new_n8805_) & (new_n3994_ | ~new_n8806_ | new_n8805_);
  assign new_n9119_ = (new_n4361_ & (\i[2880]  | \i[2881]  | \i[2882]  | \i[2883] )) | (new_n3710_ & ~\i[2880]  & ~\i[2881]  & ~\i[2882]  & ~\i[2883] );
  assign new_n9120_ = (~new_n5802_ | ~new_n7212_ | ~new_n4757_ | ~new_n4215_) & (~new_n7287_ | ~new_n6093_ | new_n4215_);
  assign new_n9121_ = ~new_n6085_ & ((\i[821]  & \i[820] ) | \i[823]  | \i[822] );
  assign new_n9122_ = (~new_n8959_ & ~new_n8973_) | (~new_n8913_ & (~new_n8959_ | ~new_n8973_));
  assign \o[65]  = ~new_n9124_ ^ new_n9125_;
  assign new_n9124_ = (~new_n9027_ & new_n9026_) | (new_n9025_ & (~new_n9027_ | new_n9026_));
  assign new_n9125_ = new_n9126_ ^ new_n9127_;
  assign new_n9126_ = (~new_n9029_ & new_n9122_) | (new_n9028_ & (~new_n9029_ | new_n9122_));
  assign new_n9127_ = new_n9128_ ? (~new_n9129_ ^ new_n9162_) : (new_n9129_ ^ new_n9162_);
  assign new_n9128_ = (~new_n9051_ & new_n9050_) | (~new_n9030_ & (~new_n9051_ | new_n9050_));
  assign new_n9129_ = new_n9130_ ? (new_n9138_ ^ new_n9139_) : (~new_n9138_ ^ new_n9139_);
  assign new_n9130_ = new_n9131_ ? (~new_n9132_ ^ new_n9133_) : (new_n9132_ ^ new_n9133_);
  assign new_n9131_ = (~new_n9055_ & new_n9054_) | (new_n9053_ & (~new_n9055_ | new_n9054_));
  assign new_n9132_ = (new_n9044_ & new_n9045_) | (~new_n9033_ & (new_n9044_ | new_n9045_));
  assign new_n9133_ = new_n9134_ ^ new_n9135_;
  assign new_n9134_ = (~new_n9036_ & new_n9035_) | (new_n9034_ & (~new_n9036_ | new_n9035_));
  assign new_n9135_ = ~new_n9136_ ^ new_n9137_;
  assign new_n9136_ = (~new_n9070_ & ~new_n9073_) | (~new_n9066_ & (~new_n9070_ | ~new_n9073_));
  assign new_n9137_ = (~new_n9041_ & ~new_n9043_) | (~new_n9037_ & (~new_n9041_ | ~new_n9043_));
  assign new_n9138_ = (~new_n9078_ & new_n9077_) | (~new_n9052_ & (~new_n9078_ | new_n9077_));
  assign new_n9139_ = new_n9140_ ? (new_n9144_ ^ new_n9145_) : (~new_n9144_ ^ new_n9145_);
  assign new_n9140_ = new_n9141_ ? (new_n9142_ ^ new_n9143_) : (~new_n9142_ ^ new_n9143_);
  assign new_n9141_ = (~new_n9082_ & new_n9081_) | (new_n9080_ & (~new_n9082_ | new_n9081_));
  assign new_n9142_ = (~new_n9065_ & new_n9076_) | (~new_n9056_ & (~new_n9065_ | new_n9076_));
  assign new_n9143_ = (~new_n9060_ & new_n9064_) | (~new_n9057_ & (~new_n9060_ | new_n9064_));
  assign new_n9144_ = (~new_n9092_ & new_n9091_) | (~new_n9079_ & (~new_n9092_ | new_n9091_));
  assign new_n9145_ = new_n9146_ ? (new_n9147_ ^ new_n9150_) : (~new_n9147_ ^ new_n9150_);
  assign new_n9146_ = (~new_n9094_ & ~new_n9109_) | (~new_n9093_ & (~new_n9094_ | ~new_n9109_));
  assign new_n9147_ = ~new_n9148_ ^ new_n9149_;
  assign new_n9148_ = (~new_n9100_ & ~new_n9105_) | (~new_n9095_ & (~new_n9100_ | ~new_n9105_));
  assign new_n9149_ = (~new_n9086_ & ~new_n9089_) | (~new_n9083_ & (~new_n9086_ | ~new_n9089_));
  assign new_n9150_ = new_n9151_ ? (~new_n9152_ ^ new_n9161_) : (new_n9152_ ^ new_n9161_);
  assign new_n9151_ = ~new_n9110_ & new_n9117_;
  assign new_n9152_ = new_n9153_ ^ new_n9159_;
  assign new_n9153_ = (new_n9155_ | new_n9154_ | ~new_n8812_) & (new_n8812_ | (new_n4215_ ? new_n9157_ : new_n9158_));
  assign new_n9154_ = ~new_n5896_ & (new_n4520_ ? (new_n8398_ ? new_n6856_ : ~new_n5626_) : ~new_n8803_);
  assign new_n9155_ = new_n5896_ & (new_n8805_ ? ~new_n9156_ : (new_n8806_ | new_n4356_));
  assign new_n9156_ = ~new_n4361_ & (\i[2880]  | \i[2881]  | \i[2882]  | \i[2883] );
  assign new_n9157_ = (new_n6101_ | new_n7212_) & (new_n5802_ | new_n5156_ | ~new_n7212_);
  assign new_n9158_ = (~new_n7810_ | ~new_n8809_ | new_n7287_) & (~new_n7287_ | (new_n6093_ ? new_n6296_ : new_n5200_));
  assign new_n9159_ = ~new_n3223_ & (new_n9160_ | (~new_n5231_ & ~new_n8363_ & ~\i[2767]  & new_n9014_));
  assign new_n9160_ = new_n6061_ & ~new_n9014_ & ~new_n6926_ & ~new_n9015_;
  assign new_n9161_ = new_n4238_ & ~new_n8836_ & ~new_n8835_ & ~new_n7442_ & ~new_n8832_;
  assign new_n9162_ = (~new_n9032_ & new_n9049_) | (new_n9031_ & (~new_n9032_ | new_n9049_));
  assign \o[66]  = ((new_n9164_ | new_n9165_) & (~new_n9166_ ^ ~new_n9167_)) | (~new_n9164_ & ~new_n9165_ & (~new_n9166_ ^ new_n9167_));
  assign new_n9164_ = ~new_n9125_ & new_n9124_;
  assign new_n9165_ = ~new_n9127_ & new_n9126_;
  assign new_n9166_ = (~new_n9129_ & new_n9162_) | (new_n9128_ & (~new_n9129_ | new_n9162_));
  assign new_n9167_ = new_n9168_ ? (~new_n9169_ ^ new_n9181_) : (new_n9169_ ^ new_n9181_);
  assign new_n9168_ = (~new_n9139_ & new_n9138_) | (~new_n9130_ & (~new_n9139_ | new_n9138_));
  assign new_n9169_ = new_n9170_ ? (new_n9174_ ^ new_n9175_) : (~new_n9174_ ^ new_n9175_);
  assign new_n9170_ = new_n9171_ ? (new_n9172_ ^ new_n9173_) : (~new_n9172_ ^ new_n9173_);
  assign new_n9171_ = (new_n9142_ & new_n9143_) | (new_n9141_ & (new_n9142_ | new_n9143_));
  assign new_n9172_ = ~new_n9135_ & new_n9134_;
  assign new_n9173_ = new_n9136_ & new_n9137_;
  assign new_n9174_ = (~new_n9145_ & new_n9144_) | (~new_n9140_ & (~new_n9145_ | new_n9144_));
  assign new_n9175_ = new_n9176_ ? (~new_n9177_ ^ new_n9180_) : (new_n9177_ ^ new_n9180_);
  assign new_n9176_ = (~new_n9147_ & ~new_n9150_) | (new_n9146_ & (~new_n9147_ | ~new_n9150_));
  assign new_n9177_ = new_n9178_ ^ new_n9179_;
  assign new_n9178_ = (new_n9152_ & new_n9161_) | (~new_n9151_ & (new_n9152_ | new_n9161_));
  assign new_n9179_ = ~new_n9159_ & new_n9153_;
  assign new_n9180_ = new_n9148_ & new_n9149_;
  assign new_n9181_ = (~new_n9133_ & new_n9132_) | (new_n9131_ & (~new_n9133_ | new_n9132_));
  assign \o[67]  = ~new_n9183_ ^ new_n9184_;
  assign new_n9183_ = (new_n9166_ | (~new_n9167_ & (new_n9165_ | new_n9164_))) & (new_n9165_ | new_n9164_ | ~new_n9167_);
  assign new_n9184_ = new_n9185_ ^ new_n9186_;
  assign new_n9185_ = (~new_n9169_ & new_n9181_) | (new_n9168_ & (~new_n9169_ | new_n9181_));
  assign new_n9186_ = new_n9187_ ? (~new_n9188_ ^ new_n9191_) : (new_n9188_ ^ new_n9191_);
  assign new_n9187_ = (~new_n9175_ & new_n9174_) | (~new_n9170_ & (~new_n9175_ | new_n9174_));
  assign new_n9188_ = ~new_n9189_ ^ new_n9190_;
  assign new_n9189_ = (~new_n9177_ & new_n9180_) | (new_n9176_ & (~new_n9177_ | new_n9180_));
  assign new_n9190_ = ~new_n9179_ & new_n9178_;
  assign new_n9191_ = (new_n9172_ & new_n9173_) | (new_n9171_ & (new_n9172_ | new_n9173_));
  assign \o[68]  = ((new_n9193_ | new_n9194_) & (~new_n9195_ ^ new_n9196_)) | (~new_n9193_ & ~new_n9194_ & (~new_n9195_ ^ ~new_n9196_));
  assign new_n9193_ = ~new_n9184_ & new_n9183_;
  assign new_n9194_ = ~new_n9186_ & new_n9185_;
  assign new_n9195_ = (~new_n9188_ & new_n9191_) | (new_n9187_ & (~new_n9188_ | new_n9191_));
  assign new_n9196_ = new_n9189_ & new_n9190_;
  assign \o[69]  = (new_n9196_ | new_n9193_ | new_n9194_) & (new_n9195_ | (new_n9196_ & (new_n9193_ | new_n9194_)));
endmodule


